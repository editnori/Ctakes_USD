 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Procedure|Health Care Activity|SIMPLE_SEGMENT|46,55|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|46,60|false|false|false|C2598112||Admission Date
Finding|Body Substance|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|80,89|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|80,94|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|136,139|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|147,154|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|147,154|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Attribute|Clinical Attribute|SIMPLE_SEGMENT|167,176|false|false|false|C1717415||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|167,176|false|false|false|C0020517|Hypersensitivity|Allergies
Finding|Body Substance|SIMPLE_SEGMENT|179,186|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|179,186|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|179,186|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Attribute|Clinical Attribute|SIMPLE_SEGMENT|215,224|true|false|false|C1717415||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|215,224|true|false|false|C0020517|Hypersensitivity|Allergies
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|228,233|false|false|false|C0013227|Pharmaceutical Preparations|Drugs
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|228,233|false|false|false|C3687832|Drugs - dental services|Drugs
Finding|Functional Concept|SIMPLE_SEGMENT|236,245|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|254,269|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|260,269|false|false|false|C3864418||Complaint
Finding|Finding|SIMPLE_SEGMENT|260,269|false|false|false|C5441521|Complaint (finding)|Complaint
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|273,282|false|false|false|C0751438|Posterior pituitary disease|posterior
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|273,300|false|false|false|C0554595|Tibialis posterior tendinitis|posterior tibial tendonitis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|283,289|false|false|false|C0040184|Bone structure of tibia|tibial
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|290,300|false|false|false|C0039503|Tendinitis|tendonitis
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|301,305|false|false|false|C0043246;C3203359|Laceration;Rupture|tear
Finding|Body Substance|SIMPLE_SEGMENT|301,305|false|false|false|C0039409|Tears (substance)|tear
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|308,314|false|false|false|C1550316|Tarsal|tarsal
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|308,321|false|false|false|C0225150|Structure of tarsal canal|tarsal tunnel
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|308,329|false|false|false|C0196577|Decompression of tarsal tunnel|tarsal tunnel release
Finding|Functional Concept|SIMPLE_SEGMENT|322,329|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|release
Procedure|Health Care Activity|SIMPLE_SEGMENT|322,329|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|322,329|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|release
Finding|Classification|SIMPLE_SEGMENT|332,337|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|338,346|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|338,346|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|350,368|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|359,368|false|false|false|C0945766||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|359,368|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|359,368|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|359,368|false|false|false|C0184661|Interventional procedure|Procedure
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|376,382|false|false|false|C0039508|Tendon structure|tendon
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|376,389|false|false|false|C0565350|Plastic repair of tendon|tendon repair
Finding|Functional Concept|SIMPLE_SEGMENT|383,389|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Finding|Organism Function|SIMPLE_SEGMENT|383,389|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Procedure|Health Care Activity|SIMPLE_SEGMENT|383,389|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|383,389|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|392,398|false|false|false|C1550316|Tarsal|tarsal
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|392,405|false|false|false|C0225150|Structure of tarsal canal|tarsal tunnel
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|392,413|false|false|false|C0196577|Decompression of tarsal tunnel|tarsal tunnel release
Finding|Functional Concept|SIMPLE_SEGMENT|406,413|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|release
Procedure|Health Care Activity|SIMPLE_SEGMENT|406,413|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|406,413|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|release
Finding|Conceptual Entity|SIMPLE_SEGMENT|417,424|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|417,424|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|417,424|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|417,427|false|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|417,443|false|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|417,443|false|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|428,435|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|428,435|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|428,443|false|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|436,443|false|false|false|C0221423|Illness (finding)|Illness
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|458,461|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|458,461|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|458,461|false|false|false|C1504769|DFFB protein, human|CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|458,461|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|458,461|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|458,461|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|458,461|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|463,466|false|false|false|C0020538|Hypertensive disease|HTN
Finding|Functional Concept|SIMPLE_SEGMENT|503,513|false|false|false|C1947976|Correction (change)|correction
Finding|Functional Concept|SIMPLE_SEGMENT|521,525|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|526,535|false|false|false|C0751438|Posterior pituitary disease|posterior
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|536,542|false|false|false|C0040184|Bone structure of tibia|tibial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|543,549|false|false|false|C0039508|Tendon structure|tendon
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|556,562|false|false|false|C1550316|Tarsal|tarsal
Finding|Functional Concept|SIMPLE_SEGMENT|570,577|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|release
Procedure|Health Care Activity|SIMPLE_SEGMENT|570,577|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|570,577|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|release
Finding|Intellectual Product|SIMPLE_SEGMENT|587,595|false|false|false|C2984058|Have Pain|had pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|591,595|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|591,595|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|591,595|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Functional Concept|SIMPLE_SEGMENT|603,607|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|603,612|false|false|false|C0230461|Structure of left foot|left foot
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|608,612|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|608,612|false|false|false|C0555980|Foot problem|foot
Finding|Finding|SIMPLE_SEGMENT|628,632|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|628,632|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|628,632|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Gene or Genome|SIMPLE_SEGMENT|637,640|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|637,640|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|SIMPLE_SEGMENT|637,640|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Finding|Finding|SIMPLE_SEGMENT|652,660|false|false|false|C0332149|Possible|possible
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|661,665|false|false|false|C0043246;C3203359|Laceration;Rupture|tear
Finding|Body Substance|SIMPLE_SEGMENT|661,665|false|false|false|C0039409|Tears (substance)|tear
Finding|Gene or Genome|SIMPLE_SEGMENT|697,702|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|703,712|false|false|false|C0751438|Posterior pituitary disease|posterior
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|713,717|false|false|false|C0043246;C3203359|Laceration;Rupture|tear
Finding|Body Substance|SIMPLE_SEGMENT|713,717|false|false|false|C0039409|Tears (substance)|tear
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|729,735|false|false|false|C0039508|Tendon structure|tendon
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|746,752|false|false|false|C1550316|Tarsal|tarsal
Finding|Functional Concept|SIMPLE_SEGMENT|760,767|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|release
Procedure|Health Care Activity|SIMPLE_SEGMENT|760,767|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|760,767|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|release
Finding|Finding|SIMPLE_SEGMENT|781,785|false|false|false|C0241158;C1419736;C2004491|Cicatrix;RPS4X gene;Scar Tissue|scar
Finding|Gene or Genome|SIMPLE_SEGMENT|781,785|false|false|false|C0241158;C1419736;C2004491|Cicatrix;RPS4X gene;Scar Tissue|scar
Finding|Pathologic Function|SIMPLE_SEGMENT|781,785|false|false|false|C0241158;C1419736;C2004491|Cicatrix;RPS4X gene;Scar Tissue|scar
Finding|Finding|SIMPLE_SEGMENT|781,792|false|false|false|C0241158;C2004491|Cicatrix;Scar Tissue|scar tissue
Finding|Pathologic Function|SIMPLE_SEGMENT|781,792|false|false|false|C0241158;C2004491|Cicatrix;Scar Tissue|scar tissue
Anatomy|Tissue|SIMPLE_SEGMENT|786,792|false|false|false|C0040300|Body tissue|tissue
Finding|Intellectual Product|SIMPLE_SEGMENT|786,792|false|false|false|C1547928|Tissue Specimen Code|tissue
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|811,817|false|false|false|C0040184|Bone structure of tibia|tibial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|818,823|false|false|false|C0027740|Nerve|nerve
Finding|Conceptual Entity|SIMPLE_SEGMENT|835,842|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|835,842|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|835,842|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|835,845|false|false|false|C0262926|Medical History|history of
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|846,855|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|846,855|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|846,855|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Body Substance|SIMPLE_SEGMENT|885,892|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|885,892|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|885,892|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|SIMPLE_SEGMENT|933,937|false|false|false|C0947322;C1881534|Make - Instruction Imperative;Manufacturer Name|make
Finding|Intellectual Product|SIMPLE_SEGMENT|933,937|false|false|false|C0947322;C1881534|Make - Instruction Imperative;Manufacturer Name|make
Finding|Intellectual Product|SIMPLE_SEGMENT|939,943|false|false|false|C4724437|SURE Test|sure
Finding|Idea or Concept|SIMPLE_SEGMENT|962,970|false|true|false|C1546466|Problems - What subject filter|problems
Finding|Finding|SIMPLE_SEGMENT|977,997|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Finding|Functional Concept|SIMPLE_SEGMENT|982,989|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|982,989|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|982,989|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|982,989|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|982,997|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|990,997|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|990,997|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|990,997|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|999,1005|false|false|false|C0004096|Asthma|asthma
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1007,1016|false|false|false|C0034067|Pulmonary Emphysema|emphysema
Finding|Pathologic Function|SIMPLE_SEGMENT|1007,1016|false|false|false|C0013990|Pathological accumulation of air in tissues|emphysema
Finding|Intellectual Product|SIMPLE_SEGMENT|1018,1025|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|1018,1025|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1018,1036|false|false|false|C0008677|Bronchitis, Chronic|chronic bronchitis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1026,1036|false|false|false|C0006277;C0149514|Acute bronchitis;Bronchitis|bronchitis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1038,1041|false|false|false|C0020538|Hypertensive disease|HTN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1043,1046|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1043,1046|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|1043,1046|false|false|false|C1504769|DFFB protein, human|CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|1043,1046|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1043,1046|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|1043,1046|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1043,1046|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1056,1063|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|1056,1063|false|false|false|C1314974|Cardiac attachment|cardiac
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1076,1085|false|false|false|C0149931|Migraine Disorders|migraines
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1087,1091|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1103,1108|false|false|false|C0994475|Pills|pills
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1113,1120|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|1113,1120|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1113,1120|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|1113,1120|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1113,1120|false|false|false|C0202098|Insulin measurement|insulin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1123,1129|false|false|false|C0002871|Anemia|Anemia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1131,1141|false|false|false|C0442874|Neuropathy|neuropathy
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1143,1150|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|1143,1150|false|false|false|C0860603|Anxiety symptoms|anxiety
Finding|Functional Concept|SIMPLE_SEGMENT|1154,1160|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|1154,1168|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1161,1168|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1161,1168|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1161,1168|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|1174,1180|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|1174,1180|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|1174,1180|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|1174,1180|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|1174,1188|false|false|false|C0241889|Family Medical History|Family History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1181,1188|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1181,1188|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1181,1188|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1218,1221|false|false|false|C0020538|Hypertensive disease|htn
Finding|Finding|SIMPLE_SEGMENT|1227,1235|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|1227,1235|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1227,1235|false|false|false|C0031809|Physical Examination|Physical
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1241,1251|false|false|false|C0550215||Appearance
Procedure|Health Care Activity|SIMPLE_SEGMENT|1241,1251|false|false|false|C2051406|patient appearance regarding mental status exam|Appearance
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1253,1256|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1253,1256|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1253,1256|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|1253,1256|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1253,1256|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Finding|Finding|SIMPLE_SEGMENT|1253,1256|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1257,1262|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1270,1275|false|false|false|C0018787;C4037974|Chest>Heart;Heart|Heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1270,1275|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|Heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|1270,1275|false|false|false|C0795691|HEART PROBLEM|Heart
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1281,1286|false|false|false|C0024109|Lung|Lungs
Finding|Finding|SIMPLE_SEGMENT|1288,1293|false|false|false|C0039070;C4554554|Faint - appearance;Syncope|faint
Finding|Sign or Symptom|SIMPLE_SEGMENT|1288,1293|false|false|false|C0039070;C4554554|Faint - appearance;Syncope|faint
Finding|Sign or Symptom|SIMPLE_SEGMENT|1294,1301|false|false|false|C0043144|Wheezing|wheezes
Finding|Idea or Concept|SIMPLE_SEGMENT|1312,1317|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1318,1325|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1318,1325|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Finding|Finding|SIMPLE_SEGMENT|1318,1325|false|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1327,1332|false|false|false|C0028754|Obesity|obese
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1340,1348|false|false|false|C0005847|Blood Vessel|VASCULAR
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1349,1354|false|false|false|C0016504;C0687080|Foot;Paw|Pedal
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|1349,1361|false|false|false|C0232157|Pedal pulse|Pedal Pulses
Drug|Food|SIMPLE_SEGMENT|1355,1361|false|false|false|C5890763||Pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|1355,1361|false|false|false|C0391850|Physiologic pulse|Pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|1355,1361|false|false|false|C0034107|Pulse taking|Pulses
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1425,1428|false|false|false|C0059387;C0074289|selenocysteine;staphylococcal enterotoxin C|sec
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1425,1428|false|false|false|C0059387;C0074289|selenocysteine;staphylococcal enterotoxin C|sec
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|1425,1428|false|false|false|C0059387;C0074289|selenocysteine;staphylococcal enterotoxin C|sec
Drug|Immunologic Factor|SIMPLE_SEGMENT|1425,1428|false|false|false|C0059387;C0074289|selenocysteine;staphylococcal enterotoxin C|sec
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1438,1441|false|false|false|C0059387;C0074289|selenocysteine;staphylococcal enterotoxin C|sec
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1438,1441|false|false|false|C0059387;C0074289|selenocysteine;staphylococcal enterotoxin C|sec
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|1438,1441|false|false|false|C0059387;C0074289|selenocysteine;staphylococcal enterotoxin C|sec
Drug|Immunologic Factor|SIMPLE_SEGMENT|1438,1441|false|false|false|C0059387;C0074289|selenocysteine;staphylococcal enterotoxin C|sec
Finding|Idea or Concept|SIMPLE_SEGMENT|1446,1455|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Finding|Intellectual Product|SIMPLE_SEGMENT|1446,1455|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Finding|Finding|SIMPLE_SEGMENT|1475,1484|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|1475,1484|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Procedure|Health Care Activity|SIMPLE_SEGMENT|1475,1484|false|false|false|C2229507|sensory exam|Sensation
Finding|Finding|SIMPLE_SEGMENT|1495,1501|false|false|false|C1554187|Gender Status - Intact|Intact
Finding|Functional Concept|SIMPLE_SEGMENT|1506,1512|false|false|false|C0332197|Absent|Absent
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1506,1512|false|false|false|C5237010|Expression Negative|Absent
Finding|Mental Process|SIMPLE_SEGMENT|1532,1546|false|false|false|C0033499|Proprioception|Proprioception
Finding|Finding|SIMPLE_SEGMENT|1551,1557|false|false|false|C1554187|Gender Status - Intact|Intact
Finding|Functional Concept|SIMPLE_SEGMENT|1563,1569|false|false|false|C0332197|Absent|Absent
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1563,1569|false|false|false|C5237010|Expression Negative|Absent
Procedure|Health Care Activity|SIMPLE_SEGMENT|1592,1601|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1602,1606|false|false|false|C0587081|Laboratory test finding|Labs
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1620,1625|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|1620,1625|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|1626,1629|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|1634,1637|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1634,1637|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1634,1637|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1644,1647|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1644,1647|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|1644,1647|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1644,1647|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1653,1656|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1653,1656|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|1664,1667|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1664,1667|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1664,1667|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1664,1667|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|1671,1674|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1671,1674|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|1671,1674|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|1671,1674|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1671,1674|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1681,1685|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1702,1705|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1722,1727|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|1722,1727|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Inorganic Chemical|SIMPLE_SEGMENT|1767,1771|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1767,1771|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1767,1771|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1796,1801|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|1796,1801|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1802,1805|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1802,1805|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|1802,1805|false|false|false|C0001899|Alanine Transaminase|ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|1802,1805|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|1802,1805|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|1802,1805|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1802,1805|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|1809,1812|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1809,1812|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1809,1812|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1809,1812|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|1809,1812|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Finding|Gene or Genome|SIMPLE_SEGMENT|1809,1812|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1828,1833|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|1828,1833|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1858,1863|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|1858,1863|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1865,1870|false|false|false|C0019018|Glycosylated hemoglobin A|HbA1c
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1865,1870|false|false|false|C0019018|Glycosylated hemoglobin A|HbA1c
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1865,1870|false|false|false|C0202054|Glucohemoglobin measurement|HbA1c
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1889,1894|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|1889,1894|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1908,1911|false|false|false|C0023821|High Density Lipoproteins|HDL
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1908,1911|false|false|false|C0023821|High Density Lipoproteins|HDL
Finding|Gene or Genome|SIMPLE_SEGMENT|1908,1911|false|false|false|C3715113|HSD11B1 wt Allele|HDL
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1908,1911|false|false|false|C0392885|High density lipoprotein measurement|HDL
Finding|Intellectual Product|SIMPLE_SEGMENT|1942,1947|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|1948,1956|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1948,1963|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|1948,1963|false|false|false|C0489547|Hospital course|Hospital Course
Finding|Body Substance|SIMPLE_SEGMENT|1969,1976|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1969,1976|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1969,1976|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|SIMPLE_SEGMENT|2017,2023|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Finding|Organism Function|SIMPLE_SEGMENT|2017,2023|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Procedure|Health Care Activity|SIMPLE_SEGMENT|2017,2023|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2017,2023|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2031,2037|false|false|false|C1550316|Tarsal|tarsal
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|2031,2044|false|false|false|C0225150|Structure of tarsal canal|tarsal tunnel
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2031,2052|false|false|false|C0196577|Decompression of tarsal tunnel|tarsal tunnel release
Finding|Functional Concept|SIMPLE_SEGMENT|2045,2052|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|release
Procedure|Health Care Activity|SIMPLE_SEGMENT|2045,2052|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2045,2052|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|release
Finding|Body Substance|SIMPLE_SEGMENT|2059,2066|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|2059,2066|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|2059,2066|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2086,2090|false|false|false|C0671954|CD3EAP protein, human|cast
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2086,2090|false|false|false|C0671954|CD3EAP protein, human|cast
Finding|Body Substance|SIMPLE_SEGMENT|2086,2090|false|false|false|C0302143;C0687709;C1413137;C1539080;C1705948;C1825060;C4284789|CAST gene;Childhood Autism Spectrum Test;Children of Alcoholics Screening Test;ERC2 gene;POLR1G gene;POLR1G wt Allele;cast body substance|cast
Finding|Gene or Genome|SIMPLE_SEGMENT|2086,2090|false|false|false|C0302143;C0687709;C1413137;C1539080;C1705948;C1825060;C4284789|CAST gene;Childhood Autism Spectrum Test;Children of Alcoholics Screening Test;ERC2 gene;POLR1G gene;POLR1G wt Allele;cast body substance|cast
Finding|Intellectual Product|SIMPLE_SEGMENT|2086,2090|false|false|false|C0302143;C0687709;C1413137;C1539080;C1705948;C1825060;C4284789|CAST gene;Childhood Autism Spectrum Test;Children of Alcoholics Screening Test;ERC2 gene;POLR1G gene;POLR1G wt Allele;cast body substance|cast
Finding|Conceptual Entity|SIMPLE_SEGMENT|2124,2128|false|false|false|C0868928;C1706256|Case - situation;Clinical Study Case|case
Finding|Functional Concept|SIMPLE_SEGMENT|2124,2128|false|false|false|C0868928;C1706256|Case - situation;Clinical Study Case|case
Finding|Body Substance|SIMPLE_SEGMENT|2135,2142|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|2135,2142|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|2135,2142|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2158,2167|false|false|false|C0945766||procedure
Event|Occupational Activity|SIMPLE_SEGMENT|2158,2167|false|false|false|C1546467|Act Class - procedure|procedure
Finding|Functional Concept|SIMPLE_SEGMENT|2158,2167|false|false|false|C2700391|Procedure (set of actions)|procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2158,2167|false|false|false|C0184661|Interventional procedure|procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2172,2182|false|false|false|C2926599||anesthesia
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2172,2182|false|false|false|C4049933|Anesthesia substance|anesthesia
Finding|Finding|SIMPLE_SEGMENT|2172,2182|false|false|false|C0278134;C2219802|Absence of sensation|anesthesia
Finding|Sign or Symptom|SIMPLE_SEGMENT|2172,2182|false|false|false|C0278134;C2219802|Absence of sensation|anesthesia
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2172,2182|false|false|false|C0002903;C0002912|Anesthesia procedures;Dental anesthesia|anesthesia
Finding|Finding|SIMPLE_SEGMENT|2183,2187|false|false|false|C5575035|Well (answer to question)|well
Finding|Idea or Concept|SIMPLE_SEGMENT|2196,2204|false|false|false|C0750489|apparent|apparent
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2205,2218|true|false|false|C0802632||complications
Finding|Functional Concept|SIMPLE_SEGMENT|2205,2218|true|false|false|C0009566;C1171258|Complication;complication aspects|complications
Finding|Pathologic Function|SIMPLE_SEGMENT|2205,2218|true|false|false|C0009566;C1171258|Complication;complication aspects|complications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2228,2234|false|false|false|C4255046||report
Finding|Intellectual Product|SIMPLE_SEGMENT|2228,2234|false|false|false|C0684224|Report (document)|report
Procedure|Health Care Activity|SIMPLE_SEGMENT|2228,2234|false|false|false|C0700287|Reporting|report
Finding|Gene or Genome|SIMPLE_SEGMENT|2258,2262|false|false|false|C1420638;C1539127;C1710283|CORO7 gene;TCF21 gene;TCF21 wt Allele|POD1
Drug|Organic Chemical|SIMPLE_SEGMENT|2281,2289|false|false|false|C0700899|Benadryl|benadryl
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2281,2289|false|false|false|C0700899|Benadryl|benadryl
Drug|Organic Chemical|SIMPLE_SEGMENT|2294,2297|false|false|false|C0939812|Ruta graveolens preparation|RUE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2294,2297|false|false|false|C0939812|Ruta graveolens preparation|RUE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2298,2302|false|false|false|C5779629|Eruption of skin (disorder)|rash
Finding|Pathologic Function|SIMPLE_SEGMENT|2298,2302|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|SIMPLE_SEGMENT|2298,2302|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Finding|SIMPLE_SEGMENT|2340,2351|false|false|false|C0020649|Hypotension|hypotension
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2357,2360|false|false|false|C0871470|Systolic Pressure|SBP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2357,2360|false|false|false|C0085805|Androgen Binding Protein|SBP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2357,2360|false|false|false|C0085805|Androgen Binding Protein|SBP
Finding|Gene or Genome|SIMPLE_SEGMENT|2357,2360|false|false|false|C1705296;C3274833|CCHCR1 wt Allele;SHBG wt Allele|SBP
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2357,2360|false|false|false|C1306620|Systolic blood pressure measurement|SBP
Finding|Finding|SIMPLE_SEGMENT|2376,2388|false|false|false|C0231221;C0332151|Asymptomatic (finding);Asymptomatic diagnosis of|asymptomatic
Drug|Food|SIMPLE_SEGMENT|2401,2406|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|vital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2401,2412|false|false|false|C0488614;C0518766|Vital signs|vital signs
Procedure|Health Care Activity|SIMPLE_SEGMENT|2401,2412|false|false|false|C0150404|Taking vital signs|vital signs
Finding|Finding|SIMPLE_SEGMENT|2407,2412|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|2407,2412|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Intellectual Product|SIMPLE_SEGMENT|2413,2419|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Finding|SIMPLE_SEGMENT|2432,2436|false|false|false|C5575035|Well (answer to question)|well
Finding|Finding|SIMPLE_SEGMENT|2437,2448|false|false|false|C2709070|on room air|on room air
Drug|Inorganic Chemical|SIMPLE_SEGMENT|2440,2448|false|false|false|C3846005|Room Air|room air
Drug|Inorganic Chemical|SIMPLE_SEGMENT|2445,2448|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2445,2448|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|SIMPLE_SEGMENT|2445,2448|false|false|false|C0001861;C3536832|Air (substance);air|air
Finding|Finding|SIMPLE_SEGMENT|2445,2448|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|SIMPLE_SEGMENT|2445,2448|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|SIMPLE_SEGMENT|2445,2448|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Finding|SIMPLE_SEGMENT|2511,2520|false|false|false|C0460139|Pressure (finding)|pressures
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|2511,2520|false|false|false|C0033095||pressures
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|2531,2539|false|false|false|C0039155|Systole|systolic
Drug|Organic Chemical|SIMPLE_SEGMENT|2553,2561|false|false|false|C0700899|Benadryl|Benadryl
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2553,2561|false|false|false|C0700899|Benadryl|Benadryl
Finding|Finding|SIMPLE_SEGMENT|2562,2568|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|2562,2568|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|2605,2614|false|false|false|C0027415|Narcotics|narcotics
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2605,2614|false|false|false|C0027415|Narcotics|narcotics
Finding|Finding|SIMPLE_SEGMENT|2623,2630|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|2623,2630|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|2623,2630|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2623,2630|false|false|false|C0543467|Operative Surgical Procedures|surgery
Finding|Body Substance|SIMPLE_SEGMENT|2640,2647|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|2640,2647|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|2640,2647|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2672,2678|false|false|false|C5889824||status
Finding|Idea or Concept|SIMPLE_SEGMENT|2672,2678|false|false|false|C1546481|What subject filter - Status|status
Finding|Body Substance|SIMPLE_SEGMENT|2700,2709|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|2700,2709|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|2700,2709|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|2700,2709|false|false|false|C0030685|Patient Discharge|discharge
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2700,2714|false|false|false|C0184713|Discharge to home|discharge home
Finding|Idea or Concept|SIMPLE_SEGMENT|2710,2714|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|2710,2714|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|2710,2714|false|false|false|C1553498|home health encounter|home
Finding|Body Substance|SIMPLE_SEGMENT|2720,2727|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|2720,2727|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|2720,2727|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2734,2738|false|false|false|C0671954|CD3EAP protein, human|cast
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2734,2738|false|false|false|C0671954|CD3EAP protein, human|cast
Finding|Body Substance|SIMPLE_SEGMENT|2734,2738|false|false|false|C0302143;C0687709;C1413137;C1539080;C1705948;C1825060;C4284789|CAST gene;Childhood Autism Spectrum Test;Children of Alcoholics Screening Test;ERC2 gene;POLR1G gene;POLR1G wt Allele;cast body substance|cast
Finding|Gene or Genome|SIMPLE_SEGMENT|2734,2738|false|false|false|C0302143;C0687709;C1413137;C1539080;C1705948;C1825060;C4284789|CAST gene;Childhood Autism Spectrum Test;Children of Alcoholics Screening Test;ERC2 gene;POLR1G gene;POLR1G wt Allele;cast body substance|cast
Finding|Intellectual Product|SIMPLE_SEGMENT|2734,2738|false|false|false|C0302143;C0687709;C1413137;C1539080;C1705948;C1825060;C4284789|CAST gene;Childhood Autism Spectrum Test;Children of Alcoholics Screening Test;ERC2 gene;POLR1G gene;POLR1G wt Allele;cast body substance|cast
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2768,2771|false|false|false|C1452534|ACE protein, human|ACE
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2768,2771|false|false|false|C1452534|ACE protein, human|ACE
Finding|Gene or Genome|SIMPLE_SEGMENT|2768,2771|false|false|false|C1413931;C4284014|ACE gene;Adverse Childhood Experience questionnaire|ACE
Finding|Intellectual Product|SIMPLE_SEGMENT|2768,2771|false|false|false|C1413931;C4284014|ACE gene;Adverse Childhood Experience questionnaire|ACE
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2768,2771|false|false|false|C0050385;C0108844;C0279078;C1879921|CDE Regimen;CDE protocol;cisplatin, cytarabine, and etoposide chemotherapy protocol;cyclophosphamide/doxorubicin protocol|ACE
Finding|Body Substance|SIMPLE_SEGMENT|2777,2784|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|2777,2784|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|2777,2784|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2802,2814|false|false|false|C3263700||instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|2802,2814|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|instructions
Finding|Body Substance|SIMPLE_SEGMENT|2840,2849|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|2840,2849|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|2840,2849|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|2840,2849|false|false|false|C0030685|Patient Discharge|discharge
Finding|Idea or Concept|SIMPLE_SEGMENT|2933,2937|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2938,2947|false|false|false|C3864998||condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2938,2947|false|false|false|C0012634|Disease|condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|2938,2947|false|false|false|C1705253|Logical Condition|condition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2961,2972|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2961,2972|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|2961,2972|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|2961,2985|false|false|false|C1627937|Medications on admission|Medications on Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|2976,2985|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Organic Chemical|SIMPLE_SEGMENT|3007,3016|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3007,3016|false|false|false|C0001927|albuterol|Albuterol
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3017,3024|false|false|false|C1112870|Aerosol Dose Form|Aerosol
Finding|Gene or Genome|SIMPLE_SEGMENT|3025,3028|false|false|false|C1422467|CIAO3 gene|prn
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3033,3036|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Enzyme|SIMPLE_SEGMENT|3033,3036|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Organic Chemical|SIMPLE_SEGMENT|3033,3036|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3033,3036|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Finding|Gene or Genome|SIMPLE_SEGMENT|3033,3036|false|false|false|C1412553|ARSA gene|ASA
Drug|Organic Chemical|SIMPLE_SEGMENT|3038,3046|false|false|false|C0004147|atenolol|Atenolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3038,3046|false|false|false|C0004147|atenolol|Atenolol
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3052,3059|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Hormone|SIMPLE_SEGMENT|3052,3059|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3052,3059|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|3052,3059|false|false|false|C1337112|INS gene|Insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3052,3059|false|false|false|C0202098|Insulin measurement|Insulin
Drug|Organic Chemical|SIMPLE_SEGMENT|3095,3105|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3095,3105|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|SIMPLE_SEGMENT|3095,3117|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3095,3117|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3124,3134|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3124,3134|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Organic Chemical|SIMPLE_SEGMENT|3139,3148|false|false|false|C0025598|metformin|Metformin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3139,3148|false|false|false|C0025598|metformin|Metformin
Drug|Organic Chemical|SIMPLE_SEGMENT|3150,3160|false|false|false|C0591573|Glucophage|Glucophage
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3150,3160|false|false|false|C0591573|Glucophage|Glucophage
Drug|Organic Chemical|SIMPLE_SEGMENT|3174,3187|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3174,3187|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Organic Chemical|SIMPLE_SEGMENT|3193,3203|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3193,3203|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Organic Chemical|SIMPLE_SEGMENT|3217,3223|false|false|false|C0633084|Plavix|Plavix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3217,3223|false|false|false|C0633084|Plavix|Plavix
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3237,3246|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|3237,3246|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|SIMPLE_SEGMENT|3237,3246|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3237,3246|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3237,3246|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Finding|Physiologic Function|SIMPLE_SEGMENT|3237,3246|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3237,3246|false|false|false|C0202194|Potassium measurement|Potassium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|3248,3256|false|false|false|C0008203;C0596019|Chlorides;chloride ion|chloride
Finding|Physiologic Function|SIMPLE_SEGMENT|3248,3256|false|false|false|C4553021|Chloride metabolic function|chloride
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3248,3256|false|false|false|C0201952|Chloride measurement|chloride
Drug|Organic Chemical|SIMPLE_SEGMENT|3266,3277|false|false|false|C0074554|simvastatin|Simvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3266,3277|false|false|false|C0074554|simvastatin|Simvastatin
Finding|Body Substance|SIMPLE_SEGMENT|3286,3295|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|3286,3295|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|3286,3295|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|3286,3295|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|3286,3307|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3296,3307|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3296,3307|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|3296,3307|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|3312,3321|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3312,3321|false|false|false|C0001927|albuterol|Albuterol
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3339,3346|false|false|false|C1112870|Aerosol Dose Form|Aerosol
Finding|Functional Concept|SIMPLE_SEGMENT|3362,3372|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Organism Function|SIMPLE_SEGMENT|3362,3372|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Sign or Symptom|SIMPLE_SEGMENT|3408,3414|false|false|false|C0043144|Wheezing|wheeze
Drug|Organic Chemical|SIMPLE_SEGMENT|3421,3428|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3421,3428|false|false|false|C0004057|aspirin|Aspirin
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3436,3442|false|false|false|C0039225|Tablet Dosage Form|Tablet
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3444,3451|false|false|false|C1545665|Views delayed|Delayed
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3444,3459|false|false|false|C1707664|Delayed Release Dosage Form|Delayed Release
Finding|Functional Concept|SIMPLE_SEGMENT|3452,3459|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|3452,3459|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3452,3459|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3481,3487|false|false|false|C0039225|Tablet Dosage Form|Tablet
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3489,3496|false|false|false|C1545665|Views delayed|Delayed
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3489,3504|false|false|false|C1707664|Delayed Release Dosage Form|Delayed Release
Finding|Functional Concept|SIMPLE_SEGMENT|3497,3504|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|3497,3504|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3497,3504|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|SIMPLE_SEGMENT|3535,3543|false|false|false|C0004147|atenolol|Atenolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3535,3543|false|false|false|C0004147|atenolol|Atenolol
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3550,3556|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3570,3576|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Organic Chemical|SIMPLE_SEGMENT|3600,3610|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3600,3610|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|SIMPLE_SEGMENT|3600,3622|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3600,3622|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3629,3635|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Functional Concept|SIMPLE_SEGMENT|3646,3653|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|3646,3653|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3646,3653|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3674,3680|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Functional Concept|SIMPLE_SEGMENT|3691,3698|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|3691,3698|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3691,3698|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3728,3738|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3728,3738|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3745,3751|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3765,3771|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Organic Chemical|SIMPLE_SEGMENT|3796,3805|false|false|false|C0025598|metformin|Metformin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3796,3805|false|false|false|C0025598|metformin|Metformin
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3813,3819|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3833,3839|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Finding|SIMPLE_SEGMENT|3848,3855|false|false|false|C4035626|3 times|3 times
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3850,3855|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|SIMPLE_SEGMENT|3859,3862|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|3859,3862|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|SIMPLE_SEGMENT|3870,3883|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3870,3883|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3891,3897|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3891,3909|false|false|false|C0991582|Sublingual Tablet|Tablet, Sublingual
Finding|Finding|SIMPLE_SEGMENT|3899,3909|false|false|false|C0001565;C4521982|Sublingual (intended site);Sublingual Route of Administration|Sublingual
Finding|Functional Concept|SIMPLE_SEGMENT|3899,3909|false|false|false|C0001565;C4521982|Sublingual (intended site);Sublingual Route of Administration|Sublingual
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3910,3913|false|false|false|C0262329|Short insular gyrus|Sig
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3910,3913|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Immunologic Factor|SIMPLE_SEGMENT|3910,3913|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Finding|Receptor|SIMPLE_SEGMENT|3910,3913|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3923,3929|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Finding|SIMPLE_SEGMENT|3932,3942|false|false|false|C0001565;C4521982|Sublingual (intended site);Sublingual Route of Administration|Sublingual
Finding|Functional Concept|SIMPLE_SEGMENT|3932,3942|false|false|false|C0001565;C4521982|Sublingual (intended site);Sublingual Route of Administration|Sublingual
Finding|Finding|SIMPLE_SEGMENT|3943,3953|false|false|false|C0001565;C4521982|Sublingual (intended site);Sublingual Route of Administration|Sublingual
Finding|Functional Concept|SIMPLE_SEGMENT|3943,3953|false|false|false|C0001565;C4521982|Sublingual (intended site);Sublingual Route of Administration|Sublingual
Finding|Gene or Genome|SIMPLE_SEGMENT|3954,3957|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|SIMPLE_SEGMENT|3976,3986|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3976,3986|false|false|false|C0028978|omeprazole|Omeprazole
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3993,4000|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|3993,4000|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3993,4000|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4002,4009|false|false|false|C1545665|Views delayed|Delayed
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4002,4017|false|false|false|C1707664|Delayed Release Dosage Form|Delayed Release
Finding|Functional Concept|SIMPLE_SEGMENT|4010,4017|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|4010,4017|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4010,4017|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4038,4045|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|4038,4045|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4038,4045|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4047,4054|false|false|false|C1545665|Views delayed|Delayed
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4047,4062|false|false|false|C1707664|Delayed Release Dosage Form|Delayed Release
Finding|Functional Concept|SIMPLE_SEGMENT|4055,4062|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|4055,4062|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4055,4062|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|SIMPLE_SEGMENT|4092,4103|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4092,4103|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4110,4116|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4130,4136|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4162,4171|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4162,4171|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|SIMPLE_SEGMENT|4162,4171|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4162,4171|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4162,4171|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Finding|Physiologic Function|SIMPLE_SEGMENT|4162,4171|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4162,4171|false|false|false|C0202194|Potassium measurement|Potassium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4162,4180|false|false|false|C0032825|potassium chloride|Potassium Chloride
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4162,4180|false|false|false|C0032825|potassium chloride|Potassium Chloride
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4172,4180|false|false|false|C0008203;C0596019|Chlorides;chloride ion|Chloride
Finding|Physiologic Function|SIMPLE_SEGMENT|4172,4180|false|false|false|C4553021|Chloride metabolic function|Chloride
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4172,4180|false|false|false|C0201952|Chloride measurement|Chloride
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4188,4191|false|false|false|C0039225|Tablet Dosage Form|Tab
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4197,4200|false|false|false|C0919436|REL Protein|Rel
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4197,4200|false|false|false|C0919436|REL Protein|Rel
Finding|Gene or Genome|SIMPLE_SEGMENT|4197,4200|false|false|false|C0035018;C1704703;C1705630|Concept Relationship;REL gene;REL wt Allele|Rel
Finding|Idea or Concept|SIMPLE_SEGMENT|4197,4200|false|false|false|C0035018;C1704703;C1705630|Concept Relationship;REL gene;REL wt Allele|Rel
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|4202,4210|false|false|false|C0597177|Particle|Particle
Finding|Gene or Genome|SIMPLE_SEGMENT|4202,4210|false|false|false|C4085054|PARTICL gene|Particle
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4211,4218|false|false|false|C0025611;C0444626;C1378554;C4551577|Crystal - natural material;Crystal Structure;Crystals;methamphetamine|Crystal
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|4211,4218|false|false|false|C0025611;C0444626;C1378554;C4551577|Crystal - natural material;Crystal Structure;Crystals;methamphetamine|Crystal
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|4211,4218|false|false|false|C0025611;C0444626;C1378554;C4551577|Crystal - natural material;Crystal Structure;Crystals;methamphetamine|Crystal
Drug|Organic Chemical|SIMPLE_SEGMENT|4211,4218|false|false|false|C0025611;C0444626;C1378554;C4551577|Crystal - natural material;Crystal Structure;Crystals;methamphetamine|Crystal
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4211,4218|false|false|false|C0025611;C0444626;C1378554;C4551577|Crystal - natural material;Crystal Structure;Crystals;methamphetamine|Crystal
Finding|Body Substance|SIMPLE_SEGMENT|4211,4218|false|false|false|C0427896|Crystal - human material|Crystal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4233,4236|false|false|false|C0039225|Tablet Dosage Form|Tab
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4242,4245|false|false|false|C0919436|REL Protein|Rel
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4242,4245|false|false|false|C0919436|REL Protein|Rel
Finding|Gene or Genome|SIMPLE_SEGMENT|4242,4245|false|false|false|C0035018;C1704703;C1705630|Concept Relationship;REL gene;REL wt Allele|Rel
Finding|Idea or Concept|SIMPLE_SEGMENT|4242,4245|false|false|false|C0035018;C1704703;C1705630|Concept Relationship;REL gene;REL wt Allele|Rel
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|4247,4255|false|false|false|C0597177|Particle|Particle
Finding|Gene or Genome|SIMPLE_SEGMENT|4247,4255|false|false|false|C4085054|PARTICL gene|Particle
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4256,4263|false|false|false|C0025611;C0444626;C1378554;C4551577|Crystal - natural material;Crystal Structure;Crystals;methamphetamine|Crystal
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|4256,4263|false|false|false|C0025611;C0444626;C1378554;C4551577|Crystal - natural material;Crystal Structure;Crystals;methamphetamine|Crystal
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|4256,4263|false|false|false|C0025611;C0444626;C1378554;C4551577|Crystal - natural material;Crystal Structure;Crystals;methamphetamine|Crystal
Drug|Organic Chemical|SIMPLE_SEGMENT|4256,4263|false|false|false|C0025611;C0444626;C1378554;C4551577|Crystal - natural material;Crystal Structure;Crystals;methamphetamine|Crystal
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4256,4263|false|false|false|C0025611;C0444626;C1378554;C4551577|Crystal - natural material;Crystal Structure;Crystals;methamphetamine|Crystal
Finding|Body Substance|SIMPLE_SEGMENT|4256,4263|false|false|false|C0427896|Crystal - human material|Crystal
Drug|Organic Chemical|SIMPLE_SEGMENT|4288,4299|false|false|false|C0074554|simvastatin|Simvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4288,4299|false|false|false|C0074554|simvastatin|Simvastatin
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4306,4312|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4326,4332|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Organic Chemical|SIMPLE_SEGMENT|4358,4369|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4358,4369|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4358,4380|false|false|false|C0939232|fluticasone / salmeterol|Fluticasone-Salmeterol
Drug|Organic Chemical|SIMPLE_SEGMENT|4370,4380|false|false|false|C0073992|salmeterol|Salmeterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4370,4380|false|false|false|C0073992|salmeterol|Salmeterol
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4397,4401|false|false|false|C1556138|Disc - Body Part|Disk
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4397,4401|false|false|false|C0993608|Disk Drug Form|Disk
Finding|Functional Concept|SIMPLE_SEGMENT|4407,4413|false|false|false|C1550509|Participation Type - device|Device
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4414,4417|false|false|false|C0262329|Short insular gyrus|Sig
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4414,4417|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Immunologic Factor|SIMPLE_SEGMENT|4414,4417|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Finding|Receptor|SIMPLE_SEGMENT|4414,4417|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4428,4432|false|false|false|C1556138|Disc - Body Part|Disk
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4428,4432|false|false|false|C0993608|Disk Drug Form|Disk
Finding|Functional Concept|SIMPLE_SEGMENT|4438,4444|false|false|false|C1550509|Participation Type - device|Device
Finding|Functional Concept|SIMPLE_SEGMENT|4445,4455|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Organism Function|SIMPLE_SEGMENT|4445,4455|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|4456,4459|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4456,4459|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4456,4459|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|4456,4459|false|false|false|C1332410|BID gene|BID
Finding|Finding|SIMPLE_SEGMENT|4461,4468|false|false|false|C4035627|2 times|2 times
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4463,4468|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|SIMPLE_SEGMENT|4471,4474|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|4471,4474|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4483,4490|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Hormone|SIMPLE_SEGMENT|4483,4490|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4483,4490|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|4483,4490|false|false|false|C1337112|INS gene|Insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4483,4490|false|false|false|C0202098|Insulin measurement|Insulin
Drug|Organic Chemical|SIMPLE_SEGMENT|4533,4542|false|false|false|C0701017|Compazine|Compazine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4533,4542|false|false|false|C0701017|Compazine|Compazine
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4549,4555|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4569,4575|false|false|false|C0039225|Tablet Dosage Form|Tablet
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4614,4620|false|false|false|C4255480||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|4614,4620|false|false|false|C0027497|Nausea|nausea
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4631,4637|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|SIMPLE_SEGMENT|4642,4649|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|4658,4667|false|false|false|C0030049|oxycodone|Oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4658,4667|false|false|false|C0030049|oxycodone|Oxycodone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4658,4667|false|false|false|C0524222|Oxycodone measurement|Oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4658,4681|false|false|false|C0717368|acetaminophen / oxycodone|Oxycodone-Acetaminophen
Drug|Organic Chemical|SIMPLE_SEGMENT|4668,4681|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4668,4681|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4668,4681|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4689,4695|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4705,4712|false|false|false|C0039225|Tablet Dosage Form|Tablets
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4751,4755|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|4751,4755|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|4751,4755|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4766,4772|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|SIMPLE_SEGMENT|4777,4784|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|4793,4802|false|false|false|C0030049|oxycodone|Oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4793,4802|false|false|false|C0030049|oxycodone|Oxycodone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4793,4802|false|false|false|C0524222|Oxycodone measurement|Oxycodone
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4809,4815|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Functional Concept|SIMPLE_SEGMENT|4826,4833|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|4826,4833|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4826,4833|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4850,4856|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Functional Concept|SIMPLE_SEGMENT|4867,4874|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|4867,4874|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4867,4874|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4878,4881|false|false|false|C0751781|Dentatorubral-Pallidoluysian Atrophy|hrs
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4878,4881|false|false|false|C1568891|HGS protein, human|hrs
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4878,4881|false|false|false|C1568891|HGS protein, human|hrs
Finding|Gene or Genome|SIMPLE_SEGMENT|4878,4881|false|false|false|C1366514;C1415473;C1419996;C1708271;C5575450;C5780798|ATN1 wt Allele;HARS1 gene;HARS1 wt Allele;HGS gene;HGS wt Allele;SRSF5 gene|hrs
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4917,4923|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Functional Concept|SIMPLE_SEGMENT|4934,4941|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|4934,4941|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4934,4941|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Finding|Idea or Concept|SIMPLE_SEGMENT|4952,4959|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|4968,4976|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4968,4976|false|false|false|C1692318|docusate|Docusate
Drug|Organic Chemical|SIMPLE_SEGMENT|4968,4983|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4968,4983|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4977,4983|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4977,4983|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4977,4983|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|4977,4983|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4977,4983|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4991,4997|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5011,5017|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|SIMPLE_SEGMENT|5030,5033|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|5030,5033|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5044,5050|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|SIMPLE_SEGMENT|5055,5062|false|false|false|C0807726|refill|Refills
Finding|Body Substance|SIMPLE_SEGMENT|5070,5079|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|5070,5079|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|5070,5079|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|5070,5079|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5070,5091|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|5070,5091|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5080,5091|false|false|false|C2926604||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|5080,5091|false|false|false|C0184758|Patient disposition|Disposition
Finding|Idea or Concept|SIMPLE_SEGMENT|5093,5097|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|5093,5097|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|5093,5097|false|false|false|C1553498|home health encounter|Home
Finding|Body Substance|SIMPLE_SEGMENT|5100,5109|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|5100,5109|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|5100,5109|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|5100,5109|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|5100,5119|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5110,5119|false|false|false|C0945731||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|5110,5119|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|5110,5119|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5110,5119|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|5121,5125|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5126,5135|false|false|false|C0751438|Posterior pituitary disease|posterior
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5126,5144|false|false|false|C0224463|Tibialis posterior muscle structure|posterior tibialis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5136,5144|false|false|false|C1710422|Tibialis Muscle|tibialis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5136,5155|false|false|false|C0158321|Tibialis tendinitis|tibialis tendonitis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5145,5155|false|false|false|C0039503|Tendinitis|tendonitis
Finding|Functional Concept|SIMPLE_SEGMENT|5156,5160|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5161,5167|false|false|false|C1550316|Tarsal|tarsal
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5161,5174|false|false|false|C0225150|Structure of tarsal canal|tarsal tunnel
Finding|Body Substance|SIMPLE_SEGMENT|5178,5187|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|5178,5187|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|5178,5187|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|5178,5187|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5188,5197|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5188,5197|false|false|false|C0012634|Disease|Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|5188,5197|false|false|false|C1705253|Logical Condition|Condition
Finding|Idea or Concept|SIMPLE_SEGMENT|5199,5203|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|Good
Finding|Body Substance|SIMPLE_SEGMENT|5207,5216|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|5207,5216|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|5207,5216|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|5207,5216|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5207,5229|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|5207,5229|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|5207,5229|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5217,5229|false|false|false|C3263700||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|5217,5229|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Finding|Conceptual Entity|SIMPLE_SEGMENT|5249,5262|false|false|false|C4724283|Pre-admission Encounter|pre-admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5263,5274|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5263,5274|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|SIMPLE_SEGMENT|5263,5274|false|false|false|C4284232|Medications|medications
Finding|Finding|SIMPLE_SEGMENT|5292,5295|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|5292,5295|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5297,5310|false|false|false|C2741652||prescriptions
Procedure|Health Care Activity|SIMPLE_SEGMENT|5297,5310|false|false|false|C0033080|Prescription (procedure)|prescriptions
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5349,5357|false|false|false|C1705365|Dressing Dosage Form|dressing
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|5349,5357|false|false|false|C0518459;C1305428|Ability to dress|dressing
Finding|Finding|SIMPLE_SEGMENT|5349,5357|false|false|false|C0518459;C1305428|Ability to dress|dressing
Procedure|Health Care Activity|SIMPLE_SEGMENT|5349,5357|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5349,5357|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5358,5362|false|false|false|C0671954|CD3EAP protein, human|cast
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5358,5362|false|false|false|C0671954|CD3EAP protein, human|cast
Finding|Body Substance|SIMPLE_SEGMENT|5358,5362|false|false|false|C0302143;C0687709;C1413137;C1539080;C1705948;C1825060;C4284789|CAST gene;Childhood Autism Spectrum Test;Children of Alcoholics Screening Test;ERC2 gene;POLR1G gene;POLR1G wt Allele;cast body substance|cast
Finding|Gene or Genome|SIMPLE_SEGMENT|5358,5362|false|false|false|C0302143;C0687709;C1413137;C1539080;C1705948;C1825060;C4284789|CAST gene;Childhood Autism Spectrum Test;Children of Alcoholics Screening Test;ERC2 gene;POLR1G gene;POLR1G wt Allele;cast body substance|cast
Finding|Intellectual Product|SIMPLE_SEGMENT|5358,5362|false|false|false|C0302143;C0687709;C1413137;C1539080;C1705948;C1825060;C4284789|CAST gene;Childhood Autism Spectrum Test;Children of Alcoholics Screening Test;ERC2 gene;POLR1G gene;POLR1G wt Allele;cast body substance|cast
Event|Activity|SIMPLE_SEGMENT|5363,5368|false|false|false|C1947930|Cleaning (activity)|clean
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5384,5389|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5415,5423|true|false|false|C1705365|Dressing Dosage Form|dressing
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|5415,5423|true|false|false|C0518459;C1305428|Ability to dress|dressing
Finding|Finding|SIMPLE_SEGMENT|5415,5423|true|false|false|C0518459;C1305428|Ability to dress|dressing
Procedure|Health Care Activity|SIMPLE_SEGMENT|5415,5423|true|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5415,5423|true|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Finding|Functional Concept|SIMPLE_SEGMENT|5424,5431|false|false|false|C0392747|Changing|changes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5457,5463|false|false|false|C0944911||WEIGHT
Finding|Finding|SIMPLE_SEGMENT|5457,5463|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|WEIGHT
Finding|Sign or Symptom|SIMPLE_SEGMENT|5457,5463|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|WEIGHT
Procedure|Health Care Activity|SIMPLE_SEGMENT|5457,5463|false|false|false|C1305866|Weighing patient|WEIGHT
Finding|Functional Concept|SIMPLE_SEGMENT|5480,5484|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5480,5489|false|false|false|C0230461|Structure of left foot|left foot
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5485,5489|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|5485,5489|false|false|false|C0555980|Foot problem|foot
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5495,5499|false|false|false|C0671954|CD3EAP protein, human|cast
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5495,5499|false|false|false|C0671954|CD3EAP protein, human|cast
Finding|Body Substance|SIMPLE_SEGMENT|5495,5499|false|false|false|C0302143;C0687709;C1413137;C1539080;C1705948;C1825060;C4284789|CAST gene;Childhood Autism Spectrum Test;Children of Alcoholics Screening Test;ERC2 gene;POLR1G gene;POLR1G wt Allele;cast body substance|cast
Finding|Gene or Genome|SIMPLE_SEGMENT|5495,5499|false|false|false|C0302143;C0687709;C1413137;C1539080;C1705948;C1825060;C4284789|CAST gene;Childhood Autism Spectrum Test;Children of Alcoholics Screening Test;ERC2 gene;POLR1G gene;POLR1G wt Allele;cast body substance|cast
Finding|Intellectual Product|SIMPLE_SEGMENT|5495,5499|false|false|false|C0302143;C0687709;C1413137;C1539080;C1705948;C1825060;C4284789|CAST gene;Childhood Autism Spectrum Test;Children of Alcoholics Screening Test;ERC2 gene;POLR1G gene;POLR1G wt Allele;cast body substance|cast
Finding|Finding|SIMPLE_SEGMENT|5522,5532|false|false|false|C2135586;C4321408|Wheelchair Usually Used;has wheelchair at home (history)|wheelchair
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5540,5545|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Functional Concept|SIMPLE_SEGMENT|5558,5562|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5564,5568|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|5564,5568|false|false|false|C0555980|Foot problem|foot
Finding|Finding|SIMPLE_SEGMENT|5589,5597|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|5589,5597|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Intellectual Product|SIMPLE_SEGMENT|5611,5617|false|false|false|C2348314|Doctor - Title|doctor
Finding|Functional Concept|SIMPLE_SEGMENT|5642,5650|false|false|false|C0442805|Increase|increase
Finding|Functional Concept|SIMPLE_SEGMENT|5654,5658|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5654,5663|false|false|false|C0230461|Structure of left foot|left foot
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5659,5663|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|5659,5663|false|false|false|C0555980|Foot problem|foot
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5665,5672|false|false|false|C0041834|Erythema|redness
Finding|Finding|SIMPLE_SEGMENT|5665,5672|false|false|false|C0332575|Redness|redness
Finding|Finding|SIMPLE_SEGMENT|5674,5682|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|5674,5682|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Finding|SIMPLE_SEGMENT|5686,5703|false|false|false|C0517630|Purulent drainage|purulent drainage
Finding|Body Substance|SIMPLE_SEGMENT|5695,5703|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|SIMPLE_SEGMENT|5695,5703|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5695,5703|false|false|false|C0013103|Drainage procedure|drainage
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|5714,5719|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Finding|Body Substance|SIMPLE_SEGMENT|5714,5719|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|SIMPLE_SEGMENT|5714,5719|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|SIMPLE_SEGMENT|5714,5719|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5730,5736|false|false|false|C4255480||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|5730,5736|false|false|false|C0027497|Nausea|nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|5738,5746|false|false|false|C0042963|Vomiting|vomiting
Finding|Sign or Symptom|SIMPLE_SEGMENT|5748,5754|false|false|false|C0015967|Fever|fevers
Finding|Sign or Symptom|SIMPLE_SEGMENT|5775,5781|false|false|false|C0085593|Chills|chills
Finding|Body Substance|SIMPLE_SEGMENT|5790,5796|false|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Finding|Finding|SIMPLE_SEGMENT|5790,5796|false|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Finding|Idea or Concept|SIMPLE_SEGMENT|5804,5813|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Finding|Functional Concept|SIMPLE_SEGMENT|5814,5822|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|5814,5822|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Procedure|Health Care Activity|SIMPLE_SEGMENT|5826,5834|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5835,5847|false|false|false|C3263700||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|5835,5847|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

