 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|46,55|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|46,55|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|46,60|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|80,89|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|80,89|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|80,94|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|136,139|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|147,154|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|147,154|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|SIMPLE_SEGMENT|156,168|false|false|false|||NEUROSURGERY
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|156,168|false|false|false|C0524850|Neurosurgical Procedures|NEUROSURGERY
Disorder|Injury or Poisoning|Allergies|183,194|false|false|false|C0161486;C2876539|Poisoning by penicillin;Poisoning by, adverse effect of and underdosing of penicillins|Penicillins
Drug|Antibiotic|Allergies|183,194|false|false|false|C0030842|penicillins|Penicillins
Drug|Organic Chemical|Allergies|183,194|false|false|false|C0030842|penicillins|Penicillins
Event|Event|Allergies|183,194|false|false|false|||Penicillins
Finding|Pathologic Function|Allergies|183,194|false|false|false|C0413443|Adverse reaction to penicillins|Penicillins
Drug|Organic Chemical|Allergies|197,202|false|false|false|C0376414|Paxil|Paxil
Drug|Pharmacologic Substance|Allergies|197,202|false|false|false|C0376414|Paxil|Paxil
Drug|Organic Chemical|Allergies|205,215|false|false|false|C0085934|Wellbutrin|Wellbutrin
Drug|Pharmacologic Substance|Allergies|205,215|false|false|false|C0085934|Wellbutrin|Wellbutrin
Event|Event|Allergies|218,227|false|false|false|||Attending
Finding|Functional Concept|Allergies|218,227|false|false|false|C1999232|Attending (action)|Attending
Event|Event|Chief Complaint|261,269|false|false|false|||hardware
Finding|Classification|Chief Complaint|272,277|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|278,286|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|278,286|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|290,308|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|299,308|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|299,308|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|299,308|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|299,308|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|299,308|false|false|false|C0184661|Interventional procedure|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|318,334|false|false|false|C5453054|Hardware Removal|hardware removal
Event|Activity|Chief Complaint|327,334|false|false|false|C1883720|Removing (action)|removal
Event|Event|Chief Complaint|327,334|false|false|false|||removal
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|327,334|false|false|false|C0015252;C0185115;C0728940|Excision;Extraction;removal technique|removal
Finding|Idea or Concept|History of Present Illness|380,384|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|History of Present Illness|380,384|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|History of Present Illness|385,388|false|false|false|||old
Finding|Finding|History of Present Illness|404,417|false|false|false|C0455610|History of surgery|prior surgery
Event|Event|History of Present Illness|410,417|false|false|false|||surgery
Finding|Finding|History of Present Illness|410,417|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|History of Present Illness|410,417|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|History of Present Illness|410,417|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|410,417|false|false|false|C0543467|Operative Surgical Procedures|surgery
Finding|Finding|History of Present Illness|424,432|false|false|false|C0332149|Possible|possible
Finding|Functional Concept|History of Present Illness|434,439|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Disorder|Neoplastic Process|History of Present Illness|449,471|false|false|false|C0334579|Anaplastic astrocytoma|anaplastic astrocytoma
Disorder|Neoplastic Process|History of Present Illness|460,471|false|false|false|C0004114|Astrocytoma|astrocytoma
Event|Event|History of Present Illness|460,471|false|false|false|||astrocytoma
Event|Event|History of Present Illness|477,487|false|false|false|||craniotomy
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|477,487|false|false|false|C0010280|Craniotomy|craniotomy
Event|Event|History of Present Illness|492,501|false|false|false|||resection
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|492,501|false|false|false|C0015252;C0728940|Excision;removal technique|resection
Finding|Functional Concept|History of Present Illness|540,548|false|false|false|C1314939|Involvement with|involved
Event|Event|History of Present Illness|549,554|false|false|false|||field
Finding|Conceptual Entity|History of Present Illness|549,554|false|false|false|C1521738;C2346620;C2349184|Field;Force Field;Knowledge Field|field
Procedure|Health Care Activity|History of Present Illness|549,554|false|false|false|C1553496|field - patient encounter|field
Event|Event|History of Present Illness|556,567|false|false|false|||irradiation
Phenomenon|Natural Phenomenon or Process|History of Present Illness|556,567|false|false|false|C0851346;C1282930|Irradiation (physical force);Radiation|irradiation
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|556,567|false|false|false|C1522449|Radiation therapy (procedure)|irradiation
Event|Event|History of Present Illness|595,601|false|false|false|||cycles
Drug|Organic Chemical|History of Present Illness|606,613|false|false|false|C0876179|Temodar|Temodar
Drug|Pharmacologic Substance|History of Present Illness|606,613|false|false|false|C0876179|Temodar|Temodar
Event|Event|History of Present Illness|614,619|false|false|false|||ended
Finding|Functional Concept|History of Present Illness|630,636|false|false|false|C1522484;C1561503;C1705190|Precision - second;Second Suffix;metastatic qualifier|second
Finding|Idea or Concept|History of Present Illness|630,636|false|false|false|C1522484;C1561503;C1705190|Precision - second;Second Suffix;metastatic qualifier|second
Finding|Intellectual Product|History of Present Illness|630,636|false|false|false|C1522484;C1561503;C1705190|Precision - second;Second Suffix;metastatic qualifier|second
Event|Event|History of Present Illness|637,647|false|false|false|||craniotomy
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|637,647|false|false|false|C0010280|Craniotomy|craniotomy
Disorder|Neoplastic Process|History of Present Illness|652,657|false|false|false|C0027651|Neoplasms|tumor
Finding|Finding|History of Present Illness|652,657|false|false|false|C1578706;C3273930|Tumor Mass|tumor
Finding|Intellectual Product|History of Present Illness|652,657|false|false|false|C1578706;C3273930|Tumor Mass|tumor
Disorder|Neoplastic Process|History of Present Illness|652,668|false|false|false|C0521158|Recurrent tumor|tumor recurrence
Disorder|Neoplastic Process|History of Present Illness|658,668|false|false|false|C1458156|Recurrent Malignant Neoplasm|recurrence
Event|Event|History of Present Illness|658,668|false|false|false|||recurrence
Finding|Pathologic Function|History of Present Illness|658,668|false|false|false|C2825055|Recurrence (disease attribute)|recurrence
Phenomenon|Phenomenon or Process|History of Present Illness|658,668|false|false|false|C0034897|Recurrence|recurrence
Anatomy|Body Location or Region|History of Present Illness|700,703|false|false|false|C5239890|area PCV|PCV
Disorder|Virus|History of Present Illness|700,703|false|false|false|C0206411|Porcine circovirus|PCV
Drug|Nucleic Acid, Nucleoside, or Nucleotide|History of Present Illness|700,703|false|false|false|C0164815|penciclovir|PCV
Drug|Pharmacologic Substance|History of Present Illness|700,703|false|false|false|C0164815|penciclovir|PCV
Event|Event|History of Present Illness|700,703|false|false|false|||PCV
Procedure|Laboratory Procedure|History of Present Illness|700,703|false|false|false|C0018935;C0070167;C1882252|Hematocrit Measurement;Procarbazine-Lomustine-Vincristine (PCV) Regimen;lomustine/procarbazine/vincristine|PCV
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|700,703|false|false|false|C0018935;C0070167;C1882252|Hematocrit Measurement;Procarbazine-Lomustine-Vincristine (PCV) Regimen;lomustine/procarbazine/vincristine|PCV
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|704,708|false|false|false|C0376161|Comb (body structure)|comb
Drug|Organic Chemical|History of Present Illness|704,708|false|false|false|C0278789|Combid|comb
Drug|Pharmacologic Substance|History of Present Illness|704,708|false|false|false|C0278789|Combid|comb
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|704,708|false|false|false|C0279325;C0280054|bleomycin/cyclophosphamide/methotrexate/vincristine protocol;bleomycin/cyclophosphamide/semustine/vincristine protocol|comb
Event|Event|History of Present Illness|709,714|false|false|false|||chemo
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|709,714|false|false|false|C0392920;C3665472|Chemotherapy;Chemotherapy Regimen|chemo
Event|Event|History of Present Illness|741,750|false|false|false|||presented
Event|Event|History of Present Illness|764,772|false|false|false|||hardware
Event|Event|History of Present Illness|780,786|false|false|false|||office
Finding|Idea or Concept|History of Present Illness|780,786|false|false|false|C1549636|Address type - Office|office
Event|Event|History of Present Illness|796,802|false|false|false|||needed
Event|Event|History of Present Illness|803,812|false|false|false|||admission
Procedure|Health Care Activity|History of Present Illness|803,812|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Drug|Chemical Viewed Structurally|History of Present Illness|816,823|false|false|false|C1704241|complex (molecular entity)|complex
Event|Event|History of Present Illness|824,832|false|false|false|||revision
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|824,832|false|false|false|C0558347;C1527075|Revision procedure;Surgical revision|revision
Event|Event|History of Present Illness|855,861|false|false|false|||eroded
Anatomy|Body System|History of Present Illness|874,878|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|History of Present Illness|874,878|false|true|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|History of Present Illness|874,878|false|true|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Finding|Body Substance|History of Present Illness|874,878|false|true|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|History of Present Illness|874,878|false|true|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Drug|Substance|History of Present Illness|880,888|false|false|false|C0032167|Plastics|Plastics
Event|Event|History of Present Illness|880,888|false|false|false|||Plastics
Event|Event|History of Present Illness|895,908|false|false|false|||reconstructed
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|913,918|false|false|false|C0036270|Scalp structure|scalp
Finding|Finding|History of Present Illness|928,932|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|History of Present Illness|928,932|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|History of Present Illness|928,932|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Body Substance|History of Present Illness|939,946|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|939,946|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|939,946|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|947,955|false|false|false|||presents
Event|Event|History of Present Illness|978,985|false|false|false|||history
Finding|Conceptual Entity|History of Present Illness|978,985|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|978,985|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|978,985|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|978,988|false|false|false|C0262926|Medical History|history of
Event|Event|History of Present Illness|989,997|false|false|false|||pruritus
Finding|Sign or Symptom|History of Present Illness|989,997|false|false|false|C0033774|Pruritus|pruritus
Anatomy|Body Location or Region|History of Present Illness|1017,1021|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1017,1021|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|History of Present Illness|1017,1021|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1017,1021|false|false|false|C0876917|Procedure on head|head
Finding|Idea or Concept|History of Present Illness|1026,1031|false|false|false|C0750546|newly|newly
Event|Event|History of Present Illness|1032,1041|false|false|false|||diagnosed
Event|Event|History of Present Illness|1050,1058|false|false|false|||hardware
Event|Event|History of Present Illness|1065,1072|false|false|false|||reports
Event|Event|History of Present Illness|1098,1102|false|false|false|||look
Anatomy|Body Location or Region|History of Present Illness|1121,1125|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1121,1125|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|History of Present Illness|1121,1125|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1121,1125|false|false|false|C0876917|Procedure on head|head
Finding|Gene or Genome|History of Present Illness|1135,1138|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|History of Present Illness|1144,1147|false|false|false|||saw
Drug|Inorganic Chemical|History of Present Illness|1153,1158|false|false|false|C0025552|Metals|metal
Event|Event|History of Present Illness|1159,1167|false|false|false|||hardware
Finding|Finding|History of Present Illness|1177,1190|false|false|false|C0455610|History of surgery|prior surgery
Event|Event|History of Present Illness|1183,1190|false|false|false|||surgery
Finding|Finding|History of Present Illness|1183,1190|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|History of Present Illness|1183,1190|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|History of Present Illness|1183,1190|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1183,1190|false|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Event|History of Present Illness|1196,1203|false|false|false|||present
Finding|Finding|History of Present Illness|1196,1203|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|History of Present Illness|1196,1203|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Functional Concept|Past Medical History|1229,1234|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Disorder|Neoplastic Process|Past Medical History|1244,1266|false|false|false|C0334579|Anaplastic astrocytoma|anaplastic astrocytoma
Disorder|Neoplastic Process|Past Medical History|1255,1266|false|true|false|C0004114|Astrocytoma|astrocytoma
Event|Event|Past Medical History|1255,1266|false|false|false|||astrocytoma
Event|Event|Past Medical History|1268,1278|false|false|false|||Craniotomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1268,1278|false|false|false|C0010280|Craniotomy|Craniotomy
Event|Event|Past Medical History|1303,1314|false|false|false|||irradiation
Phenomenon|Natural Phenomenon or Process|Past Medical History|1303,1314|false|false|false|C0851346;C1282930|Irradiation (physical force);Radiation|irradiation
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1303,1314|false|false|false|C1522449|Radiation therapy (procedure)|irradiation
Event|Event|Past Medical History|1344,1350|false|false|false|||cycles
Drug|Organic Chemical|Past Medical History|1354,1361|false|false|false|C0876179|Temodar|Temodar
Drug|Pharmacologic Substance|Past Medical History|1354,1361|false|false|false|C0876179|Temodar|Temodar
Event|Event|Past Medical History|1362,1367|false|false|false|||ended
Event|Event|Past Medical History|1374,1384|false|false|false|||craniotomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1374,1384|false|false|false|C0010280|Craniotomy|craniotomy
Disorder|Injury or Poisoning|Past Medical History|1422,1427|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Event|Event|Past Medical History|1422,1427|false|false|false|||wound
Finding|Body Substance|Past Medical History|1422,1427|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|Past Medical History|1422,1427|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|Past Medical History|1422,1427|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Event|Event|Past Medical History|1428,1436|false|false|false|||revision
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1428,1436|false|false|false|C0558347;C1527075|Revision procedure;Surgical revision|revision
Event|Activity|Past Medical History|1441,1448|false|false|false|C1883720|Removing (action)|removal
Event|Event|Past Medical History|1441,1448|false|false|false|||removal
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1441,1448|false|false|false|C0015252;C0185115;C0728940|Excision;Extraction;removal technique|removal
Event|Event|Past Medical History|1474,1482|false|false|false|||hardware
Drug|Organic Chemical|Past Medical History|1484,1492|false|false|false|C0699581|Accutane|Accutane
Drug|Pharmacologic Substance|Past Medical History|1484,1492|false|false|false|C0699581|Accutane|Accutane
Event|Event|Past Medical History|1484,1492|false|false|false|||Accutane
Disorder|Disease or Syndrome|Past Medical History|1514,1521|false|false|false|C0012634|Disease|disease
Event|Event|Past Medical History|1514,1521|false|false|false|||disease
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1536,1550|false|false|false|C0520483|Tubal Ligation|tubal ligation
Event|Event|Past Medical History|1542,1550|false|false|false|||ligation
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1542,1550|false|false|false|C0023690|Ligation|ligation
Event|Event|Past Medical History|1551,1564|false|false|false|||tonsillectomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1551,1564|false|false|false|C0040423|Tonsillectomy|tonsillectomy
Disorder|Disease or Syndrome|Past Medical History|1566,1576|false|false|false|C0006277;C0149514|Acute bronchitis;Bronchitis|bronchitis
Event|Event|Past Medical History|1566,1576|false|false|false|||bronchitis
Disorder|Mental or Behavioral Dysfunction|Past Medical History|1578,1588|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|depression
Event|Event|Past Medical History|1578,1588|false|false|false|||depression
Finding|Functional Concept|Past Medical History|1578,1588|false|false|false|C0460137;C1579931|Depression - motion|depression
Finding|Sign or Symptom|Past Medical History|1578,1588|false|false|false|C0460137;C1579931|Depression - motion|depression
Event|Event|Past Medical History|1592,1600|false|false|false|||seizures
Finding|Sign or Symptom|Past Medical History|1592,1600|false|false|false|C0036572|Seizures|seizures
Disorder|Disease or Syndrome|General Exam|1669,1674|false|false|false|C0028754|Obesity|obese
Event|Event|General Exam|1669,1674|false|false|false|||obese
Event|Event|General Exam|1675,1678|false|false|false|||Gen
Finding|Classification|General Exam|1675,1678|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Finding|Gene or Genome|General Exam|1675,1678|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Event|Event|General Exam|1687,1698|false|false|false|||comfortable
Finding|Finding|General Exam|1687,1698|false|false|false|C5546696|Feeling comfortable|comfortable
Disorder|Disease or Syndrome|General Exam|1700,1703|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|1700,1703|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|1700,1703|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|1700,1703|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|1700,1703|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|General Exam|1700,1703|false|false|false|||NAD
Finding|Finding|General Exam|1700,1703|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|General Exam|1705,1710|false|false|false|C1512338|HEENT|HEENT
Event|Event|General Exam|1722,1726|false|false|false|||EOMs
Finding|Functional Concept|General Exam|1722,1726|false|false|false|C0241886|Extraocular|EOMs
Event|Event|General Exam|1728,1734|false|false|false|||intact
Finding|Finding|General Exam|1728,1734|false|false|false|C1554187|Gender Status - Intact|intact
Anatomy|Body Location or Region|General Exam|1735,1739|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|General Exam|1735,1739|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|General Exam|1735,1739|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|General Exam|1741,1747|false|false|false|||Supple
Finding|Functional Concept|General Exam|1741,1747|false|false|false|C0332254|Supple|Supple
Event|Event|General Exam|1752,1755|true|false|false|||LNN
Event|Event|General Exam|1756,1759|true|false|false|||RRR
Event|Event|General Exam|1763,1766|true|false|false|||SOB
Finding|Sign or Symptom|General Exam|1763,1766|true|false|false|C0013404|Dyspnea|SOB
Disorder|Disease or Syndrome|General Exam|1767,1772|true|false|false|C0028754|Obesity|obese
Event|Event|General Exam|1767,1772|true|false|false|||obese
Event|Event|General Exam|1781,1785|false|false|false|||Warm
Finding|Finding|General Exam|1781,1785|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|1781,1785|false|false|false|C0687712|warming process|Warm
Finding|Finding|General Exam|1790,1794|false|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|1795,1803|false|false|false|||perfused
Finding|Mental Process|General Exam|1814,1820|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|General Exam|1814,1827|false|false|false|C0488568;C0488569||Mental status
Finding|Finding|General Exam|1814,1827|false|false|false|C0278060|Mental state|Mental status
Attribute|Clinical Attribute|General Exam|1821,1827|false|false|false|C5889824||status
Event|Event|General Exam|1821,1827|false|false|false|||status
Finding|Idea or Concept|General Exam|1821,1827|false|false|false|C1546481|What subject filter - Status|status
Event|Event|General Exam|1829,1834|false|false|false|||Awake
Attribute|Clinical Attribute|General Exam|1839,1844|false|false|false|C5890168||alert
Drug|Organic Chemical|General Exam|1839,1844|false|false|false|C0718338|Alert brand of caffeine|alert
Drug|Pharmacologic Substance|General Exam|1839,1844|false|false|false|C0718338|Alert brand of caffeine|alert
Event|Event|General Exam|1839,1844|false|false|false|||alert
Finding|Finding|General Exam|1839,1844|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Functional Concept|General Exam|1839,1844|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Intellectual Product|General Exam|1839,1844|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Event|Event|General Exam|1846,1857|false|false|false|||cooperative
Event|Event|General Exam|1863,1867|false|false|false|||exam
Finding|Functional Concept|General Exam|1863,1867|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|General Exam|1863,1867|false|false|false|C0582103|Medical Examination|exam
Event|Event|General Exam|1869,1875|false|false|false|||normal
Event|Event|General Exam|1876,1882|false|false|false|||affect
Finding|Mental Process|General Exam|1876,1882|false|false|false|C0001721|Affect (mental function)|affect
Procedure|Health Care Activity|General Exam|1876,1882|false|false|false|C2237113|assessment of affect|affect
Finding|Gene or Genome|General Exam|1892,1898|false|false|false|C1424587|LITAF gene|simple
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|1899,1908|false|false|false|C0012931|Recombinant DNA|construct
Event|Event|General Exam|1899,1908|false|false|false|||construct
Finding|Idea or Concept|General Exam|1899,1908|false|false|false|C2827421|Construct|construct
Event|Event|General Exam|1910,1921|false|false|false|||Orientation
Finding|Mental Process|General Exam|1910,1921|false|false|false|C0029266|Mental Orientation|Orientation
Event|Event|General Exam|1923,1931|false|false|false|||Oriented
Finding|Finding|General Exam|1923,1931|false|false|false|C1961028|Oriented to place|Oriented
Finding|Finding|General Exam|1923,1941|false|false|false|C1961030|Oriented to person|Oriented to person
Attribute|Clinical Attribute|General Exam|1935,1941|false|false|false|C5890614||person
Event|Event|General Exam|1935,1941|false|false|false|||person
Finding|Intellectual Product|General Exam|1935,1941|false|false|false|C1522390|Person Info|person
Event|Activity|General Exam|1943,1948|false|false|false|C1882509|put - instruction imperative|place
Event|Event|General Exam|1943,1948|false|false|false|||place
Finding|Functional Concept|General Exam|1943,1948|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|General Exam|1943,1948|false|false|false|C1533810||place
Event|Event|General Exam|1960,1966|false|false|false|||Recall
Event|Governmental or Regulatory Activity|General Exam|1960,1966|false|false|false|C1705180|Recall (activity)|Recall
Finding|Mental Process|General Exam|1960,1966|false|false|false|C0034770|Mental Recall|Recall
Event|Event|General Exam|1972,1979|false|false|false|||objects
Procedure|Therapeutic or Preventive Procedure|General Exam|1983,1992|false|false|false|C0886384|5 minutes Office visit|5 minutes
Event|Event|General Exam|1985,1992|false|false|false|||minutes
Attribute|Clinical Attribute|General Exam|1994,2002|false|false|false|C2706915||Language
Event|Event|General Exam|1994,2002|false|false|false|||Language
Finding|Intellectual Product|General Exam|1994,2002|false|false|false|C0033348|Programming Languages|Language
Event|Event|General Exam|2004,2010|false|false|false|||Speech
Finding|Organism Function|General Exam|2004,2010|false|false|false|C0037817|Speech|Speech
Procedure|Diagnostic Procedure|General Exam|2004,2010|false|false|false|C0846595|Speech assessment|Speech
Finding|Idea or Concept|General Exam|2023,2027|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Event|Event|General Exam|2028,2041|false|false|false|||comprehension
Finding|Mental Process|General Exam|2028,2041|false|false|false|C0162340|Comprehension|comprehension
Event|Event|General Exam|2046,2056|false|false|false|||repetition
Finding|Finding|General Exam|2046,2056|false|false|false|C0205341;C2018025|Repeat;speech fluency repetition (physical finding)|repetition
Finding|Functional Concept|General Exam|2046,2056|false|false|false|C0205341;C2018025|Repeat;speech fluency repetition (physical finding)|repetition
Event|Event|General Exam|2058,2064|false|false|false|||Naming
Finding|Mental Process|General Exam|2058,2064|false|false|false|C0233735|Naming (function)|Naming
Event|Event|General Exam|2065,2071|false|false|false|||intact
Finding|Finding|General Exam|2065,2071|false|false|false|C1554187|Gender Status - Intact|intact
Disorder|Mental or Behavioral Dysfunction|General Exam|2076,2086|true|false|false|C0013362|Dysarthria|dysarthria
Event|Event|General Exam|2076,2086|true|false|false|||dysarthria
Event|Event|General Exam|2101,2107|true|false|false|||errors
Anatomy|Body Part, Organ, or Organ Component|General Exam|2110,2117|false|false|false|C0037303|Bone structure of cranium|Cranial
Anatomy|Body Part, Organ, or Organ Component|General Exam|2110,2124|false|false|false|C0010268|Cranial Nerves|Cranial Nerves
Disorder|Neoplastic Process|General Exam|2110,2124|false|false|false|C0004992;C0496937|Benign neoplasm of cranial nerves;Neoplasm of uncertain or unknown behavior of cranial nerves|Cranial Nerves
Anatomy|Body Part, Organ, or Organ Component|General Exam|2118,2124|false|false|false|C0027740|Nerve|Nerves
Event|Event|General Exam|2133,2139|true|false|false|||tested
Anatomy|Body Part, Organ, or Organ Component|General Exam|2144,2150|false|false|false|C0034121|Pupil|Pupils
Event|Event|General Exam|2159,2164|false|false|false|||round
Event|Event|General Exam|2169,2177|false|false|false|||reactive
Procedure|Therapeutic or Preventive Procedure|General Exam|2169,2177|false|false|false|C4722408|Reactive Therapy|reactive
Finding|Finding|General Exam|2169,2186|false|false|false|C4068744|Reactive to light|reactive to light
Drug|Amino Acid, Peptide, or Protein|General Exam|2181,2186|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|General Exam|2181,2186|false|false|false|C1570446|TNFSF14 protein, human|light
Event|Event|General Exam|2181,2186|false|false|false|||light
Finding|Finding|General Exam|2181,2186|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|General Exam|2181,2186|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|General Exam|2181,2186|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|General Exam|2181,2186|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|General Exam|2181,2186|false|false|false|C0031765|Phototherapy|light
Finding|Functional Concept|General Exam|2212,2218|false|false|false|C0234621|Visual|Visual
Event|Event|General Exam|2219,2225|false|false|false|||fields
Event|Event|General Exam|2230,2234|false|false|false|||full
Event|Event|General Exam|2238,2251|false|false|false|||confrontation
Finding|Finding|General Exam|2238,2251|false|false|false|C0518608|Social confrontation skill|confrontation
Procedure|Diagnostic Procedure|General Exam|2238,2251|false|false|false|C0700282;C1444674|Confrontation;Confrontation visual field test|confrontation
Procedure|Therapeutic or Preventive Procedure|General Exam|2238,2251|false|false|false|C0700282;C1444674|Confrontation;Confrontation visual field test|confrontation
Finding|Functional Concept|General Exam|2266,2277|true|false|false|C0241886|Extraocular|Extraocular
Procedure|Diagnostic Procedure|General Exam|2266,2287|true|false|false|C2228439|examination of extraocular movements|Extraocular movements
Event|Event|General Exam|2278,2287|true|false|false|||movements
Finding|Organism Function|General Exam|2278,2287|true|false|false|C0026649|Movement|movements
Event|Event|General Exam|2288,2294|true|false|false|||intact
Finding|Finding|General Exam|2288,2294|true|false|false|C1554187|Gender Status - Intact|intact
Disorder|Disease or Syndrome|General Exam|2315,2324|true|false|false|C0028738|Nystagmus|nystagmus
Event|Event|General Exam|2315,2324|true|false|false|||nystagmus
Anatomy|Body Part, Organ, or Organ Component|General Exam|2329,2332|false|false|false|C2338708;C3496273;C3496274|Lamina VII of gray matter of spinal cord;layer VII (Cajal);lobule VII|VII
Finding|Intellectual Product|General Exam|2329,2332|false|false|false|C0445385|Roman numeral VII|VII
Anatomy|Body Location or Region|General Exam|2334,2340|false|false|false|C0015450|Face|Facial
Event|Event|General Exam|2341,2349|false|false|false|||strength
Finding|Idea or Concept|General Exam|2341,2349|false|false|false|C0808080|Strength (attribute)|strength
Event|Event|General Exam|2354,2363|false|false|false|||sensation
Finding|Finding|General Exam|2354,2363|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|General Exam|2354,2363|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|General Exam|2354,2363|false|false|false|C2229507|sensory exam|sensation
Event|Event|General Exam|2364,2370|false|false|false|||intact
Finding|Finding|General Exam|2364,2370|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|General Exam|2375,2384|false|false|false|||symmetric
Finding|Conceptual Entity|General Exam|2375,2384|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|General Exam|2375,2384|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Anatomy|Body Part, Organ, or Organ Component|General Exam|2386,2390|false|false|false|C0228488;C2327388|Cerebellar pyramis;Lamina VIII of gray matter of spinal cord|VIII
Finding|Gene or Genome|General Exam|2386,2390|false|false|false|C0445599;C1413661|COX8A gene;Roman numeral VIII|VIII
Finding|Intellectual Product|General Exam|2386,2390|false|false|false|C0445599;C1413661|COX8A gene;Roman numeral VIII|VIII
Event|Event|General Exam|2392,2399|false|false|false|||Hearing
Finding|Finding|General Exam|2392,2399|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|Hearing
Finding|Physiologic Function|General Exam|2392,2399|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|Hearing
Event|Event|General Exam|2400,2406|false|false|false|||intact
Finding|Finding|General Exam|2400,2406|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|General Exam|2410,2415|false|false|false|||voice
Finding|Idea or Concept|General Exam|2410,2415|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Intellectual Product|General Exam|2410,2415|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Organism Function|General Exam|2410,2415|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Anatomy|Body Part, Organ, or Organ Component|General Exam|2424,2431|false|false|false|C0700374|Palate|Palatal
Event|Event|General Exam|2432,2441|false|false|false|||elevation
Procedure|Therapeutic or Preventive Procedure|General Exam|2432,2441|false|false|false|C0439775|Elevation procedure|elevation
Event|Event|General Exam|2442,2453|false|false|false|||symmetrical
Finding|Finding|General Exam|2442,2453|false|false|false|C0332516|Symmetrical|symmetrical
Anatomy|Body Part, Organ, or Organ Component|General Exam|2459,2478|false|false|false|C0224153|Structure of sternocleidomastoid muscle|Sternocleidomastoid
Anatomy|Body Part, Organ, or Organ Component|General Exam|2483,2492|false|false|false|C0224361|Structure of trapezius muscle|trapezius
Event|Event|General Exam|2493,2499|false|false|false|||normal
Anatomy|Body Part, Organ, or Organ Component|General Exam|2518,2524|true|false|false|C0040408|Tongue|Tongue
Disorder|Neoplastic Process|General Exam|2518,2524|true|false|false|C0153933|Benign neoplasm of tongue|Tongue
Procedure|Health Care Activity|General Exam|2518,2524|true|false|false|C0872394|Procedure on tongue|Tongue
Finding|Finding|General Exam|2518,2532|true|false|false|C3693372|tongue midline|Tongue midline
Anatomy|Cell Component|General Exam|2525,2532|true|false|false|C1660780|midline cell component|midline
Event|Event|General Exam|2541,2555|true|false|false|||fasciculations
Finding|Sign or Symptom|General Exam|2541,2555|true|false|false|C0015644|Muscular fasciculation|fasciculations
Event|Event|General Exam|2558,2563|false|false|false|||Motor
Finding|Functional Concept|General Exam|2558,2563|false|false|false|C1513492|motor movement|Motor
Drug|Biomedical or Dental Material|General Exam|2572,2576|false|false|false|C0012173;C1337615|Bulk (conceptual);Dietary Fiber|bulk
Drug|Food|General Exam|2572,2576|false|false|false|C0012173;C1337615|Bulk (conceptual);Dietary Fiber|bulk
Event|Event|General Exam|2572,2576|false|false|false|||bulk
Event|Event|General Exam|2581,2585|false|false|false|||tone
Finding|Finding|General Exam|2602,2610|true|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Finding|Idea or Concept|General Exam|2602,2610|true|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Disorder|Disease or Syndrome|General Exam|2602,2620|true|false|false|C0013384|Dyskinetic syndrome|abnormal movements
Finding|Finding|General Exam|2602,2620|true|false|false|C0558189|Abnormal movement|abnormal movements
Event|Event|General Exam|2611,2620|true|false|false|||movements
Finding|Organism Function|General Exam|2611,2620|true|false|false|C0026649|Movement|movements
Event|Event|General Exam|2637,2641|false|false|false|||area
Event|Governmental or Regulatory Activity|General Exam|2637,2641|false|false|false|C1510751|Academic Research Enhancement Awards|area
Event|Event|General Exam|2672,2677|false|false|false|||shows
Event|Event|General Exam|2681,2688|false|false|false|||chronic
Finding|Intellectual Product|General Exam|2681,2688|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|General Exam|2681,2688|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Anatomy|Body System|General Exam|2689,2693|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|General Exam|2689,2693|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|General Exam|2689,2693|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Finding|Body Substance|General Exam|2689,2693|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|General Exam|2689,2693|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Disorder|Disease or Syndrome|General Exam|2694,2700|false|false|false|C1861101|THYROID HORMONE PLASMA MEMBRANE TRANSPORT DEFECT|defect
Event|Event|General Exam|2694,2700|false|false|false|||defect
Finding|Functional Concept|General Exam|2694,2700|false|false|false|C1457869|Defect|defect
Finding|Finding|General Exam|2711,2721|false|false|false|C4722602|Underlying|underlying
Event|Event|General Exam|2722,2729|false|false|false|||harware
Event|Event|General Exam|2734,2740|false|false|false|||eroded
Anatomy|Body System|General Exam|2753,2757|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|General Exam|2753,2757|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|General Exam|2753,2757|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Event|Event|General Exam|2753,2757|false|false|false|||skin
Finding|Body Substance|General Exam|2753,2757|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|General Exam|2753,2757|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Event|Event|General Exam|2759,2768|false|false|false|||Different
Event|Event|General Exam|2783,2791|false|false|false|||repaired
Event|Event|General Exam|2804,2814|false|false|false|||represents
Event|Event|General Exam|2854,2863|true|false|false|||discharge
Finding|Body Substance|General Exam|2854,2863|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|General Exam|2854,2863|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|General Exam|2854,2863|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|General Exam|2854,2863|true|false|false|C0030685|Patient Discharge|discharge
Event|Event|General Exam|2882,2890|true|false|false|||swelling
Finding|Finding|General Exam|2882,2890|true|true|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|General Exam|2882,2890|true|true|false|C0013604;C0038999|Edema;Swelling|swelling
Event|Event|General Exam|2922,2930|false|false|false|||PHYSICAL
Finding|Finding|General Exam|2922,2930|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|General Exam|2922,2930|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|General Exam|2922,2930|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|General Exam|2922,2935|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|General Exam|2922,2935|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Event|Event|General Exam|2931,2935|false|false|false|||EXAM
Finding|Functional Concept|General Exam|2931,2935|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|2931,2935|false|false|false|C0582103|Medical Examination|EXAM
Event|Event|General Exam|2936,2941|false|false|false|||PRIOR
Event|Event|General Exam|2945,2954|false|false|false|||DISCHARGE
Finding|Body Substance|General Exam|2945,2954|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|2945,2954|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|2945,2954|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|2945,2954|false|false|false|C0030685|Patient Discharge|DISCHARGE
Disorder|Disease or Syndrome|General Exam|2964,2969|false|false|false|C0028754|Obesity|obese
Event|Event|General Exam|2964,2969|false|false|false|||obese
Event|Event|General Exam|2970,2973|false|false|false|||Gen
Finding|Classification|General Exam|2970,2973|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Finding|Gene or Genome|General Exam|2970,2973|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Event|Event|General Exam|2982,2993|false|false|false|||comfortable
Finding|Finding|General Exam|2982,2993|false|false|false|C5546696|Feeling comfortable|comfortable
Disorder|Disease or Syndrome|General Exam|2995,2998|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|2995,2998|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|2995,2998|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|2995,2998|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|2995,2998|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|General Exam|2995,2998|false|false|false|||NAD
Finding|Finding|General Exam|2995,2998|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|General Exam|3000,3005|false|false|false|C1512338|HEENT|HEENT
Event|Event|General Exam|3017,3021|false|false|false|||EOMs
Finding|Functional Concept|General Exam|3017,3021|false|false|false|C0241886|Extraocular|EOMs
Event|Event|General Exam|3023,3029|false|false|false|||intact
Finding|Finding|General Exam|3023,3029|false|false|false|C1554187|Gender Status - Intact|intact
Anatomy|Body Location or Region|General Exam|3030,3034|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|General Exam|3030,3034|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|General Exam|3030,3034|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|General Exam|3036,3042|false|false|false|||Supple
Finding|Functional Concept|General Exam|3036,3042|false|false|false|C0332254|Supple|Supple
Anatomy|Body Location or Region|General Exam|3044,3052|false|false|false|C2338258|Cranial incision point|Incision
Disorder|Injury or Poisoning|General Exam|3044,3052|false|false|false|C0332803|Surgical wound|Incision
Event|Event|General Exam|3044,3052|false|false|false|||Incision
Procedure|Therapeutic or Preventive Procedure|General Exam|3044,3052|false|false|false|C0184898|Surgical incisions|Incision
Event|Activity|General Exam|3054,3059|false|false|false|C1947930|Cleaning (activity)|clean
Event|Event|General Exam|3066,3072|false|false|false|||intact
Finding|Finding|General Exam|3066,3072|false|false|false|C1554187|Gender Status - Intact|intact
Disorder|Disease or Syndrome|General Exam|3077,3084|true|false|false|C0041834|Erythema|redness
Event|Event|General Exam|3077,3084|true|false|false|||redness
Finding|Finding|General Exam|3077,3084|true|false|false|C0332575|Redness|redness
Event|Event|General Exam|3086,3094|true|false|false|||swelling
Finding|Finding|General Exam|3086,3094|true|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|General Exam|3086,3094|true|false|false|C0013604;C0038999|Edema;Swelling|swelling
Disorder|Disease or Syndrome|General Exam|3096,3104|true|false|false|C0041834|Erythema|erythema
Event|Event|General Exam|3096,3104|true|false|false|||erythema
Event|Event|General Exam|3109,3118|false|false|false|||discharge
Finding|Body Substance|General Exam|3109,3118|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|General Exam|3109,3118|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|General Exam|3109,3118|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|General Exam|3109,3118|false|false|false|C0030685|Patient Discharge|discharge
Anatomy|Body Space or Junction|General Exam|3120,3127|false|false|false|C0502420|Suture Joint|Sutures
Event|Activity|General Exam|3131,3136|false|false|false|C1882509|put - instruction imperative|place
Event|Event|General Exam|3131,3136|false|false|false|||place
Finding|Functional Concept|General Exam|3131,3136|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|General Exam|3131,3136|false|false|false|C1533810||place
Event|Event|General Exam|3165,3175|false|false|false|||Hematology
Finding|Intellectual Product|General Exam|3165,3175|false|false|false|C1547985|Diagnostic Service Section ID - Hematology|Hematology
Procedure|Laboratory Procedure|General Exam|3165,3175|false|false|false|C0018941;C0200627;C2183233|Hematologic Tests;Hematology procedure;diagnostic service sources hematology (procedure)|Hematology
Drug|Organic Chemical|General Exam|3177,3185|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|COMPLETE
Drug|Pharmacologic Substance|General Exam|3177,3185|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|COMPLETE
Drug|Vitamin|General Exam|3177,3185|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|COMPLETE
Event|Event|General Exam|3177,3185|false|false|false|||COMPLETE
Finding|Functional Concept|General Exam|3177,3185|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|COMPLETE
Finding|Idea or Concept|General Exam|3177,3185|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|COMPLETE
Procedure|Laboratory Procedure|General Exam|3177,3197|false|false|false|C0009555|Complete Blood Count|COMPLETE BLOOD COUNT
Disorder|Disease or Syndrome|General Exam|3186,3191|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3186,3191|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3186,3191|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|3186,3197|false|false|false|C0005771|Blood Cell Count|BLOOD COUNT
Anatomy|Cell|General Exam|3198,3201|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|3202,3205|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|3202,3205|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|3202,3205|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|3206,3209|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|3206,3209|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|3206,3209|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|3206,3209|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|3210,3213|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|3210,3213|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|3214,3217|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|3214,3217|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|3214,3217|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|3214,3217|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|3214,3217|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|3218,3221|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|3218,3221|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|3218,3221|false|false|false|||MCH
Finding|Gene or Genome|General Exam|3218,3221|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|3218,3221|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|3218,3221|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|3222,3226|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|3231,3234|false|false|false|C0201617|Primed lymphocyte test|Plt
Drug|Chemical Viewed Functionally|General Exam|3299,3304|false|false|false|C0178499|Base|BASIC
Event|Event|General Exam|3299,3304|false|false|false|||BASIC
Finding|Functional Concept|General Exam|3299,3304|false|false|false|C1527178|Basis - conceptual entity|BASIC
Event|Event|General Exam|3305,3316|false|false|false|||COAGULATION
Finding|Organ or Tissue Function|General Exam|3305,3316|false|false|false|C0005778;C1328723|Blood coagulation;Coagulation process|COAGULATION
Finding|Physiologic Function|General Exam|3305,3316|false|false|false|C0005778;C1328723|Blood coagulation;Coagulation process|COAGULATION
Lab|Laboratory or Test Result|General Exam|3305,3316|false|false|false|C0427579|Blood coagulation pathway observation|COAGULATION
Procedure|Laboratory Procedure|General Exam|3305,3316|false|false|false|C0005790;C0441509;C1561952|Blood coagulation tests;Coagulation procedure;Observation Method - Coagulation|COAGULATION
Procedure|Therapeutic or Preventive Procedure|General Exam|3305,3316|false|false|false|C0005790;C0441509;C1561952|Blood coagulation tests;Coagulation procedure;Observation Method - Coagulation|COAGULATION
Disorder|Neoplastic Process|General Exam|3322,3325|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|General Exam|3322,3325|false|false|false|||PTT
Procedure|Laboratory Procedure|General Exam|3322,3325|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Event|Event|General Exam|3327,3330|false|false|false|||PLT
Procedure|Laboratory Procedure|General Exam|3327,3330|false|false|false|C0201617|Primed lymphocyte test|PLT
Attribute|Clinical Attribute|General Exam|3332,3335|false|false|false|C0368980|Coagulation tissue factor induced.INR|INR
Event|Event|General Exam|3332,3335|false|false|false|||INR
Procedure|Laboratory Procedure|General Exam|3332,3335|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Therapeutic or Preventive Procedure|General Exam|3332,3335|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Laboratory Procedure|General Exam|3337,3340|false|false|false|C0201617|Primed lymphocyte test|Plt
Event|Event|General Exam|3365,3374|false|false|false|||Chemistry
Finding|Finding|General Exam|3365,3374|false|false|false|C0079107;C1547978;C2183231|Chemistry Section ID;chemical aspects;diagnostic service sources chemistry (fluid analysis)|Chemistry
Finding|Functional Concept|General Exam|3365,3374|false|false|false|C0079107;C1547978;C2183231|Chemistry Section ID;chemical aspects;diagnostic service sources chemistry (fluid analysis)|Chemistry
Finding|Intellectual Product|General Exam|3365,3374|false|false|false|C0079107;C1547978;C2183231|Chemistry Section ID;chemical aspects;diagnostic service sources chemistry (fluid analysis)|Chemistry
Procedure|Laboratory Procedure|General Exam|3365,3374|false|false|false|C0201682|Chemical procedure|Chemistry
Anatomy|Body Part, Organ, or Organ Component|General Exam|3376,3381|false|false|false|C0022646|Kidney|RENAL
Disorder|Disease or Syndrome|General Exam|3376,3381|false|false|false|C0042075|Urologic Diseases|RENAL
Event|Event|General Exam|3376,3381|false|false|false|||RENAL
Drug|Biologically Active Substance|General Exam|3384,3391|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|General Exam|3384,3391|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|General Exam|3384,3391|false|false|false|C0017725|glucose|GLUCOSE
Event|Event|General Exam|3384,3391|false|false|false|||GLUCOSE
Lab|Laboratory or Test Result|General Exam|3384,3391|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|General Exam|3384,3391|false|false|false|C0337438|Glucose measurement|GLUCOSE
Drug|Biologically Active Substance|General Exam|3392,3399|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|3392,3399|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|3392,3399|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|General Exam|3392,3399|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|3392,3399|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|3420,3424|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|3420,3424|false|false|false|C0005367|Bicarbonates|HCO3
Event|Event|General Exam|3420,3424|false|false|false|||HCO3
Procedure|Laboratory Procedure|General Exam|3420,3424|false|false|false|C0202059|Bicarbonate measurement|HCO3
Finding|Body Substance|Hospital Course|3502,3509|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|3502,3509|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|3502,3509|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|3510,3519|false|false|false|||presented
Event|Occupational Activity|Hospital Course|3545,3552|false|false|false|C0557854|Services|service
Finding|Idea or Concept|Hospital Course|3545,3552|false|false|false|C3245478|ActInformationPrivacyReason - service|service
Event|Event|Hospital Course|3565,3574|false|false|false|||treatment
Finding|Conceptual Entity|Hospital Course|3565,3574|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Hospital Course|3565,3574|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Hospital Course|3565,3574|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3565,3574|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Event|Event|Hospital Course|3586,3594|false|false|false|||hardware
Event|Event|Hospital Course|3612,3619|false|false|false|||surgery
Finding|Finding|Hospital Course|3612,3619|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Hospital Course|3612,3619|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Hospital Course|3612,3619|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3612,3619|false|false|false|C0543467|Operative Surgical Procedures|surgery
Anatomy|Body Location or Region|Hospital Course|3627,3631|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|3627,3631|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|Hospital Course|3627,3631|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3627,3631|false|false|false|C0876917|Procedure on head|head
Event|Event|Hospital Course|3637,3641|false|false|false|||went
Event|Activity|Hospital Course|3684,3691|false|false|false|C1883720|Removing (action)|removal
Event|Event|Hospital Course|3684,3691|false|false|false|||removal
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3684,3691|false|false|false|C0015252;C0185115;C0728940|Excision;Extraction;removal technique|removal
Event|Event|Hospital Course|3703,3711|false|false|false|||hardware
Finding|Body Substance|Hospital Course|3746,3753|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|3746,3753|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|3746,3753|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|3758,3764|false|false|false|||stable
Finding|Intellectual Product|Hospital Course|3758,3764|false|false|false|C1547311|Patient Condition Code - Stable|stable
Disorder|Disease or Syndrome|Hospital Course|3766,3776|false|false|false|C0009450|Communicable Diseases|Infectious
Disorder|Disease or Syndrome|Hospital Course|3766,3784|false|false|false|C0009450|Communicable Diseases|Infectious disease
Disorder|Disease or Syndrome|Hospital Course|3777,3784|false|false|false|C0012634|Disease|disease
Event|Event|Hospital Course|3777,3784|false|false|false|||disease
Event|Event|Hospital Course|3786,3795|false|false|false|||consulted
Finding|Body Substance|Hospital Course|3800,3807|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|3800,3807|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|3800,3807|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|3812,3823|false|false|false|||recommended
Drug|Clinical Drug|Hospital Course|3824,3835|false|false|false|C0016277;C0812735|INJECTION FLUCONAZOLE, 200 MG ADMINISTERED;fluconazole|fluconazole
Drug|Organic Chemical|Hospital Course|3824,3835|false|false|false|C0016277;C0812735|INJECTION FLUCONAZOLE, 200 MG ADMINISTERED;fluconazole|fluconazole
Drug|Pharmacologic Substance|Hospital Course|3824,3835|false|false|false|C0016277;C0812735|INJECTION FLUCONAZOLE, 200 MG ADMINISTERED;fluconazole|fluconazole
Event|Event|Hospital Course|3824,3835|false|false|false|||fluconazole
Event|Event|Hospital Course|3853,3857|false|false|false|||days
Drug|Food|Hospital Course|3862,3867|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|yeast
Drug|Immunologic Factor|Hospital Course|3862,3867|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|yeast
Drug|Indicator, Reagent, or Diagnostic Aid|Hospital Course|3862,3867|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|yeast
Drug|Pharmacologic Substance|Hospital Course|3862,3867|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|yeast
Disorder|Disease or Syndrome|Hospital Course|3862,3877|false|false|false|C0750466|Yeast infection|yeast infection
Disorder|Disease or Syndrome|Hospital Course|3868,3877|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|Hospital Course|3868,3877|false|false|false|||infection
Finding|Pathologic Function|Hospital Course|3868,3877|false|false|false|C3714514|Infection|infection
Drug|Antibiotic|Hospital Course|3882,3888|false|false|false|C0700517|Keflex|Keflex
Drug|Organic Chemical|Hospital Course|3882,3888|false|false|false|C0700517|Keflex|Keflex
Disorder|Mental or Behavioral Dysfunction|Hospital Course|3899,3902|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|3899,3902|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|3899,3902|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|3899,3902|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|3899,3902|false|false|false|C1332410|BID gene|BID
Anatomy|Body Location or Region|Hospital Course|3920,3923|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Hospital Course|3920,3923|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Hospital Course|3920,3923|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3920,3935|false|false|false|C0853245|DVT prophylaxis|DVT prophylaxis
Event|Event|Hospital Course|3924,3935|false|false|false|||prophylaxis
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3924,3935|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Finding|Body Substance|Hospital Course|3941,3948|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|3941,3948|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|3941,3948|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|Hospital Course|3958,3970|false|false|false|C1522438|Subcutaneous Route of Administration|subcutaneous
Drug|Organic Chemical|Hospital Course|3958,3978|false|false|false|C0353681|subcutaneous heparin|subcutaneous heparin
Drug|Pharmacologic Substance|Hospital Course|3958,3978|false|false|false|C0353681|subcutaneous heparin|subcutaneous heparin
Drug|Biologically Active Substance|Hospital Course|3971,3978|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|Hospital Course|3971,3978|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|Hospital Course|3971,3978|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Event|Event|Hospital Course|3971,3978|false|false|false|||heparin
Disorder|Disease or Syndrome|Hospital Course|3984,3987|false|false|false|C0002895;C0271287;C0342788|Anemia, Sickle Cell;Renal carnitine transport defect;Schnyder crystalline corneal dystrophy|SCD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|3984,3987|false|false|false|C5441731|SCD protein, human|SCD
Drug|Enzyme|Hospital Course|3984,3987|false|false|false|C5441731|SCD protein, human|SCD
Finding|Gene or Genome|Hospital Course|3984,3987|false|false|false|C0085298;C1419846;C1420140;C1549989|Doctor of Science;SCD gene;SLC22A5 gene;Sudden Cardiac Death|SCD
Finding|Intellectual Product|Hospital Course|3984,3987|false|false|false|C0085298;C1419846;C1420140;C1549989|Doctor of Science;SCD gene;SLC22A5 gene;Sudden Cardiac Death|SCD
Finding|Pathologic Function|Hospital Course|3984,3987|false|false|false|C0085298;C1419846;C1420140;C1549989|Doctor of Science;SCD gene;SLC22A5 gene;Sudden Cardiac Death|SCD
Event|Event|Hospital Course|3984,3989|false|false|false|||SCD's
Event|Event|Hospital Course|4001,4005|false|false|false|||stay
Finding|Finding|Hospital Course|4015,4019|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Hospital Course|4015,4019|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Hospital Course|4015,4019|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|Hospital Course|4023,4032|false|false|false|||discharge
Finding|Body Substance|Hospital Course|4023,4032|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|4023,4032|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|4023,4032|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|4023,4032|false|false|false|C0030685|Patient Discharge|discharge
Finding|Body Substance|Hospital Course|4038,4045|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|4038,4045|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|4038,4045|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|4050,4054|false|false|false|||able
Finding|Finding|Hospital Course|4050,4054|false|false|false|C1299581|Able (qualifier value)|able
Event|Event|Hospital Course|4090,4094|false|false|false|||able
Finding|Finding|Hospital Course|4090,4094|false|false|false|C1299581|Able (qualifier value)|able
Event|Event|Hospital Course|4098,4102|false|false|false|||void
Event|Event|Hospital Course|4126,4130|false|false|false|||able
Finding|Finding|Hospital Course|4126,4130|false|false|false|C1299581|Able (qualifier value)|able
Attribute|Clinical Attribute|Hospital Course|4145,4154|false|false|false|C4255433||agreement
Event|Event|Hospital Course|4145,4154|false|false|false|||agreement
Finding|Intellectual Product|Hospital Course|4145,4154|false|false|false|C0680240;C4255373|Agreement;Agreement (document)|agreement
Finding|Social Behavior|Hospital Course|4145,4154|false|false|false|C0680240;C4255373|Agreement;Agreement (document)|agreement
Event|Event|Hospital Course|4159,4172|false|false|false|||understanding
Finding|Mental Process|Hospital Course|4159,4172|false|false|false|C0162340|Comprehension|understanding
Finding|Body Substance|Hospital Course|4180,4189|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|4180,4189|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|4180,4189|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|4180,4189|false|false|false|C0030685|Patient Discharge|discharge
Attribute|Clinical Attribute|Hospital Course|4180,4194|false|false|false|C2745873||discharge plan
Finding|Intellectual Product|Hospital Course|4180,4194|false|false|false|C2735970|Discharge plan|discharge plan
Procedure|Health Care Activity|Hospital Course|4180,4194|false|false|false|C0012622|Discharge Planning|discharge plan
Disorder|Disease or Syndrome|Hospital Course|4190,4194|false|false|false|C0270724|Infantile Neuroaxonal Dystrophy|plan
Event|Event|Hospital Course|4190,4194|false|false|false|||plan
Finding|Functional Concept|Hospital Course|4190,4194|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Intellectual Product|Hospital Course|4190,4194|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Mental Process|Hospital Course|4190,4194|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Attribute|Clinical Attribute|Hospital Course|4198,4209|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|4198,4209|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|4198,4209|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|4198,4209|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|4198,4222|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|4213,4222|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|4213,4222|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|Hospital Course|4241,4251|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Hospital Course|4241,4251|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|Hospital Course|4241,4256|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|Hospital Course|4252,4256|false|false|false|||list
Finding|Intellectual Product|Hospital Course|4252,4256|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|Hospital Course|4264,4274|false|false|false|||inaccurate
Event|Event|Hospital Course|4279,4287|false|false|false|||requires
Event|Event|Hospital Course|4296,4309|false|false|false|||investigation
Finding|Intellectual Product|Hospital Course|4296,4309|false|false|false|C1552578|Act Class - investigation|investigation
Procedure|Health Care Activity|Hospital Course|4296,4309|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|investigation
Drug|Organic Chemical|Hospital Course|4314,4324|false|false|false|C0002333|alprazolam|ALPRAZolam
Drug|Pharmacologic Substance|Hospital Course|4314,4324|false|false|false|C0002333|alprazolam|ALPRAZolam
Event|Event|Hospital Course|4335,4338|false|false|false|||TID
Drug|Hazardous or Poisonous Substance|Hospital Course|4343,4355|false|false|false|C0004482|azathioprine|Azathioprine
Drug|Organic Chemical|Hospital Course|4343,4355|false|false|false|C0004482|azathioprine|Azathioprine
Drug|Pharmacologic Substance|Hospital Course|4343,4355|false|false|false|C0004482|azathioprine|Azathioprine
Disorder|Mental or Behavioral Dysfunction|Hospital Course|4366,4369|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4366,4369|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|4366,4369|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|4366,4369|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|4366,4369|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|4374,4385|false|false|false|C0012125|dicyclomine|DiCYCLOmine
Drug|Pharmacologic Substance|Hospital Course|4374,4385|false|false|false|C0012125|dicyclomine|DiCYCLOmine
Finding|Gene or Genome|Hospital Course|4399,4402|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Location or Region|Hospital Course|4403,4412|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|Hospital Course|4403,4417|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|Hospital Course|4413,4417|false|false|false|C2598155||pain
Event|Event|Hospital Course|4413,4417|false|false|false|||pain
Finding|Functional Concept|Hospital Course|4413,4417|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|4413,4417|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|4422,4433|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|4422,4433|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|4422,4444|false|false|false|C0939232|fluticasone / salmeterol|Fluticasone-Salmeterol
Drug|Organic Chemical|Hospital Course|4422,4451|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Pharmacologic Substance|Hospital Course|4422,4451|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Organic Chemical|Hospital Course|4434,4444|false|false|false|C0073992|salmeterol|Salmeterol
Drug|Pharmacologic Substance|Hospital Course|4434,4444|false|false|false|C0073992|salmeterol|Salmeterol
Event|Event|Hospital Course|4445,4451|false|false|false|||Diskus
Drug|Biomedical or Dental Material|Hospital Course|4464,4467|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Organic Chemical|Hospital Course|4464,4467|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Pharmacologic Substance|Hospital Course|4464,4467|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Event|Event|Hospital Course|4464,4467|false|false|false|||INH
Finding|Functional Concept|Hospital Course|4464,4467|false|false|false|C0205535|Inhalation Route of Administration|INH
Disorder|Mental or Behavioral Dysfunction|Hospital Course|4471,4474|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4471,4474|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|4471,4474|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|4471,4474|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|4471,4474|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|4479,4490|false|false|false|C0020264|hydrocodone|Hydrocodone
Drug|Pharmacologic Substance|Hospital Course|4479,4490|false|false|false|C0020264|hydrocodone|Hydrocodone
Drug|Organic Chemical|Hospital Course|4491,4504|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|4491,4504|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Hospital Course|4491,4504|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|4491,4504|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Biomedical or Dental Material|Hospital Course|4519,4522|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|Hospital Course|4519,4522|false|false|false|||TAB
Event|Event|Hospital Course|4526,4529|false|false|false|||Q4H
Finding|Gene or Genome|Hospital Course|4530,4533|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|4534,4538|false|false|false|C2598155||pain
Event|Event|Hospital Course|4534,4538|false|false|false|||pain
Finding|Functional Concept|Hospital Course|4534,4538|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|4534,4538|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4543,4553|false|false|false|C0666743|infliximab|Infliximab
Drug|Immunologic Factor|Hospital Course|4543,4553|false|false|false|C0666743|infliximab|Infliximab
Drug|Pharmacologic Substance|Hospital Course|4543,4553|false|false|false|C0666743|infliximab|Infliximab
Event|Event|Hospital Course|4543,4553|false|false|false|||Infliximab
Procedure|Laboratory Procedure|Hospital Course|4543,4553|false|false|false|C5201962|Drug assay infliximab|Infliximab
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4577,4590|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Hormone|Hospital Course|4577,4590|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Organic Chemical|Hospital Course|4577,4590|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Pharmacologic Substance|Hospital Course|4577,4590|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Event|Event|Hospital Course|4577,4590|false|false|false|||Levothyroxine
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4577,4597|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Hormone|Hospital Course|4577,4597|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Pharmacologic Substance|Hospital Course|4577,4597|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Biologically Active Substance|Hospital Course|4591,4597|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|4591,4597|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|4591,4597|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|4591,4597|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|4591,4597|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|4591,4597|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Organic Chemical|Hospital Course|4618,4628|false|false|false|C0127615|mesalamine|Mesalamine
Drug|Pharmacologic Substance|Hospital Course|4618,4628|false|false|false|C0127615|mesalamine|Mesalamine
Drug|Organic Chemical|Hospital Course|4647,4657|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Pharmacologic Substance|Hospital Course|4647,4657|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Organic Chemical|Hospital Course|4678,4690|false|false|false|C0033405|promethazine|Promethazine
Drug|Pharmacologic Substance|Hospital Course|4678,4690|false|false|false|C0033405|promethazine|Promethazine
Event|Event|Hospital Course|4704,4707|false|false|false|||PRN
Finding|Gene or Genome|Hospital Course|4704,4707|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|Hospital Course|4717,4727|false|false|false|C0076829|topiramate|Topiramate
Drug|Pharmacologic Substance|Hospital Course|4717,4727|false|false|false|C0076829|topiramate|Topiramate
Event|Event|Hospital Course|4717,4727|false|false|false|||Topiramate
Procedure|Laboratory Procedure|Hospital Course|4717,4727|false|false|false|C0519827|Topiramate measurement|Topiramate
Drug|Organic Chemical|Hospital Course|4717,4737|false|false|false|C0723778|Topamax|Topiramate (Topamax)
Drug|Pharmacologic Substance|Hospital Course|4717,4737|false|false|false|C0723778|Topamax|Topiramate (Topamax)
Drug|Organic Chemical|Hospital Course|4729,4736|false|false|false|C0723778|Topamax|Topamax
Drug|Pharmacologic Substance|Hospital Course|4729,4736|false|false|false|C0723778|Topamax|Topamax
Disorder|Mental or Behavioral Dysfunction|Hospital Course|4748,4751|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4748,4751|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|4748,4751|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|4748,4751|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|4748,4751|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|4757,4768|false|false|false|C0078569|venlafaxine|Venlafaxine
Drug|Pharmacologic Substance|Hospital Course|4757,4768|false|false|false|C0078569|venlafaxine|Venlafaxine
Event|Event|Hospital Course|4757,4768|false|false|false|||Venlafaxine
Drug|Organic Chemical|Hospital Course|4793,4801|false|false|false|C0078839|zolpidem|Zolpidem
Drug|Pharmacologic Substance|Hospital Course|4793,4801|false|false|false|C0078839|zolpidem|Zolpidem
Event|Event|Hospital Course|4793,4801|false|false|false|||Zolpidem
Drug|Organic Chemical|Hospital Course|4793,4810|false|false|false|C0724725|zolpidem tartrate|Zolpidem Tartrate
Drug|Pharmacologic Substance|Hospital Course|4793,4810|false|false|false|C0724725|zolpidem tartrate|Zolpidem Tartrate
Drug|Organic Chemical|Hospital Course|4802,4810|false|false|false|C0039328;C0144544|Tartrates;tartrate|Tartrate
Drug|Pharmacologic Substance|Hospital Course|4802,4810|false|false|false|C0039328;C0144544|Tartrates;tartrate|Tartrate
Event|Event|Hospital Course|4827,4836|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|4827,4836|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|4827,4836|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|4827,4836|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|4827,4836|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|4827,4848|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|4837,4848|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|4837,4848|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|4837,4848|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|4837,4848|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|4853,4863|false|false|false|C0002333|alprazolam|ALPRAZolam
Drug|Pharmacologic Substance|Hospital Course|4853,4863|false|false|false|C0002333|alprazolam|ALPRAZolam
Event|Event|Hospital Course|4874,4877|false|false|false|||TID
Drug|Hazardous or Poisonous Substance|Hospital Course|4882,4894|false|false|false|C0004482|azathioprine|Azathioprine
Drug|Organic Chemical|Hospital Course|4882,4894|false|false|false|C0004482|azathioprine|Azathioprine
Drug|Pharmacologic Substance|Hospital Course|4882,4894|false|false|false|C0004482|azathioprine|Azathioprine
Disorder|Mental or Behavioral Dysfunction|Hospital Course|4905,4908|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4905,4908|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|4905,4908|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|4905,4908|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|4905,4908|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|4913,4924|false|false|false|C0012125|dicyclomine|DiCYCLOmine
Drug|Pharmacologic Substance|Hospital Course|4913,4924|false|false|false|C0012125|dicyclomine|DiCYCLOmine
Finding|Gene or Genome|Hospital Course|4938,4941|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Location or Region|Hospital Course|4942,4951|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|Hospital Course|4942,4956|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|Hospital Course|4952,4956|false|false|false|C2598155||pain
Event|Event|Hospital Course|4952,4956|false|false|false|||pain
Finding|Functional Concept|Hospital Course|4952,4956|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|4952,4956|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4961,4974|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Hormone|Hospital Course|4961,4974|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Organic Chemical|Hospital Course|4961,4974|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Pharmacologic Substance|Hospital Course|4961,4974|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Event|Event|Hospital Course|4961,4974|false|false|false|||Levothyroxine
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4961,4981|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Hormone|Hospital Course|4961,4981|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Pharmacologic Substance|Hospital Course|4961,4981|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Biologically Active Substance|Hospital Course|4975,4981|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|4975,4981|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|4975,4981|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|4975,4981|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|4975,4981|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|4975,4981|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Organic Chemical|Hospital Course|5002,5012|false|false|false|C0127615|mesalamine|Mesalamine
Drug|Pharmacologic Substance|Hospital Course|5002,5012|false|false|false|C0127615|mesalamine|Mesalamine
Drug|Organic Chemical|Hospital Course|5031,5041|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Pharmacologic Substance|Hospital Course|5031,5041|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Organic Chemical|Hospital Course|5061,5071|false|false|false|C0076829|topiramate|Topiramate
Drug|Pharmacologic Substance|Hospital Course|5061,5071|false|false|false|C0076829|topiramate|Topiramate
Event|Event|Hospital Course|5061,5071|false|false|false|||Topiramate
Procedure|Laboratory Procedure|Hospital Course|5061,5071|false|false|false|C0519827|Topiramate measurement|Topiramate
Drug|Organic Chemical|Hospital Course|5061,5081|false|false|false|C0723778|Topamax|Topiramate (Topamax)
Drug|Pharmacologic Substance|Hospital Course|5061,5081|false|false|false|C0723778|Topamax|Topiramate (Topamax)
Drug|Organic Chemical|Hospital Course|5073,5080|false|false|false|C0723778|Topamax|Topamax
Drug|Pharmacologic Substance|Hospital Course|5073,5080|false|false|false|C0723778|Topamax|Topamax
Disorder|Mental or Behavioral Dysfunction|Hospital Course|5092,5095|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5092,5095|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|5092,5095|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|5092,5095|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|5092,5095|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|5100,5111|false|false|false|C0078569|venlafaxine|Venlafaxine
Drug|Pharmacologic Substance|Hospital Course|5100,5111|false|false|false|C0078569|venlafaxine|Venlafaxine
Event|Event|Hospital Course|5100,5111|false|false|false|||Venlafaxine
Drug|Organic Chemical|Hospital Course|5135,5143|false|false|false|C0078839|zolpidem|Zolpidem
Drug|Pharmacologic Substance|Hospital Course|5135,5143|false|false|false|C0078839|zolpidem|Zolpidem
Event|Event|Hospital Course|5135,5143|false|false|false|||Zolpidem
Drug|Organic Chemical|Hospital Course|5135,5152|false|false|false|C0724725|zolpidem tartrate|Zolpidem Tartrate
Drug|Pharmacologic Substance|Hospital Course|5135,5152|false|false|false|C0724725|zolpidem tartrate|Zolpidem Tartrate
Drug|Organic Chemical|Hospital Course|5144,5152|false|false|false|C0039328;C0144544|Tartrates;tartrate|Tartrate
Drug|Pharmacologic Substance|Hospital Course|5144,5152|false|false|false|C0039328;C0144544|Tartrates;tartrate|Tartrate
Drug|Organic Chemical|Hospital Course|5170,5181|false|false|false|C0020264|hydrocodone|Hydrocodone
Drug|Pharmacologic Substance|Hospital Course|5170,5181|false|false|false|C0020264|hydrocodone|Hydrocodone
Drug|Organic Chemical|Hospital Course|5182,5195|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|5182,5195|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Hospital Course|5182,5195|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|5182,5195|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Biomedical or Dental Material|Hospital Course|5210,5213|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|Hospital Course|5210,5213|false|false|false|||TAB
Event|Event|Hospital Course|5217,5220|false|false|false|||Q4H
Finding|Gene or Genome|Hospital Course|5221,5224|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|5225,5229|false|false|false|C2598155||pain
Event|Event|Hospital Course|5225,5229|false|false|false|||pain
Finding|Functional Concept|Hospital Course|5225,5229|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|5225,5229|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|5235,5248|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|5235,5248|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Hospital Course|5235,5248|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|5235,5248|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|Hospital Course|5267,5270|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|5271,5282|false|false|false|||temperature
Procedure|Health Care Activity|Hospital Course|5271,5282|false|false|false|C0886414|Body temperature measurement|temperature
Attribute|Clinical Attribute|Hospital Course|5284,5288|false|false|false|C2598155||pain
Event|Event|Hospital Course|5284,5288|false|false|false|||pain
Finding|Functional Concept|Hospital Course|5284,5288|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|5284,5288|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|5294,5302|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|5294,5302|false|false|false|C1692318|docusate|Docusate
Event|Event|Hospital Course|5294,5302|false|false|false|||Docusate
Drug|Organic Chemical|Hospital Course|5294,5309|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|Hospital Course|5294,5309|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|Hospital Course|5303,5309|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|5303,5309|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|5303,5309|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|5303,5309|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|5303,5309|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|5303,5309|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|Hospital Course|5320,5323|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5320,5323|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|5320,5323|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|5320,5323|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|5320,5323|false|false|false|C1332410|BID gene|BID
Finding|Gene or Genome|Hospital Course|5324,5327|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|5328,5340|false|false|false|||constipation
Finding|Sign or Symptom|Hospital Course|5328,5340|false|false|false|C0009806|Constipation|constipation
Drug|Organic Chemical|Hospital Course|5346,5354|false|false|false|C1692318|docusate|docusate
Drug|Pharmacologic Substance|Hospital Course|5346,5354|false|false|false|C1692318|docusate|docusate
Drug|Organic Chemical|Hospital Course|5346,5361|false|false|false|C0243237|docusate sodium|docusate sodium
Drug|Pharmacologic Substance|Hospital Course|5346,5361|false|false|false|C0243237|docusate sodium|docusate sodium
Drug|Biologically Active Substance|Hospital Course|5355,5361|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|Hospital Course|5355,5361|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|Hospital Course|5355,5361|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Event|Event|Hospital Course|5355,5361|false|false|false|||sodium
Finding|Physiologic Function|Hospital Course|5355,5361|false|false|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|Hospital Course|5355,5361|false|false|false|C0337443|Sodium measurement|sodium
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5373,5380|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|Hospital Course|5373,5380|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|Hospital Course|5373,5380|false|false|false|C0006935|capsule (pharmacologic)|capsule
Finding|Functional Concept|Hospital Course|5384,5392|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|5387,5392|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|5387,5392|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|Hospital Course|5401,5404|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|5401,5404|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5416,5423|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|5416,5423|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|5416,5423|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Event|Event|Hospital Course|5424,5431|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|5424,5431|false|false|false|C0807726|refill|Refills
Drug|Clinical Drug|Hospital Course|5439,5450|false|false|false|C0016277;C0812735|INJECTION FLUCONAZOLE, 200 MG ADMINISTERED;fluconazole|Fluconazole
Drug|Organic Chemical|Hospital Course|5439,5450|false|false|false|C0016277;C0812735|INJECTION FLUCONAZOLE, 200 MG ADMINISTERED;fluconazole|Fluconazole
Drug|Pharmacologic Substance|Hospital Course|5439,5450|false|false|false|C0016277;C0812735|INJECTION FLUCONAZOLE, 200 MG ADMINISTERED;fluconazole|Fluconazole
Drug|Pharmacologic Substance|Hospital Course|5466,5474|false|false|false|C0720099|Duration brand of oxymetazoline|Duration
Event|Event|Hospital Course|5466,5474|false|false|false|||Duration
Drug|Clinical Drug|Hospital Course|5488,5499|false|false|false|C0016277;C0812735|INJECTION FLUCONAZOLE, 200 MG ADMINISTERED;fluconazole|fluconazole
Drug|Organic Chemical|Hospital Course|5488,5499|false|false|false|C0016277;C0812735|INJECTION FLUCONAZOLE, 200 MG ADMINISTERED;fluconazole|fluconazole
Drug|Pharmacologic Substance|Hospital Course|5488,5499|false|false|false|C0016277;C0812735|INJECTION FLUCONAZOLE, 200 MG ADMINISTERED;fluconazole|fluconazole
Event|Event|Hospital Course|5488,5499|false|false|false|||fluconazole
Drug|Biomedical or Dental Material|Hospital Course|5509,5515|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|5519,5527|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|5522,5527|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|5522,5527|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Biomedical or Dental Material|Hospital Course|5544,5550|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|5551,5558|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|5551,5558|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|5566,5575|false|false|false|C0030049|oxycodone|OxycoDONE
Drug|Pharmacologic Substance|Hospital Course|5566,5575|false|false|false|C0030049|oxycodone|OxycoDONE
Event|Event|Hospital Course|5566,5575|false|false|false|||OxycoDONE
Procedure|Laboratory Procedure|Hospital Course|5566,5575|false|false|false|C0524222|Oxycodone measurement|OxycoDONE
Finding|Idea or Concept|Hospital Course|5577,5586|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Finding|Intellectual Product|Hospital Course|5577,5586|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Drug|Biomedical or Dental Material|Hospital Course|5577,5594|false|false|false|C1708470|Immediate Release Dosage Form|Immediate Release
Event|Event|Hospital Course|5587,5594|false|false|false|||Release
Finding|Functional Concept|Hospital Course|5587,5594|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|5587,5594|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5587,5594|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Finding|Gene or Genome|Hospital Course|5609,5612|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Finding|Hospital Course|5617,5625|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|Hospital Course|5617,5625|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Attribute|Clinical Attribute|Hospital Course|5627,5631|false|false|false|C2598155||pain
Event|Event|Hospital Course|5627,5631|false|false|false|||pain
Finding|Functional Concept|Hospital Course|5627,5631|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|5627,5631|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|5633,5635|false|false|false|||RX
Drug|Organic Chemical|Hospital Course|5637,5646|false|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|Hospital Course|5637,5646|false|false|false|C0030049|oxycodone|oxycodone
Event|Event|Hospital Course|5637,5646|false|false|false|||oxycodone
Procedure|Laboratory Procedure|Hospital Course|5637,5646|false|false|false|C0524222|Oxycodone measurement|oxycodone
Drug|Biomedical or Dental Material|Hospital Course|5656,5662|false|false|false|C0039225|Tablet Dosage Form|tablet
Event|Event|Hospital Course|5656,5662|false|false|false|||tablet
Finding|Functional Concept|Hospital Course|5666,5674|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|5669,5674|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|5669,5674|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Biomedical or Dental Material|Hospital Course|5706,5712|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|5713,5720|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|5713,5720|false|false|false|C0807726|refill|Refills
Drug|Antibiotic|Hospital Course|5728,5738|false|false|false|C0007716|cephalexin|Cephalexin
Drug|Organic Chemical|Hospital Course|5728,5738|false|false|false|C0007716|cephalexin|Cephalexin
Drug|Pharmacologic Substance|Hospital Course|5754,5762|false|false|false|C0720099|Duration brand of oxymetazoline|Duration
Event|Event|Hospital Course|5754,5762|false|false|false|||Duration
Drug|Antibiotic|Hospital Course|5776,5786|false|false|false|C0007716|cephalexin|cephalexin
Drug|Organic Chemical|Hospital Course|5776,5786|false|false|false|C0007716|cephalexin|cephalexin
Event|Event|Hospital Course|5776,5786|false|false|false|||cephalexin
Drug|Biomedical or Dental Material|Hospital Course|5796,5802|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|5806,5814|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|5809,5814|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|5809,5814|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|Hospital Course|5823,5826|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|5823,5826|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biomedical or Dental Material|Hospital Course|5838,5844|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|5845,5852|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|5845,5852|false|false|false|C0807726|refill|Refills
Event|Event|Hospital Course|5859,5868|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|5859,5868|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|5859,5868|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|5859,5868|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|5859,5868|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|5859,5880|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|5859,5880|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|5869,5880|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|5869,5880|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|5869,5880|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|Hospital Course|5882,5886|false|false|false|||Home
Finding|Idea or Concept|Hospital Course|5882,5886|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|5882,5886|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|5882,5886|false|false|false|C1553498|home health encounter|Home
Event|Event|Hospital Course|5889,5898|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|5889,5898|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|5889,5898|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|5889,5898|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|5889,5898|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|5889,5908|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|5899,5908|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|5899,5908|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|5899,5908|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|5899,5908|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|5899,5908|false|false|false|C0011900|Diagnosis|Diagnosis
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5910,5926|false|false|false|C5453054|Hardware Removal|Hardware removal
Event|Activity|Hospital Course|5919,5926|false|false|false|C1883720|Removing (action)|removal
Event|Event|Hospital Course|5919,5926|false|false|false|||removal
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5919,5926|false|false|false|C0015252;C0185115;C0728940|Excision;Extraction;removal technique|removal
Finding|Mental Process|Discharge Condition|5951,5957|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|5951,5964|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|5951,5964|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|5958,5964|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|5958,5964|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|5966,5971|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|5966,5971|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|5976,5984|false|false|false|||coherent
Finding|Finding|Discharge Condition|5976,5984|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|5986,5991|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|5986,6008|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|5986,6008|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|5995,6008|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|5995,6008|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|5995,6008|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|6010,6015|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|6010,6015|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|6010,6015|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|6010,6015|false|false|false|||Alert
Finding|Finding|Discharge Condition|6010,6015|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|6010,6015|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|6010,6015|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|6020,6031|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|6020,6031|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|6033,6041|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|6033,6041|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|6033,6041|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|6042,6048|false|false|false|C5889824||Status
Event|Event|Discharge Condition|6042,6048|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|6042,6048|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|6050,6060|false|false|false|||Ambulatory
Finding|Functional Concept|Discharge Condition|6050,6060|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|6050,6060|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|6050,6060|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|6050,6060|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|6063,6074|false|false|false|||Independent
Finding|Finding|Discharge Condition|6063,6074|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Condition|6063,6074|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Event|Event|Discharge Instructions|6112,6116|false|false|false|||take
Drug|Clinical Drug|Discharge Instructions|6117,6128|false|false|false|C0016277;C0812735|INJECTION FLUCONAZOLE, 200 MG ADMINISTERED;fluconazole|Fluconazole
Drug|Organic Chemical|Discharge Instructions|6117,6128|false|false|false|C0016277;C0812735|INJECTION FLUCONAZOLE, 200 MG ADMINISTERED;fluconazole|Fluconazole
Drug|Pharmacologic Substance|Discharge Instructions|6117,6128|false|false|false|C0016277;C0812735|INJECTION FLUCONAZOLE, 200 MG ADMINISTERED;fluconazole|Fluconazole
Event|Event|Discharge Instructions|6129,6134|false|false|false|||200mg
Finding|Intellectual Product|Discharge Instructions|6135,6139|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Antibiotic|Discharge Instructions|6171,6177|false|false|false|C0700517|Keflex|Keflex
Drug|Organic Chemical|Discharge Instructions|6171,6177|false|false|false|C0700517|Keflex|Keflex
Event|Event|Discharge Instructions|6171,6177|false|false|false|||Keflex
Disorder|Injury or Poisoning|Discharge Instructions|6193,6198|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Event|Event|Discharge Instructions|6193,6198|false|false|false|||wound
Finding|Body Substance|Discharge Instructions|6193,6198|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|Discharge Instructions|6193,6198|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|Discharge Instructions|6193,6198|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Pathologic Function|Discharge Instructions|6193,6208|false|false|false|C0043241|Wound Infection|wound infection
Disorder|Disease or Syndrome|Discharge Instructions|6199,6208|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|Discharge Instructions|6199,6208|false|false|false|||infection
Finding|Pathologic Function|Discharge Instructions|6199,6208|false|false|false|C3714514|Infection|infection
Attribute|Clinical Attribute|Discharge Instructions|6212,6221|false|false|false|C1382187|Clearance of substance|Clearance
Event|Event|Discharge Instructions|6212,6221|false|false|false|||Clearance
Phenomenon|Natural Phenomenon or Process|Discharge Instructions|6212,6221|false|false|false|C2825073|Clearance [PK]|Clearance
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|6212,6221|false|false|false|C4554548|Clearance procedure|Clearance
Event|Event|Discharge Instructions|6225,6230|false|false|false|||drive
Finding|Mental Process|Discharge Instructions|6225,6230|false|false|false|C0013126|Intrinsic drive|drive
Event|Event|Discharge Instructions|6235,6241|false|false|false|||return
Event|Occupational Activity|Discharge Instructions|6245,6249|false|false|false|C0043227|Work|work
Event|Event|Discharge Instructions|6258,6267|false|false|false|||addressed
Event|Event|Discharge Instructions|6292,6298|false|false|false|||office
Finding|Idea or Concept|Discharge Instructions|6292,6298|false|false|false|C1549636|Address type - Office|office
Procedure|Health Care Activity|Discharge Instructions|6292,6304|false|false|false|C0028900|Office Visits|office visit
Event|Event|Discharge Instructions|6299,6304|false|false|false|||visit
Finding|Social Behavior|Discharge Instructions|6299,6304|false|false|false|C0545082|Visit|visit
Event|Event|Discharge Instructions|6306,6310|false|false|false|||CALL
Finding|Functional Concept|Discharge Instructions|6306,6310|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|CALL
Finding|Gene or Genome|Discharge Instructions|6306,6310|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|CALL
Finding|Intellectual Product|Discharge Instructions|6306,6310|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|CALL
Finding|Mental Process|Discharge Instructions|6306,6310|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|CALL
Attribute|Clinical Attribute|Discharge Instructions|6316,6323|false|false|false|C5444295||SURGEON
Event|Event|Discharge Instructions|6316,6323|false|false|false|||SURGEON
Event|Event|Discharge Instructions|6343,6353|true|false|false|||EXPERIENCE
Finding|Mental Process|Discharge Instructions|6343,6353|true|false|false|C0237607;C0596545|Experience;Experience (Practice)|EXPERIENCE
Event|Event|Discharge Instructions|6354,6357|false|false|false|||ANY
Finding|Finding|Discharge Instructions|6378,6381|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Finding|Idea or Concept|Discharge Instructions|6378,6381|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Finding|Finding|Discharge Instructions|6378,6387|false|false|false|C0746890|new onset|New onset
Event|Event|Discharge Instructions|6382,6387|false|false|false|||onset
Event|Event|Discharge Instructions|6391,6398|false|false|false|||tremors
Finding|Sign or Symptom|Discharge Instructions|6391,6398|false|false|false|C0040822|Tremor|tremors
Event|Event|Discharge Instructions|6402,6410|false|false|false|||seizures
Finding|Sign or Symptom|Discharge Instructions|6402,6410|false|false|false|C0036572|Seizures|seizures
Disorder|Mental or Behavioral Dysfunction|Discharge Instructions|6417,6426|true|false|false|C0009676|Confusion|confusion
Event|Event|Discharge Instructions|6417,6426|true|false|false|||confusion
Finding|Finding|Discharge Instructions|6417,6426|true|false|false|C0683369|Clouded consciousness|confusion
Event|Event|Discharge Instructions|6430,6436|true|false|false|||change
Finding|Functional Concept|Discharge Instructions|6430,6436|true|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|6430,6436|true|false|false|C4319952|Change - procedure|change
Finding|Functional Concept|Discharge Instructions|6430,6439|true|false|false|C0392747|Changing|change in
Attribute|Clinical Attribute|Discharge Instructions|6430,6453|true|false|false|C5774124||change in mental status
Finding|Finding|Discharge Instructions|6430,6453|true|false|false|C0856054|Mental status changes|change in mental status
Finding|Mental Process|Discharge Instructions|6440,6446|true|false|false|C0229992|Psyche structure|mental
Attribute|Clinical Attribute|Discharge Instructions|6440,6453|true|false|false|C0488568;C0488569||mental status
Finding|Finding|Discharge Instructions|6440,6453|true|false|false|C0278060|Mental state|mental status
Attribute|Clinical Attribute|Discharge Instructions|6447,6453|true|false|false|C5889824||status
Event|Event|Discharge Instructions|6447,6453|true|false|false|||status
Finding|Idea or Concept|Discharge Instructions|6447,6453|true|false|false|C1546481|What subject filter - Status|status
Event|Event|Discharge Instructions|6461,6469|true|false|false|||numbness
Finding|Finding|Discharge Instructions|6461,6469|true|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|Discharge Instructions|6461,6469|true|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Disorder|Disease or Syndrome|Discharge Instructions|6471,6479|true|false|false|C0030554|Paresthesia|tingling
Event|Event|Discharge Instructions|6471,6479|true|false|false|||tingling
Finding|Sign or Symptom|Discharge Instructions|6471,6479|true|false|false|C2242996|Has tingling sensation|tingling
Event|Event|Discharge Instructions|6481,6489|true|false|false|||weakness
Finding|Sign or Symptom|Discharge Instructions|6481,6489|true|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|6498,6509|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Attribute|Clinical Attribute|Discharge Instructions|6512,6516|false|false|false|C2598155||Pain
Event|Event|Discharge Instructions|6512,6516|false|false|false|||Pain
Finding|Functional Concept|Discharge Instructions|6512,6516|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Discharge Instructions|6512,6516|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Event|Event|Discharge Instructions|6520,6528|true|false|false|||headache
Finding|Sign or Symptom|Discharge Instructions|6520,6528|true|false|false|C0018681|Headache|headache
Event|Event|Discharge Instructions|6549,6559|true|false|false|||increasing
Event|Event|Discharge Instructions|6569,6577|true|false|false|||relieved
Attribute|Clinical Attribute|Discharge Instructions|6581,6585|true|false|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|6581,6585|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|6581,6585|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Pharmacologic Substance|Discharge Instructions|6586,6596|true|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Discharge Instructions|6586,6596|true|false|false|||medication
Finding|Intellectual Product|Discharge Instructions|6586,6596|true|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Discharge Instructions|6603,6608|true|false|false|||signs
Finding|Finding|Discharge Instructions|6603,6608|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Discharge Instructions|6603,6608|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Disorder|Disease or Syndrome|Discharge Instructions|6612,6621|true|false|false|C0009450|Communicable Diseases|infection
Event|Event|Discharge Instructions|6612,6621|true|false|false|||infection
Finding|Pathologic Function|Discharge Instructions|6612,6621|true|false|false|C3714514|Infection|infection
Disorder|Injury or Poisoning|Discharge Instructions|6629,6634|true|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Event|Event|Discharge Instructions|6629,6634|true|false|false|||wound
Finding|Body Substance|Discharge Instructions|6629,6634|true|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|Discharge Instructions|6629,6634|true|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|Discharge Instructions|6629,6634|true|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Anatomy|Body Location or Region|Discharge Instructions|6635,6639|true|false|false|C1515974|Anatomic Site|site
Finding|Intellectual Product|Discharge Instructions|6635,6639|true|false|false|C1546778||site
Disorder|Disease or Syndrome|Discharge Instructions|6652,6659|false|false|false|C0041834|Erythema|redness
Event|Event|Discharge Instructions|6652,6659|false|false|false|||redness
Finding|Finding|Discharge Instructions|6652,6659|false|false|false|C0332575|Redness|redness
Event|Event|Discharge Instructions|6672,6680|false|false|false|||swelling
Finding|Finding|Discharge Instructions|6672,6680|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|Discharge Instructions|6672,6680|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Event|Event|Discharge Instructions|6692,6702|false|false|false|||tenderness
Finding|Mental Process|Discharge Instructions|6692,6702|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|Discharge Instructions|6692,6702|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Event|Discharge Instructions|6707,6715|false|false|false|||drainage
Finding|Body Substance|Discharge Instructions|6707,6715|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|Discharge Instructions|6707,6715|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|6707,6715|false|false|false|C0013103|Drainage procedure|drainage
Finding|Finding|Discharge Instructions|6718,6723|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Finding|Sign or Symptom|Discharge Instructions|6718,6723|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Event|Event|Discharge Instructions|6740,6745|false|false|false|||equal
Finding|Intellectual Product|Discharge Instructions|6740,6745|false|false|false|C1549782|Relational Operator - Equal|equal
Procedure|Health Care Activity|Discharge Instructions|6762,6770|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|6771,6783|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|6771,6783|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|6771,6783|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

