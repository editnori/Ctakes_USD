 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|42,51|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|42,51|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|42,56|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|76,85|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|76,85|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|76,90|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|132,135|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|143,150|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|143,150|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|152,160|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Drug|Indicator, Reagent, or Diagnostic Aid|Allergies|178,181|false|false|false|C0013343|Dyes|Dye
Event|Event|Allergies|178,181|false|false|false|||Dye
Drug|Biologically Active Substance|Allergies|183,189|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Drug|Element, Ion, or Isotope|Allergies|183,189|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Drug|Pharmacologic Substance|Allergies|183,189|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Event|Activity|Allergies|190,200|false|false|false|C2700400|Contain (action)|Containing
Finding|Functional Concept|Allergies|190,200|false|false|false|C0332256|Containing (qualifier value)|Containing
Drug|Indicator, Reagent, or Diagnostic Aid|Allergies|201,209|false|false|false|C0009924|Contrast Media|Contrast
Drug|Indicator, Reagent, or Diagnostic Aid|Allergies|201,215|false|false|false|C0009924|Contrast Media|Contrast Media
Anatomy|Tissue|Allergies|210,215|false|false|false|C0162867;C1254021|Media layer;Tunica Media|Media
Finding|Intellectual Product|Allergies|210,215|false|false|false|C0009458;C0677540|Communications Media;PAMS Media|Media
Drug|Organic Chemical|Allergies|218,227|false|false|false|C0030049|oxycodone|Oxycodone
Drug|Pharmacologic Substance|Allergies|218,227|false|false|false|C0030049|oxycodone|Oxycodone
Event|Event|Allergies|218,227|false|false|false|||Oxycodone
Procedure|Laboratory Procedure|Allergies|218,227|false|false|false|C0524222|Oxycodone measurement|Oxycodone
Drug|Organic Chemical|Allergies|231,241|false|false|false|C0055729|cilostazol|cilostazol
Drug|Pharmacologic Substance|Allergies|231,241|false|false|false|C0055729|cilostazol|cilostazol
Event|Event|Allergies|231,241|false|false|false|||cilostazol
Drug|Organic Chemical|Allergies|244,255|false|false|false|C1569608|varenicline|Varenicline
Drug|Pharmacologic Substance|Allergies|244,255|false|false|false|C1569608|varenicline|Varenicline
Event|Event|Allergies|244,255|false|false|false|||Varenicline
Event|Event|Allergies|258,267|false|false|false|||Attending
Finding|Functional Concept|Allergies|258,267|false|false|false|C1999232|Attending (action)|Attending
Drug|Organic Chemical|Chief Complaint|293,298|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|Chief Complaint|293,298|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|Chief Complaint|293,298|false|false|false|||cough
Finding|Sign or Symptom|Chief Complaint|293,298|false|false|false|C0010200|Coughing|cough
Event|Event|Chief Complaint|300,307|false|false|false|||dyspnea
Finding|Finding|Chief Complaint|300,307|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|Chief Complaint|300,307|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Classification|Chief Complaint|310,315|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|316,324|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|316,324|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|328,346|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|337,346|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|337,346|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|337,346|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|337,346|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|337,346|false|false|false|C0184661|Interventional procedure|Procedure
Disorder|Disease or Syndrome|History of Present Illness|384,387|true|false|false|C0268529|Proline dehydrogenase deficiency|HPI
Event|Event|History of Present Illness|384,387|true|false|false|||HPI
Finding|Finding|History of Present Illness|384,387|true|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Finding|Molecular Function|History of Present Illness|384,387|true|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Finding|Idea or Concept|History of Present Illness|393,397|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|History of Present Illness|393,397|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|History of Present Illness|398,401|false|false|false|||old
Event|Event|History of Present Illness|414,421|false|false|false|||history
Finding|Conceptual Entity|History of Present Illness|414,421|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|414,421|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|414,421|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|414,424|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|History of Present Illness|425,429|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|History of Present Illness|425,429|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|History of Present Illness|425,429|false|false|false|||COPD
Finding|Gene or Genome|History of Present Illness|425,429|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Idea or Concept|History of Present Illness|434,438|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|History of Present Illness|434,438|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|History of Present Illness|434,438|false|false|false|C1553498|home health encounter|home
Disorder|Disease or Syndrome|History of Present Illness|444,447|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|History of Present Illness|444,447|false|false|false|||HTN
Event|Event|History of Present Illness|455,463|false|false|false|||admitted
Event|Event|History of Present Illness|469,476|false|false|false|||dyspnea
Finding|Finding|History of Present Illness|469,476|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|History of Present Illness|469,476|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Drug|Organic Chemical|History of Present Illness|481,486|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|481,486|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|History of Present Illness|481,486|false|false|false|||cough
Finding|Sign or Symptom|History of Present Illness|481,486|false|false|false|C0010200|Coughing|cough
Event|Event|History of Present Illness|494,500|false|false|false|||states
Anatomy|Body Location or Region|History of Present Illness|501,504|false|false|false|C2338258|Cranial incision point|inc
Event|Event|History of Present Illness|505,512|false|false|false|||dyspnea
Finding|Finding|History of Present Illness|505,512|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|History of Present Illness|505,512|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Event|Event|History of Present Illness|537,544|false|false|false|||episode
Anatomy|Body Location or Region|History of Present Illness|562,567|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|562,567|false|false|false|C0741025|Chest problem|chest
Finding|Sign or Symptom|History of Present Illness|562,576|false|false|false|C0438716|Chest pressure|chest pressure
Event|Event|History of Present Illness|568,576|false|false|false|||pressure
Finding|Finding|History of Present Illness|568,576|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|History of Present Illness|568,576|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|History of Present Illness|568,576|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|History of Present Illness|568,576|false|false|false|C0033095||pressure
Event|Event|History of Present Illness|585,592|false|false|false|||2minuts
Event|Event|History of Present Illness|628,632|false|false|false|||home
Finding|Idea or Concept|History of Present Illness|628,632|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|History of Present Illness|628,632|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|History of Present Illness|628,632|false|false|false|C1553498|home health encounter|home
Event|Event|History of Present Illness|640,646|true|false|false|||fevers
Finding|Sign or Symptom|History of Present Illness|640,646|true|false|false|C0015967|Fever|fevers
Event|Event|History of Present Illness|647,653|true|false|false|||chills
Finding|Sign or Symptom|History of Present Illness|647,653|true|false|false|C0085593|Chills|chills
Anatomy|Body Location or Region|History of Present Illness|657,660|true|false|false|C0000726;C0449202|ABD (body structure);Abdomen|abd
Disorder|Cell or Molecular Dysfunction|History of Present Illness|657,660|true|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|abd
Finding|Body Substance|History of Present Illness|668,675|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|668,675|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|668,675|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|History of Present Illness|689,697|false|false|false|||admitted
Disorder|Disease or Syndrome|History of Present Illness|712,716|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|History of Present Illness|712,716|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|History of Present Illness|712,716|false|false|false|||COPD
Finding|Gene or Genome|History of Present Illness|712,716|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|History of Present Illness|717,722|false|false|false|||flare
Finding|Finding|History of Present Illness|717,722|false|false|false|C1517205;C3540542|Exacerbation of cGVHD;Flare|flare
Finding|Sign or Symptom|History of Present Illness|717,722|false|false|false|C1517205;C3540542|Exacerbation of cGVHD;Flare|flare
Disorder|Disease or Syndrome|History of Present Illness|728,732|false|false|false|C0004238|Atrial Fibrillation|afib
Event|Event|History of Present Illness|728,732|false|false|false|||afib
Lab|Laboratory or Test Result|History of Present Illness|728,732|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|afib
Event|Event|History of Present Illness|738,741|false|false|false|||RVR
Finding|Finding|History of Present Illness|738,741|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Finding|Gene or Genome|History of Present Illness|738,741|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Drug|Antibiotic|History of Present Illness|765,777|true|true|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|History of Present Illness|765,777|true|true|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|History of Present Illness|765,777|true|true|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Event|Event|History of Present Illness|765,777|true|false|false|||azithromycin
Event|Event|History of Present Illness|786,793|true|false|false|||concern
Finding|Idea or Concept|History of Present Illness|786,793|true|false|false|C2699424|Concern|concern
Event|Event|History of Present Illness|802,814|false|false|false|||prolongation
Event|Event|History of Present Illness|826,833|false|false|false|||treated
Drug|Antibiotic|History of Present Illness|840,851|false|false|false|C0007561|ceftriaxone|ceftriaxone
Drug|Organic Chemical|History of Present Illness|840,851|false|false|false|C0007561|ceftriaxone|ceftriaxone
Event|Event|History of Present Illness|840,851|false|false|false|||ceftriaxone
Drug|Antibiotic|History of Present Illness|852,863|false|false|false|C0055011|cefpodoxime|cefpodoxime
Drug|Organic Chemical|History of Present Illness|852,863|false|false|false|C0055011|cefpodoxime|cefpodoxime
Event|Event|History of Present Illness|852,863|false|false|false|||cefpodoxime
Event|Event|History of Present Illness|873,880|false|false|false|||treated
Drug|Hormone|History of Present Illness|894,904|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|History of Present Illness|894,904|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|History of Present Illness|894,904|false|false|false|C0032952|prednisone|prednisone
Event|Event|History of Present Illness|894,904|false|false|false|||prednisone
Event|Event|History of Present Illness|910,920|false|false|false|||discharged
Drug|Hormone|History of Present Illness|928,938|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|History of Present Illness|928,938|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|History of Present Illness|928,938|false|false|false|C0032952|prednisone|prednisone
Event|Event|History of Present Illness|939,944|false|false|false|||taper
Procedure|Health Care Activity|History of Present Illness|939,944|false|false|false|C0441640||taper
Finding|Finding|History of Present Illness|954,962|false|false|false|C0392756|Reduced|decrease
Finding|Intellectual Product|History of Present Illness|984,988|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|History of Present Illness|989,993|false|false|false|||stay
Procedure|Health Care Activity|History of Present Illness|1009,1013|false|false|false|C1315068|Pulmonary ventilator management|pulm
Event|Event|History of Present Illness|1014,1020|false|false|false|||follow
Finding|Functional Concept|History of Present Illness|1014,1020|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|History of Present Illness|1014,1020|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|History of Present Illness|1014,1023|false|false|false|C0589120|Follow-up status|follow up
Procedure|Health Care Activity|History of Present Illness|1014,1023|false|false|false|C1522577|follow-up|follow up
Event|Event|History of Present Illness|1039,1048|false|false|false|||counseled
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1055,1064|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|History of Present Illness|1055,1064|false|false|false|C2707265||pulmonary
Finding|Finding|History of Present Illness|1055,1064|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Event|Event|History of Present Illness|1065,1070|false|false|false|||rehab
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1065,1070|false|false|false|C0034991|Rehabilitation therapy|rehab
Event|Event|History of Present Illness|1075,1081|false|false|false|||follow
Event|Event|History of Present Illness|1108,1118|false|false|false|||discharged
Event|Event|History of Present Illness|1122,1124|false|false|false|||2L
Event|Event|History of Present Illness|1125,1137|false|false|false|||supplemental
Finding|Functional Concept|History of Present Illness|1125,1137|false|false|false|C2348609|Supplement|supplemental
Disorder|Disease or Syndrome|History of Present Illness|1160,1165|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Event|Event|History of Present Illness|1160,1165|false|false|false|||times
Drug|Organic Chemical|History of Present Illness|1170,1182|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|History of Present Illness|1170,1182|false|false|false|C0039771|theophylline|theophylline
Event|Event|History of Present Illness|1170,1182|false|false|false|||theophylline
Procedure|Laboratory Procedure|History of Present Illness|1170,1182|false|false|false|C0039773|Assay of theophylline|theophylline
Event|Event|History of Present Illness|1187,1196|false|false|false|||decreased
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|1209,1212|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1209,1212|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|History of Present Illness|1209,1212|false|false|false|C1530795|BID protein, human|BID
Event|Event|History of Present Illness|1209,1212|false|false|false|||BID
Finding|Gene or Genome|History of Present Illness|1209,1212|false|false|false|C1332410|BID gene|BID
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|1224,1227|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1224,1227|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|History of Present Illness|1224,1227|false|false|false|C1530795|BID protein, human|BID
Event|Event|History of Present Illness|1224,1227|false|false|false|||BID
Finding|Gene or Genome|History of Present Illness|1224,1227|false|false|false|C1332410|BID gene|BID
Disorder|Disease or Syndrome|History of Present Illness|1239,1243|false|false|false|C0004238|Atrial Fibrillation|afib
Event|Event|History of Present Illness|1239,1243|false|false|false|||afib
Lab|Laboratory or Test Result|History of Present Illness|1239,1243|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|afib
Event|Event|History of Present Illness|1249,1252|false|false|false|||RVR
Finding|Finding|History of Present Illness|1249,1252|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Finding|Gene or Genome|History of Present Illness|1249,1252|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Event|Event|History of Present Illness|1270,1274|false|false|false|||seen
Event|Event|History of Present Illness|1307,1314|false|false|false|||dyspnea
Finding|Finding|History of Present Illness|1307,1314|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|History of Present Illness|1307,1314|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Event|Event|History of Present Illness|1326,1330|false|false|false|||felt
Event|Event|History of Present Illness|1339,1351|false|false|false|||continuation
Disorder|Disease or Syndrome|History of Present Illness|1359,1363|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|History of Present Illness|1359,1363|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|History of Present Illness|1359,1363|false|false|false|||COPD
Finding|Gene or Genome|History of Present Illness|1359,1363|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|History of Present Illness|1364,1369|true|false|false|||flare
Finding|Finding|History of Present Illness|1364,1369|true|false|false|C1517205;C3540542|Exacerbation of cGVHD;Flare|flare
Finding|Sign or Symptom|History of Present Illness|1364,1369|true|false|false|C1517205;C3540542|Exacerbation of cGVHD;Flare|flare
Event|Event|History of Present Illness|1378,1385|true|false|false|||setting
Finding|Mental Process|History of Present Illness|1378,1385|true|false|false|C0542559|contextual factors|setting
Finding|Body Substance|History of Present Illness|1389,1396|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1389,1396|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1389,1396|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|1401,1407|true|false|false|||taking
Finding|Idea or Concept|History of Present Illness|1412,1416|true|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|History of Present Illness|1412,1416|true|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|History of Present Illness|1412,1416|true|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|History of Present Illness|1417,1428|true|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|History of Present Illness|1417,1428|true|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|History of Present Illness|1417,1428|true|false|false|||medications
Finding|Intellectual Product|History of Present Illness|1417,1428|true|false|false|C4284232|Medications|medications
Drug|Pharmacologic Substance|History of Present Illness|1445,1455|false|false|false|C2064916|nebulizers (medication)|nebulizers
Event|Event|History of Present Illness|1445,1455|false|false|false|||nebulizers
Event|Event|History of Present Illness|1460,1468|false|false|false|||improved
Event|Event|History of Present Illness|1478,1482|false|false|false|||DCed
Event|Event|History of Present Illness|1483,1487|false|false|false|||home
Finding|Idea or Concept|History of Present Illness|1483,1487|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|History of Present Illness|1483,1487|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|History of Present Illness|1483,1487|false|false|false|C1553498|home health encounter|home
Event|Event|History of Present Illness|1502,1512|false|false|false|||assistance
Finding|Social Behavior|History of Present Illness|1502,1512|false|false|false|C0018896|Helping Behavior|assistance
Attribute|Clinical Attribute|History of Present Illness|1518,1529|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|History of Present Illness|1518,1529|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|History of Present Illness|1518,1529|false|false|false|||medications
Finding|Intellectual Product|History of Present Illness|1518,1529|false|false|false|C4284232|Medications|medications
Event|Event|History of Present Illness|1535,1543|false|false|false|||declined
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1544,1553|true|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|History of Present Illness|1544,1553|true|false|false|C2707265||pulmonary
Finding|Finding|History of Present Illness|1544,1553|true|false|false|C4522268|Pulmonary (intended site)|pulmonary
Event|Event|History of Present Illness|1554,1559|true|false|false|||rehab
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1554,1559|true|false|false|C0034991|Rehabilitation therapy|rehab
Finding|Intellectual Product|History of Present Illness|1561,1569|true|false|false|C4695111|ADMIN.FACILITY|facility
Attribute|Clinical Attribute|History of Present Illness|1570,1581|true|false|false|C2926604||disposition
Event|Event|History of Present Illness|1570,1581|true|false|false|||disposition
Procedure|Health Care Activity|History of Present Illness|1570,1581|true|false|false|C0184758|Patient disposition|disposition
Finding|Idea or Concept|History of Present Illness|1597,1604|false|false|false|C1555582|Initial (abbreviation)|initial
Event|Event|History of Present Illness|1605,1611|false|false|false|||vitals
Event|Event|History of Present Illness|1617,1621|false|false|false|||Exam
Finding|Functional Concept|History of Present Illness|1617,1621|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|History of Present Illness|1617,1621|false|false|false|C0582103|Medical Examination|Exam
Event|Event|History of Present Illness|1622,1629|false|false|false|||notable
Finding|Gene or Genome|History of Present Illness|1648,1651|false|false|false|C0015373;C1421982|Extrasensory Perception;PTPRVP gene|esp
Finding|Mental Process|History of Present Illness|1648,1651|false|false|false|C0015373;C1421982|Extrasensory Perception;PTPRVP gene|esp
Event|Event|History of Present Illness|1652,1660|false|false|false|||wheezing
Finding|Sign or Symptom|History of Present Illness|1652,1660|false|false|false|C0043144|Wheezing|wheezing
Anatomy|Body Location or Region|History of Present Illness|1666,1676|false|false|false|C0521367|Oropharyngeal|oropharynx
Lab|Laboratory or Test Result|History of Present Illness|1681,1685|false|false|false|C0587081|Laboratory test finding|Labs
Event|Event|History of Present Illness|1686,1693|false|false|false|||notable
Anatomy|Cell|History of Present Illness|1702,1705|false|false|false|C0023516|Leukocytes|WBC
Event|Event|History of Present Illness|1715,1718|false|false|false|||neg
Finding|Finding|History of Present Illness|1715,1718|false|false|false|C5848551|Neg - answer|neg
Event|Event|History of Present Illness|1720,1723|false|false|false|||EKG
Finding|Intellectual Product|History of Present Illness|1720,1723|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|History of Present Illness|1720,1723|false|false|false|C1623258|Electrocardiography|EKG
Anatomy|Body Space or Junction|History of Present Illness|1727,1732|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|History of Present Illness|1727,1732|false|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|History of Present Illness|1727,1732|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|History of Present Illness|1727,1732|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Event|Event|History of Present Illness|1736,1743|false|false|false|||Imaging
Finding|Finding|History of Present Illness|1736,1743|false|false|false|C0740845|Imaging problem|Imaging
Procedure|Diagnostic Procedure|History of Present Illness|1736,1743|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|Imaging
Event|Event|History of Present Illness|1744,1751|false|false|false|||notable
Event|Event|History of Present Illness|1757,1760|true|false|false|||CXR
Procedure|Diagnostic Procedure|History of Present Illness|1757,1760|true|false|false|C0039985|Plain chest X-ray|CXR
Finding|Intellectual Product|History of Present Illness|1764,1769|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1770,1777|true|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|History of Present Illness|1770,1777|true|false|false|C1951340|Process Pharmacologic Substance|process
Event|Event|History of Present Illness|1770,1777|true|false|false|||process
Finding|Functional Concept|History of Present Illness|1770,1777|true|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|History of Present Illness|1770,1777|true|false|false|C1522240|Process|process
Drug|Organic Chemical|History of Present Illness|1792,1798|false|false|false|C0939692|DuoNeb|duoneb
Drug|Pharmacologic Substance|History of Present Illness|1792,1798|false|false|false|C0939692|DuoNeb|duoneb
Event|Event|History of Present Illness|1792,1798|false|false|false|||duoneb
Event|Event|History of Present Illness|1815,1820|false|false|false|||125mg
Drug|Organic Chemical|History of Present Illness|1822,1829|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|History of Present Illness|1822,1829|false|false|false|C0004057|aspirin|Aspirin
Drug|Antibiotic|History of Present Illness|1849,1861|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|History of Present Illness|1849,1861|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|History of Present Illness|1849,1861|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Event|Event|History of Present Illness|1862,1867|false|false|false|||500mg
Finding|Finding|History of Present Illness|1869,1878|false|false|false|C0857465|Peak flow|Peak flow
Event|Event|History of Present Illness|1874,1878|false|false|false|||flow
Phenomenon|Natural Phenomenon or Process|History of Present Illness|1874,1878|false|false|false|C0806140|Flow|flow
Drug|Biomedical or Dental Material|History of Present Illness|1884,1892|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|History of Present Illness|1884,1892|false|false|false|||baseline
Finding|Idea or Concept|History of Present Illness|1884,1892|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|History of Present Illness|1901,1909|false|false|false|||Symptoms
Finding|Functional Concept|History of Present Illness|1901,1909|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|Symptoms
Finding|Sign or Symptom|History of Present Illness|1901,1909|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|Symptoms
Finding|Intellectual Product|History of Present Illness|1911,1918|false|false|false|C0282416|Overall Publication Type|overall
Event|Event|History of Present Illness|1919,1927|false|false|false|||improved
Drug|Biomedical or Dental Material|History of Present Illness|1934,1938|false|false|false|C1300458|Nebulizer solution|nebs
Event|Event|History of Present Illness|1934,1938|false|false|false|||nebs
Event|Event|History of Present Illness|1959,1967|false|false|false|||transfer
Finding|Functional Concept|History of Present Illness|1959,1967|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|History of Present Illness|1959,1967|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|History of Present Illness|1959,1967|false|false|false|C4706767|Transfer (immobility management)|transfer
Event|Activity|History of Present Illness|1999,2006|false|false|false|C1706079||arrival
Event|Event|History of Present Illness|1999,2006|false|false|false|||arrival
Finding|Functional Concept|History of Present Illness|1999,2006|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Anatomy|Anatomical Structure|History of Present Illness|2014,2019|false|false|false|C3714591|Floor (anatomic)|floor
Event|Event|History of Present Illness|2024,2031|false|false|false|||reports
Event|Event|History of Present Illness|2032,2039|false|false|false|||feeling
Finding|Finding|History of Present Illness|2040,2044|false|false|false|C4281574|Much|much
Event|Event|History of Present Illness|2045,2053|false|false|false|||improved
Finding|Finding|History of Present Illness|2045,2053|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Finding|Intellectual Product|History of Present Illness|2045,2053|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Event|Event|History of Present Illness|2067,2075|false|false|false|||wheezing
Finding|Sign or Symptom|History of Present Illness|2067,2075|false|false|false|C0043144|Wheezing|wheezing
Event|Event|Review of Systems|2088,2094|true|false|false|||fevers
Finding|Sign or Symptom|Review of Systems|2088,2094|true|false|false|C0015967|Fever|fevers
Event|Event|Review of Systems|2096,2102|true|false|false|||chills
Finding|Sign or Symptom|Review of Systems|2096,2102|true|false|false|C0085593|Chills|chills
Finding|Sign or Symptom|Review of Systems|2104,2116|true|false|false|C0028081|Night sweats|night sweats
Event|Event|Review of Systems|2110,2116|true|false|false|||sweats
Finding|Body Substance|Review of Systems|2110,2116|true|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Finding|Finding|Review of Systems|2110,2116|true|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Attribute|Clinical Attribute|Review of Systems|2121,2127|false|false|false|C0944911||weight
Event|Event|Review of Systems|2121,2127|false|false|false|||weight
Finding|Finding|Review of Systems|2121,2127|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|Review of Systems|2121,2127|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|Review of Systems|2121,2127|false|false|false|C1305866|Weighing patient|weight
Finding|Finding|Review of Systems|2121,2135|true|false|false|C0005911|Body Weight Changes|weight changes
Event|Event|Review of Systems|2128,2135|false|false|false|||changes
Finding|Functional Concept|Review of Systems|2128,2135|true|false|false|C0392747|Changing|changes
Event|Event|Review of Systems|2140,2147|true|false|false|||changes
Finding|Functional Concept|Review of Systems|2140,2147|true|false|false|C0392747|Changing|changes
Attribute|Clinical Attribute|Review of Systems|2152,2158|true|false|false|C2707266||vision
Event|Event|Review of Systems|2152,2158|true|false|false|||vision
Finding|Organism Function|Review of Systems|2152,2158|true|false|false|C0042789|Vision|vision
Event|Event|Review of Systems|2162,2169|true|false|false|||hearing
Finding|Finding|Review of Systems|2162,2169|true|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|hearing
Finding|Physiologic Function|Review of Systems|2162,2169|true|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|hearing
Event|Event|Review of Systems|2174,2181|true|false|false|||changes
Finding|Functional Concept|Review of Systems|2174,2181|true|false|false|C0392747|Changing|changes
Drug|Organic Chemical|Review of Systems|2185,2192|true|false|false|C4319618|Balance (substance)|balance
Drug|Pharmacologic Substance|Review of Systems|2185,2192|true|false|false|C4319618|Balance (substance)|balance
Event|Event|Review of Systems|2185,2192|true|false|false|||balance
Finding|Finding|Review of Systems|2185,2192|true|false|false|C0014653;C0560184|Ability to balance;Equilibrium|balance
Finding|Organism Function|Review of Systems|2185,2192|true|false|false|C0014653;C0560184|Ability to balance;Equilibrium|balance
Procedure|Diagnostic Procedure|Review of Systems|2185,2192|true|false|false|C2174421|examination of balance|balance
Drug|Organic Chemical|Review of Systems|2197,2202|true|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|Review of Systems|2197,2202|true|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|Review of Systems|2197,2202|true|false|false|||cough
Finding|Sign or Symptom|Review of Systems|2197,2202|true|false|false|C0010200|Coughing|cough
Event|Event|Review of Systems|2204,2206|true|false|false|||no
Event|Event|Review of Systems|2208,2217|true|false|false|||shortness
Attribute|Clinical Attribute|Review of Systems|2208,2227|true|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|Review of Systems|2208,2227|true|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|Review of Systems|2221,2227|true|false|false|C0225386|Breath|breath
Event|Event|Review of Systems|2232,2239|true|false|false|||dyspnea
Finding|Finding|Review of Systems|2232,2239|true|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|Review of Systems|2232,2239|true|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|Review of Systems|2232,2251|true|false|false|C0231807|Dyspnea on exertion|dyspnea on exertion
Event|Event|Review of Systems|2243,2251|true|false|false|||exertion
Finding|Organism Function|Review of Systems|2243,2251|true|false|false|C0015264|Exertion|exertion
Anatomy|Body Location or Region|Review of Systems|2256,2261|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Review of Systems|2256,2261|true|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Review of Systems|2256,2266|true|false|false|C2926613||chest pain
Finding|Sign or Symptom|Review of Systems|2256,2266|true|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Review of Systems|2262,2266|true|false|false|C2598155||pain
Event|Event|Review of Systems|2262,2266|true|false|false|||pain
Finding|Functional Concept|Review of Systems|2262,2266|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Review of Systems|2262,2266|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Review of Systems|2271,2283|true|false|false|||palpitations
Finding|Finding|Review of Systems|2271,2283|true|false|false|C0030252|Palpitations|palpitations
Attribute|Clinical Attribute|Review of Systems|2288,2294|true|false|false|C4255480||nausea
Event|Event|Review of Systems|2288,2294|true|false|false|||nausea
Finding|Sign or Symptom|Review of Systems|2288,2294|true|false|false|C0027497|Nausea|nausea
Finding|Finding|Review of Systems|2288,2306|true|false|false|C3843946|Nausea or vomiting|nausea or vomiting
Event|Event|Review of Systems|2298,2306|true|false|false|||vomiting
Finding|Sign or Symptom|Review of Systems|2298,2306|true|false|false|C0042963|Vomiting|vomiting
Event|Event|Review of Systems|2311,2319|true|false|false|||diarrhea
Finding|Finding|Review of Systems|2311,2319|true|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|Review of Systems|2311,2319|true|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Event|Event|Review of Systems|2324,2336|true|false|false|||constipation
Finding|Sign or Symptom|Review of Systems|2324,2336|true|false|false|C0009806|Constipation|constipation
Event|Event|Review of Systems|2341,2348|true|false|false|||dysuria
Finding|Sign or Symptom|Review of Systems|2341,2348|true|false|false|C0013428|Dysuria|dysuria
Disorder|Disease or Syndrome|Review of Systems|2352,2361|true|false|false|C0018965|Hematuria|hematuria
Event|Event|Review of Systems|2352,2361|true|false|false|||hematuria
Disorder|Disease or Syndrome|Review of Systems|2366,2378|true|false|false|C0018932|Hematochezia|hematochezia
Event|Event|Review of Systems|2366,2378|true|false|false|||hematochezia
Finding|Sign or Symptom|Review of Systems|2366,2378|true|false|false|C1321898|Blood in stool|hematochezia
Event|Event|Review of Systems|2384,2390|true|false|false|||melena
Finding|Pathologic Function|Review of Systems|2384,2390|true|false|false|C0025222|Melena|melena
Event|Event|Review of Systems|2395,2403|true|false|false|||numbness
Finding|Finding|Review of Systems|2395,2403|true|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|Review of Systems|2395,2403|true|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Event|Event|Review of Systems|2407,2415|true|false|false|||weakness
Finding|Sign or Symptom|Review of Systems|2407,2415|true|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Event|Event|Review of Systems|2426,2434|true|false|false|||deficits
Disorder|Disease or Syndrome|Past Medical History|2463,2469|false|false|false|C0004096|Asthma|ASTHMA
Event|Event|Past Medical History|2463,2469|false|false|false|||ASTHMA
Disorder|Disease or Syndrome|Past Medical History|2470,2474|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Past Medical History|2470,2474|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Past Medical History|2470,2474|false|false|false|||COPD
Finding|Gene or Genome|Past Medical History|2470,2474|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Finding|Past Medical History|2478,2486|false|false|false|C0741302|atypia morphology|ATYPICAL
Finding|Sign or Symptom|Past Medical History|2478,2497|false|false|false|C0262384|Atypical chest pain|ATYPICAL CHEST PAIN
Anatomy|Body Location or Region|Past Medical History|2487,2492|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|CHEST
Finding|Finding|Past Medical History|2487,2492|false|false|false|C0741025|Chest problem|CHEST
Attribute|Clinical Attribute|Past Medical History|2487,2497|false|false|false|C2926613||CHEST PAIN
Finding|Sign or Symptom|Past Medical History|2487,2497|false|false|false|C0008031|Chest Pain|CHEST PAIN
Attribute|Clinical Attribute|Past Medical History|2493,2497|false|true|false|C2598155||PAIN
Event|Event|Past Medical History|2493,2497|false|false|false|||PAIN
Finding|Functional Concept|Past Medical History|2493,2497|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|PAIN
Finding|Sign or Symptom|Past Medical History|2493,2497|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|PAIN
Anatomy|Body Location or Region|Past Medical History|2501,2509|false|false|false|C0027530|Neck|CERVICAL
Disorder|Disease or Syndrome|Past Medical History|2501,2521|false|false|false|C0263884|Cervical radiculitis|CERVICAL RADICULITIS
Disorder|Disease or Syndrome|Past Medical History|2510,2521|false|false|false|C0034544|Radiculitis|RADICULITIS
Event|Event|Past Medical History|2510,2521|false|false|false|||RADICULITIS
Anatomy|Body Location or Region|Past Medical History|2525,2533|false|false|false|C0027530|Neck|CERVICAL
Disorder|Disease or Syndrome|Past Medical History|2525,2545|false|false|false|C0158241;C1384641|Cervical spondylosis;Cervical spondylosis without myelopathy|CERVICAL SPONDYLOSIS
Disorder|Disease or Syndrome|Past Medical History|2534,2545|false|false|false|C0038019|Spondylosis|SPONDYLOSIS
Event|Event|Past Medical History|2534,2545|false|false|false|||SPONDYLOSIS
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2549,2557|false|false|false|C0018787|Heart|CORONARY
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2549,2564|false|false|false|C0205042|Coronary artery|CORONARY ARTERY
Disorder|Disease or Syndrome|Past Medical History|2549,2572|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|CORONARY ARTERY DISEASE
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2558,2564|false|false|false|C0003842;C0226004|Arterial system;Arteries|ARTERY
Anatomy|Body System|Past Medical History|2558,2564|false|false|false|C0003842;C0226004|Arterial system;Arteries|ARTERY
Disorder|Disease or Syndrome|Past Medical History|2558,2572|false|false|false|C0852949|Arteriopathic disease|ARTERY DISEASE
Disorder|Disease or Syndrome|Past Medical History|2565,2572|false|false|false|C0012634|Disease|DISEASE
Event|Event|Past Medical History|2565,2572|false|false|false|||DISEASE
Finding|Sign or Symptom|Past Medical History|2576,2584|false|false|false|C0018681|Headache|HEADACHE
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2588,2591|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|HIP
Drug|Amino Acid, Peptide, or Protein|Past Medical History|2588,2591|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|HIP
Drug|Biologically Active Substance|Past Medical History|2588,2591|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|HIP
Drug|Pharmacologic Substance|Past Medical History|2588,2591|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|HIP
Event|Event|Past Medical History|2588,2591|false|false|false|||HIP
Finding|Gene or Genome|Past Medical History|2588,2591|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|HIP
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2588,2591|false|false|false|C1292890|Procedure on hip|HIP
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2588,2603|false|false|false|C0392806|Prosthetic arthroplasty of hip (procedure)|HIP REPLACEMENT
Event|Event|Past Medical History|2592,2603|false|false|false|||REPLACEMENT
Finding|Functional Concept|Past Medical History|2592,2603|false|false|false|C0559956|Replacement|REPLACEMENT
Procedure|Health Care Activity|Past Medical History|2592,2603|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|REPLACEMENT
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2592,2603|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|REPLACEMENT
Disorder|Disease or Syndrome|Past Medical History|2607,2621|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|HYPERLIPIDEMIA
Event|Event|Past Medical History|2607,2621|false|false|false|||HYPERLIPIDEMIA
Finding|Finding|Past Medical History|2607,2621|false|false|false|C0428465|Serum lipids high (finding)|HYPERLIPIDEMIA
Disorder|Disease or Syndrome|Past Medical History|2625,2637|false|false|false|C0020538|Hypertensive disease|HYPERTENSION
Event|Event|Past Medical History|2625,2637|false|false|false|||HYPERTENSION
Disorder|Disease or Syndrome|Past Medical History|2641,2655|false|false|false|C0029408|Degenerative polyarthritis|OSTEOARTHRITIS
Event|Event|Past Medical History|2641,2655|false|false|false|||OSTEOARTHRITIS
Disorder|Disease or Syndrome|Past Medical History|2659,2665|false|false|false|C0019340;C0854331|Herpes simplex dermatitis|HERPES
Disorder|Disease or Syndrome|Past Medical History|2659,2672|false|false|false|C0019360;C0042338|Herpes zoster (disorder);herpesvirus 3, human|HERPES ZOSTER
Disorder|Virus|Past Medical History|2659,2672|false|false|false|C0019360;C0042338|Herpes zoster (disorder);herpesvirus 3, human|HERPES ZOSTER
Disorder|Disease or Syndrome|Past Medical History|2666,2672|false|false|false|C0019360|Herpes zoster (disorder)|ZOSTER
Event|Event|Past Medical History|2666,2672|false|false|false|||ZOSTER
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2676,2682|false|false|false|C0018792|Heart Atrium|ATRIAL
Attribute|Clinical Attribute|Past Medical History|2676,2695|false|false|false|C2926591||ATRIAL FIBRILLATION
Disorder|Disease or Syndrome|Past Medical History|2676,2695|false|false|false|C0004238|Atrial Fibrillation|ATRIAL FIBRILLATION
Lab|Laboratory or Test Result|Past Medical History|2676,2695|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|ATRIAL FIBRILLATION
Disorder|Disease or Syndrome|Past Medical History|2683,2695|false|false|false|C0232197|Fibrillation|FIBRILLATION
Event|Event|Past Medical History|2683,2695|false|false|false|||FIBRILLATION
Disorder|Mental or Behavioral Dysfunction|Past Medical History|2699,2706|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|ANXIETY
Event|Event|Past Medical History|2699,2706|false|false|false|||ANXIETY
Finding|Sign or Symptom|Past Medical History|2699,2706|false|false|false|C0860603|Anxiety symptoms|ANXIETY
Finding|Intellectual Product|Past Medical History|2710,2726|false|false|false|C1314977|Gastrointestinal attachment|GASTROINTESTINAL
Finding|Pathologic Function|Past Medical History|2710,2735|false|false|false|C0017181|Gastrointestinal Hemorrhage|GASTROINTESTINAL BLEEDING
Finding|Pathologic Function|Past Medical History|2727,2735|false|false|false|C0019080|Hemorrhage|BLEEDING
Disorder|Disease or Syndrome|Past Medical History|2739,2753|false|false|false|C0029408|Degenerative polyarthritis|OSTEOARTHRITIS
Event|Event|Past Medical History|2739,2753|false|false|false|||OSTEOARTHRITIS
Finding|Functional Concept|Past Medical History|2757,2772|false|false|false|C0333482|atherosclerotic|ATHEROSCLEROTIC
Disorder|Disease or Syndrome|Past Medical History|2757,2795|false|false|false|C0004153|Atherosclerosis|ATHEROSCLEROTIC CARDIOVASCULAR DISEASE
Anatomy|Body System|Past Medical History|2773,2787|false|false|false|C0007226;C3887460|Cardiovascular;Cardiovascular system|CARDIOVASCULAR
Disorder|Disease or Syndrome|Past Medical History|2773,2795|false|false|false|C0007222|Cardiovascular Diseases|CARDIOVASCULAR DISEASE
Disorder|Disease or Syndrome|Past Medical History|2788,2795|false|false|false|C0012634|Disease|DISEASE
Event|Event|Past Medical History|2788,2795|false|false|false|||DISEASE
Disorder|Disease or Syndrome|Past Medical History|2799,2826|false|false|false|C0085096|Peripheral Vascular Diseases|PERIPHERAL VASCULAR DISEASE
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2810,2818|false|false|false|C0005847|Blood Vessel|VASCULAR
Disorder|Disease or Syndrome|Past Medical History|2810,2826|false|false|false|C0042373|Vascular Diseases|VASCULAR DISEASE
Disorder|Disease or Syndrome|Past Medical History|2819,2826|false|false|false|C0012634|Disease|DISEASE
Event|Event|Past Medical History|2819,2826|false|false|false|||DISEASE
Finding|Idea or Concept|Family Medical History|2865,2871|false|false|false|C1546508|Relationship - Mother|Mother
Disorder|Disease or Syndrome|Family Medical History|2878,2881|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|Family Medical History|2878,2881|false|false|false|||HTN
Finding|Conceptual Entity|Family Medical History|2884,2890|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|Family Medical History|2884,2890|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Event|Event|Family Medical History|2901,2908|false|false|false|||Brother
Finding|Conceptual Entity|Family Medical History|2901,2908|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Idea or Concept|Family Medical History|2901,2908|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Event|Event|Family Medical History|2916,2923|false|false|false|||Brother
Finding|Conceptual Entity|Family Medical History|2916,2923|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Idea or Concept|Family Medical History|2916,2923|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Event|Event|Family Medical History|2932,2940|false|false|false|||Physical
Finding|Finding|Family Medical History|2932,2940|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|Family Medical History|2932,2940|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|Family Medical History|2932,2940|false|false|false|C0031809|Physical Examination|Physical
Event|Event|Family Medical History|2946,2955|false|false|false|||Admission
Procedure|Health Care Activity|Family Medical History|2946,2955|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Event|Event|Family Medical History|2988,2995|false|false|false|||General
Finding|Classification|Family Medical History|2988,2995|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|Family Medical History|2988,2995|false|false|false|C3812897|General medical service|General
Attribute|Clinical Attribute|Family Medical History|2997,3002|true|false|false|C5890168||Alert
Drug|Organic Chemical|Family Medical History|2997,3002|true|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Family Medical History|2997,3002|true|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Family Medical History|2997,3002|true|false|false|||Alert
Finding|Finding|Family Medical History|2997,3002|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Family Medical History|2997,3002|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Family Medical History|2997,3002|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Family Medical History|3004,3012|true|false|false|||oriented
Finding|Intellectual Product|Family Medical History|3017,3022|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|Family Medical History|3023,3031|true|false|false|||distress
Finding|Finding|Family Medical History|3023,3031|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|Family Medical History|3023,3031|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Event|Event|Family Medical History|3033,3040|true|false|false|||appears
Drug|Amino Acid, Peptide, or Protein|Family Medical History|3046,3050|true|true|false|C1366910|Calmodulin 1|calm
Drug|Biologically Active Substance|Family Medical History|3046,3050|true|true|false|C1366910|Calmodulin 1|calm
Event|Event|Family Medical History|3046,3050|true|false|false|||calm
Finding|Gene or Genome|Family Medical History|3046,3050|true|true|false|C0522165;C1423112;C1423544;C2827449;C5551289|Feeling calm;PICALM gene;PICALM wt Allele;SNAP91 gene;SNAP91 wt Allele|calm
Finding|Mental Process|Family Medical History|3046,3050|true|true|false|C0522165;C1423112;C1423544;C2827449;C5551289|Feeling calm;PICALM gene;PICALM wt Allele;SNAP91 gene;SNAP91 wt Allele|calm
Procedure|Therapeutic or Preventive Procedure|Family Medical History|3046,3050|true|true|false|C5552882|Cancer and Living Meaningfully Therapy|calm
Event|Event|Family Medical History|3060,3064|false|false|false|||talk
Event|Event|Family Medical History|3073,3082|false|false|false|||sentences
Finding|Intellectual Product|Family Medical History|3073,3082|false|false|true|C0876929|Sentence|sentences
Anatomy|Body Location or Region|Family Medical History|3084,3089|false|false|false|C1512338|HEENT|HEENT
Event|Event|Family Medical History|3099,3108|false|false|false|||anicteric
Finding|Finding|Family Medical History|3099,3108|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3110,3113|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|Family Medical History|3110,3113|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Location or Region|Family Medical History|3115,3125|false|false|false|C0521367|Oropharyngeal|oropharynx
Event|Event|Family Medical History|3126,3131|false|false|false|||clear
Finding|Idea or Concept|Family Medical History|3126,3131|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Location or Region|Family Medical History|3134,3138|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|Family Medical History|3134,3138|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|Family Medical History|3134,3138|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|Family Medical History|3140,3146|true|false|false|||supple
Finding|Functional Concept|Family Medical History|3140,3146|true|false|false|C0332254|Supple|supple
Event|Event|Family Medical History|3148,3151|true|false|false|||JVP
Finding|Finding|Family Medical History|3148,3151|true|false|false|C0428897|Jugular venous pressure|JVP
Event|Event|Family Medical History|3156,3164|true|false|false|||elevated
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3169,3172|true|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|Family Medical History|3169,3172|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|Family Medical History|3169,3172|true|false|false|||LAD
Finding|Gene or Genome|Family Medical History|3169,3172|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3175,3180|true|false|false|C0024109|Lung|Lungs
Event|Event|Family Medical History|3192,3200|false|false|false|||wheezing
Finding|Sign or Symptom|Family Medical History|3192,3200|false|false|false|C0043144|Wheezing|wheezing
Finding|Organ or Tissue Function|Family Medical History|3218,3226|false|false|false|C0039155|Systole|systolic
Finding|Finding|Family Medical History|3218,3233|true|false|false|C0232257|Systolic Murmurs|systolic murmur
Event|Event|Family Medical History|3227,3233|true|false|false|||murmur
Finding|Finding|Family Medical History|3227,3233|true|false|false|C0018808|Heart murmur|murmur
Event|Event|Family Medical History|3249,3252|true|false|false|||MRG
Finding|Gene or Genome|Family Medical History|3249,3252|true|false|false|C1422304|MAS1L gene|MRG
Anatomy|Body Location or Region|Family Medical History|3255,3262|true|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|Family Medical History|3255,3262|true|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Event|Event|Family Medical History|3255,3262|true|false|false|||Abdomen
Finding|Finding|Family Medical History|3255,3262|true|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|Family Medical History|3264,3268|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|Family Medical History|3264,3268|false|false|false|||soft
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3276,3281|true|false|false|C0021853|Intestines|bowel
Finding|Finding|Family Medical History|3276,3288|true|false|false|C0232693|Bowel sounds|bowel sounds
Event|Event|Family Medical History|3282,3288|true|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|Family Medical History|3282,3288|true|false|false|C0037709||sounds
Finding|Finding|Family Medical History|3289,3296|true|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|Family Medical History|3289,3296|true|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Sign or Symptom|Family Medical History|3301,3319|true|false|false|C0234246|Rebound tenderness|rebound tenderness
Event|Event|Family Medical History|3309,3319|true|false|false|||tenderness
Finding|Mental Process|Family Medical History|3309,3319|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|Family Medical History|3309,3319|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Event|Family Medical History|3324,3332|true|false|false|||guarding
Finding|Finding|Family Medical History|3324,3332|true|false|false|C0427198|Protective muscle spasm|guarding
Event|Event|Family Medical History|3337,3349|true|false|false|||organomegaly
Finding|Finding|Family Medical History|3337,3349|true|false|false|C4054315|Organomegaly|organomegaly
Event|Event|Family Medical History|3359,3364|true|false|false|||foley
Disorder|Congenital Abnormality|Family Medical History|3367,3370|true|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|Family Medical History|3367,3370|true|false|false|||Ext
Finding|Gene or Genome|Family Medical History|3367,3370|true|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|Family Medical History|3372,3376|false|false|false|||warm
Finding|Finding|Family Medical History|3372,3376|false|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|Family Medical History|3372,3376|false|false|false|C0687712|warming process|warm
Finding|Finding|Family Medical History|3378,3382|true|false|false|C5575035|Well (answer to question)|well
Event|Event|Family Medical History|3383,3391|true|false|false|||perfused
Drug|Food|Family Medical History|3396,3402|true|false|false|C5890763||pulses
Event|Event|Family Medical History|3396,3402|true|false|false|||pulses
Finding|Physiologic Function|Family Medical History|3396,3402|true|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|Family Medical History|3396,3402|true|false|false|C0034107|Pulse taking|pulses
Disorder|Anatomical Abnormality|Family Medical History|3407,3415|true|false|false|C0149651|Clubbing|clubbing
Event|Event|Family Medical History|3407,3415|true|false|false|||clubbing
Event|Event|Family Medical History|3417,3425|true|false|false|||cyanosis
Finding|Sign or Symptom|Family Medical History|3417,3425|true|false|false|C0010520|Cyanosis|cyanosis
Attribute|Clinical Attribute|Family Medical History|3431,3436|false|false|false|C1717255||edema
Event|Event|Family Medical History|3431,3436|false|false|false|||edema
Finding|Pathologic Function|Family Medical History|3431,3436|false|false|false|C0013604|Edema|edema
Finding|Gene or Genome|Family Medical History|3448,3451|true|false|false|C1539110|CNDP2 gene|CN2
Event|Event|Family Medical History|3455,3461|true|false|false|||intact
Finding|Finding|Family Medical History|3455,3461|true|false|false|C1554187|Gender Status - Intact|intact
Event|Event|Family Medical History|3472,3480|true|false|false|||deficits
Event|Event|Family Medical History|3531,3538|false|false|false|||General
Finding|Classification|Family Medical History|3531,3538|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|Family Medical History|3531,3538|false|false|false|C3812897|General medical service|General
Attribute|Clinical Attribute|Family Medical History|3540,3545|true|false|false|C5890168||Alert
Drug|Organic Chemical|Family Medical History|3540,3545|true|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Family Medical History|3540,3545|true|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Family Medical History|3540,3545|true|false|false|||Alert
Finding|Finding|Family Medical History|3540,3545|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Family Medical History|3540,3545|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Family Medical History|3540,3545|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Family Medical History|3547,3555|true|false|false|||oriented
Finding|Intellectual Product|Family Medical History|3560,3565|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|Family Medical History|3566,3574|true|false|false|||distress
Finding|Finding|Family Medical History|3566,3574|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|Family Medical History|3566,3574|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Event|Event|Family Medical History|3576,3583|true|false|false|||appears
Drug|Amino Acid, Peptide, or Protein|Family Medical History|3589,3593|true|true|false|C1366910|Calmodulin 1|calm
Drug|Biologically Active Substance|Family Medical History|3589,3593|true|true|false|C1366910|Calmodulin 1|calm
Event|Event|Family Medical History|3589,3593|true|false|false|||calm
Finding|Gene or Genome|Family Medical History|3589,3593|true|true|false|C0522165;C1423112;C1423544;C2827449;C5551289|Feeling calm;PICALM gene;PICALM wt Allele;SNAP91 gene;SNAP91 wt Allele|calm
Finding|Mental Process|Family Medical History|3589,3593|true|true|false|C0522165;C1423112;C1423544;C2827449;C5551289|Feeling calm;PICALM gene;PICALM wt Allele;SNAP91 gene;SNAP91 wt Allele|calm
Procedure|Therapeutic or Preventive Procedure|Family Medical History|3589,3593|true|true|false|C5552882|Cancer and Living Meaningfully Therapy|calm
Event|Event|Family Medical History|3603,3607|false|false|false|||talk
Event|Event|Family Medical History|3616,3625|false|false|false|||sentences
Finding|Intellectual Product|Family Medical History|3616,3625|false|false|true|C0876929|Sentence|sentences
Anatomy|Body Location or Region|Family Medical History|3627,3632|false|false|false|C1512338|HEENT|HEENT
Event|Event|Family Medical History|3642,3651|false|false|false|||anicteric
Finding|Finding|Family Medical History|3642,3651|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3653,3656|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|Family Medical History|3653,3656|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Location or Region|Family Medical History|3658,3668|false|false|false|C0521367|Oropharyngeal|oropharynx
Event|Event|Family Medical History|3669,3674|false|false|false|||clear
Finding|Idea or Concept|Family Medical History|3669,3674|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Location or Region|Family Medical History|3677,3681|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|Family Medical History|3677,3681|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|Family Medical History|3677,3681|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|Family Medical History|3683,3689|true|false|false|||supple
Finding|Functional Concept|Family Medical History|3683,3689|true|false|false|C0332254|Supple|supple
Event|Event|Family Medical History|3691,3694|true|false|false|||JVP
Finding|Finding|Family Medical History|3691,3694|true|false|false|C0428897|Jugular venous pressure|JVP
Event|Event|Family Medical History|3699,3707|true|false|false|||elevated
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3712,3715|true|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|Family Medical History|3712,3715|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|Family Medical History|3712,3715|true|false|false|||LAD
Finding|Gene or Genome|Family Medical History|3712,3715|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3718,3723|true|false|false|C0024109|Lung|Lungs
Event|Event|Family Medical History|3735,3743|false|false|false|||wheezing
Finding|Sign or Symptom|Family Medical History|3735,3743|false|false|false|C0043144|Wheezing|wheezing
Finding|Organ or Tissue Function|Family Medical History|3761,3769|false|false|false|C0039155|Systole|systolic
Finding|Finding|Family Medical History|3761,3776|true|false|false|C0232257|Systolic Murmurs|systolic murmur
Event|Event|Family Medical History|3770,3776|true|false|false|||murmur
Finding|Finding|Family Medical History|3770,3776|true|false|false|C0018808|Heart murmur|murmur
Event|Event|Family Medical History|3792,3795|true|false|false|||MRG
Finding|Gene or Genome|Family Medical History|3792,3795|true|false|false|C1422304|MAS1L gene|MRG
Anatomy|Body Location or Region|Family Medical History|3798,3805|true|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|Family Medical History|3798,3805|true|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Event|Event|Family Medical History|3798,3805|true|false|false|||Abdomen
Finding|Finding|Family Medical History|3798,3805|true|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|Family Medical History|3807,3811|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|Family Medical History|3807,3811|false|false|false|||soft
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3819,3824|true|false|false|C0021853|Intestines|bowel
Finding|Finding|Family Medical History|3819,3831|true|false|false|C0232693|Bowel sounds|bowel sounds
Event|Event|Family Medical History|3825,3831|true|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|Family Medical History|3825,3831|true|false|false|C0037709||sounds
Finding|Finding|Family Medical History|3832,3839|true|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|Family Medical History|3832,3839|true|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Sign or Symptom|Family Medical History|3844,3862|true|false|false|C0234246|Rebound tenderness|rebound tenderness
Event|Event|Family Medical History|3852,3862|true|false|false|||tenderness
Finding|Mental Process|Family Medical History|3852,3862|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|Family Medical History|3852,3862|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Event|Family Medical History|3867,3875|true|false|false|||guarding
Finding|Finding|Family Medical History|3867,3875|true|false|false|C0427198|Protective muscle spasm|guarding
Event|Event|Family Medical History|3880,3892|true|false|false|||organomegaly
Finding|Finding|Family Medical History|3880,3892|true|false|false|C4054315|Organomegaly|organomegaly
Event|Event|Family Medical History|3902,3907|true|false|false|||foley
Disorder|Congenital Abnormality|Family Medical History|3910,3913|true|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|Family Medical History|3910,3913|true|false|false|||Ext
Finding|Gene or Genome|Family Medical History|3910,3913|true|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|Family Medical History|3915,3919|false|false|false|||warm
Finding|Finding|Family Medical History|3915,3919|false|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|Family Medical History|3915,3919|false|false|false|C0687712|warming process|warm
Finding|Finding|Family Medical History|3921,3925|true|false|false|C5575035|Well (answer to question)|well
Event|Event|Family Medical History|3926,3934|true|false|false|||perfused
Drug|Food|Family Medical History|3939,3945|true|false|false|C5890763||pulses
Event|Event|Family Medical History|3939,3945|true|false|false|||pulses
Finding|Physiologic Function|Family Medical History|3939,3945|true|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|Family Medical History|3939,3945|true|false|false|C0034107|Pulse taking|pulses
Disorder|Anatomical Abnormality|Family Medical History|3950,3958|true|false|false|C0149651|Clubbing|clubbing
Event|Event|Family Medical History|3950,3958|true|false|false|||clubbing
Event|Event|Family Medical History|3960,3968|true|false|false|||cyanosis
Finding|Sign or Symptom|Family Medical History|3960,3968|true|false|false|C0010520|Cyanosis|cyanosis
Attribute|Clinical Attribute|Family Medical History|3974,3979|false|false|false|C1717255||edema
Event|Event|Family Medical History|3974,3979|false|false|false|||edema
Finding|Pathologic Function|Family Medical History|3974,3979|false|false|false|C0013604|Edema|edema
Finding|Gene or Genome|Family Medical History|3991,3994|true|false|false|C1539110|CNDP2 gene|CN2
Event|Event|Family Medical History|3998,4004|true|false|false|||intact
Finding|Finding|Family Medical History|3998,4004|true|false|false|C1554187|Gender Status - Intact|intact
Event|Event|Family Medical History|4015,4023|true|false|false|||deficits
Event|Event|Family Medical History|4045,4054|false|false|false|||Admission
Procedure|Health Care Activity|Family Medical History|4045,4054|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Disorder|Disease or Syndrome|Family Medical History|4068,4073|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|4068,4073|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|4068,4073|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|Family Medical History|4074,4077|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|Family Medical History|4082,4085|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|Family Medical History|4082,4085|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|Family Medical History|4082,4085|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|Family Medical History|4091,4094|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Family Medical History|4091,4094|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|Family Medical History|4091,4094|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Family Medical History|4091,4094|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|Family Medical History|4101,4104|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|Family Medical History|4101,4104|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|Family Medical History|4111,4114|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|Family Medical History|4111,4114|false|false|false|||MCV
Lab|Laboratory or Test Result|Family Medical History|4111,4114|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|Family Medical History|4111,4114|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|Family Medical History|4111,4114|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|Family Medical History|4119,4122|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|Family Medical History|4119,4122|false|false|false|C0600370|methacholine|MCH
Event|Event|Family Medical History|4119,4122|false|false|false|||MCH
Finding|Gene or Genome|Family Medical History|4119,4122|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|Family Medical History|4119,4122|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|Family Medical History|4119,4122|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|Family Medical History|4129,4133|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|Family Medical History|4162,4165|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|Family Medical History|4182,4187|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|4182,4187|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|4182,4187|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Body Substance|Family Medical History|4200,4206|false|false|false|C0024202|Lymph|Lymphs
Drug|Antibiotic|Family Medical History|4212,4217|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|Family Medical History|4212,4217|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|Family Medical History|4212,4217|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|Family Medical History|4224,4227|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Event|Event|Family Medical History|4224,4227|false|false|false|||Eos
Finding|Gene or Genome|Family Medical History|4224,4227|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|Family Medical History|4330,4335|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|4330,4335|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|4330,4335|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|Family Medical History|4340,4343|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|Family Medical History|4340,4343|false|false|false|||PTT
Procedure|Laboratory Procedure|Family Medical History|4340,4343|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|Family Medical History|4365,4370|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|4365,4370|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|4365,4370|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|Family Medical History|4365,4378|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|Family Medical History|4365,4378|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|Family Medical History|4365,4378|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|Family Medical History|4371,4378|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|Family Medical History|4371,4378|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|Family Medical History|4371,4378|false|false|false|C0017725|glucose|Glucose
Event|Event|Family Medical History|4371,4378|false|false|false|||Glucose
Lab|Laboratory or Test Result|Family Medical History|4371,4378|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|Family Medical History|4371,4378|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|Family Medical History|4424,4428|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|Family Medical History|4424,4428|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|Family Medical History|4424,4428|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|Family Medical History|4453,4458|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|4453,4458|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|4453,4458|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|Family Medical History|4485,4490|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|4485,4490|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|4485,4490|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|Family Medical History|4485,4498|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|Family Medical History|4491,4498|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|Family Medical History|4491,4498|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|Family Medical History|4491,4498|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|Family Medical History|4491,4498|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|Family Medical History|4491,4498|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|Family Medical History|4491,4498|false|false|false|||Calcium
Finding|Physiologic Function|Family Medical History|4491,4498|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|Family Medical History|4491,4498|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|Family Medical History|4532,4537|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|4532,4537|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|4532,4537|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|Family Medical History|4532,4545|false|false|false|C3824990|lactate in blood (lab test)|BLOOD Lactate
Drug|Organic Chemical|Family Medical History|4538,4545|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Drug|Pharmacologic Substance|Family Medical History|4538,4545|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Event|Event|Family Medical History|4538,4545|false|false|false|||Lactate
Procedure|Laboratory Procedure|Family Medical History|4538,4545|false|false|false|C0202115|Lactic acid measurement|Lactate
Finding|Body Substance|Family Medical History|4551,4560|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|Family Medical History|4551,4560|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|Family Medical History|4551,4560|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|Family Medical History|4551,4560|false|false|false|C0030685|Patient Discharge|DISCHARGE
Disorder|Disease or Syndrome|Family Medical History|4574,4579|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|4574,4579|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|4574,4579|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|Family Medical History|4580,4583|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|Family Medical History|4591,4594|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|Family Medical History|4591,4594|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|Family Medical History|4591,4594|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|Family Medical History|4601,4604|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Family Medical History|4601,4604|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|Family Medical History|4601,4604|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Family Medical History|4601,4604|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|Family Medical History|4610,4613|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|Family Medical History|4610,4613|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|Family Medical History|4621,4624|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|Family Medical History|4621,4624|false|false|false|||MCV
Lab|Laboratory or Test Result|Family Medical History|4621,4624|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|Family Medical History|4621,4624|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|Family Medical History|4621,4624|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|Family Medical History|4629,4632|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|Family Medical History|4629,4632|false|false|false|C0600370|methacholine|MCH
Event|Event|Family Medical History|4629,4632|false|false|false|||MCH
Finding|Gene or Genome|Family Medical History|4629,4632|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|Family Medical History|4629,4632|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|Family Medical History|4629,4632|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|Family Medical History|4639,4643|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|Family Medical History|4672,4675|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|Family Medical History|4692,4697|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|4692,4697|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|4692,4697|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|Family Medical History|4692,4705|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|Family Medical History|4692,4705|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|Family Medical History|4692,4705|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|Family Medical History|4698,4705|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|Family Medical History|4698,4705|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|Family Medical History|4698,4705|false|false|false|C0017725|glucose|Glucose
Event|Event|Family Medical History|4698,4705|false|false|false|||Glucose
Lab|Laboratory or Test Result|Family Medical History|4698,4705|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|Family Medical History|4698,4705|false|false|false|C0337438|Glucose measurement|Glucose
Event|Event|Family Medical History|4771,4774|true|false|false|||CXR
Procedure|Diagnostic Procedure|Family Medical History|4771,4774|true|false|false|C0039985|Plain chest X-ray|CXR
Finding|Intellectual Product|Impression|4800,4805|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Location or Region|Impression|4806,4821|true|false|false|C0553534|Cardiopulmonary|cardiopulmonary
Disorder|Disease or Syndrome|Impression|4806,4821|true|false|false|C4072686|Cardiovascular disease+Pulmonary disease|cardiopulmonary
Anatomy|Body Part, Organ, or Organ Component|Impression|4822,4829|true|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|Impression|4822,4829|true|false|false|C1951340|Process Pharmacologic Substance|process
Event|Event|Impression|4822,4829|true|false|false|||process
Finding|Functional Concept|Impression|4822,4829|true|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|Impression|4822,4829|true|false|false|C1522240|Process|process
Finding|Idea or Concept|Hospital Course|4862,4866|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|Hospital Course|4862,4866|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|Hospital Course|4867,4870|false|false|false|||old
Event|Event|Hospital Course|4883,4890|false|false|false|||history
Finding|Conceptual Entity|Hospital Course|4883,4890|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|4883,4890|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|4883,4890|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|4883,4893|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|Hospital Course|4894,4898|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|4894,4898|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|4894,4898|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|4894,4898|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Idea or Concept|Hospital Course|4903,4907|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|4903,4907|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|4903,4907|false|false|false|C1553498|home health encounter|home
Disorder|Disease or Syndrome|Hospital Course|4913,4916|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|Hospital Course|4913,4916|false|false|false|||HTN
Disorder|Disease or Syndrome|Hospital Course|4918,4922|false|false|false|C0004238|Atrial Fibrillation|Afib
Event|Event|Hospital Course|4918,4922|false|false|false|||Afib
Lab|Laboratory or Test Result|Hospital Course|4918,4922|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Afib
Event|Event|Hospital Course|4924,4932|false|false|false|||admitted
Event|Event|Hospital Course|4938,4945|false|false|false|||dyspnea
Finding|Finding|Hospital Course|4938,4945|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|Hospital Course|4938,4945|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Drug|Organic Chemical|Hospital Course|4950,4955|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|Hospital Course|4950,4955|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|Hospital Course|4950,4955|false|false|false|||cough
Finding|Sign or Symptom|Hospital Course|4950,4955|false|false|false|C0010200|Coughing|cough
Disorder|Disease or Syndrome|Hospital Course|4963,4967|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|4963,4967|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|4963,4967|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|4963,4967|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|Hospital Course|4963,4980|false|false|false|C0740304|COPD exacerbation|COPD exacerbation
Event|Event|Hospital Course|4968,4980|false|false|false|||exacerbation
Finding|Finding|Hospital Course|4968,4980|false|false|false|C4086268|Exacerbation|exacerbation
Event|Event|Hospital Course|4982,4992|false|false|false|||Presenting
Finding|Idea or Concept|Hospital Course|4982,4992|false|false|false|C0449450|Presentation|Presenting
Drug|Organic Chemical|Hospital Course|4998,5003|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|Hospital Course|4998,5003|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|Hospital Course|4998,5003|false|false|false|||cough
Finding|Sign or Symptom|Hospital Course|4998,5003|false|false|false|C0010200|Coughing|cough
Event|Event|Hospital Course|5005,5016|false|false|false|||significant
Finding|Idea or Concept|Hospital Course|5005,5016|false|false|false|C0750502|Significant|significant
Event|Event|Hospital Course|5018,5026|false|false|false|||wheezing
Finding|Sign or Symptom|Hospital Course|5018,5026|false|false|false|C0043144|Wheezing|wheezing
Finding|Intellectual Product|Hospital Course|5031,5035|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Drug|Inorganic Chemical|Hospital Course|5036,5039|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|Hospital Course|5036,5039|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|Hospital Course|5036,5039|false|false|false|C0001861;C3536832|Air (substance);air|air
Finding|Finding|Hospital Course|5036,5039|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|Hospital Course|5036,5039|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|Hospital Course|5036,5039|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Phenomenon|Natural Phenomenon or Process|Hospital Course|5036,5048|false|false|false|C0001868|Air Movements|air movement
Event|Event|Hospital Course|5040,5048|false|false|false|||movement
Finding|Organism Function|Hospital Course|5040,5048|false|false|false|C0026649|Movement|movement
Event|Event|Hospital Course|5059,5069|false|false|false|||consistent
Finding|Idea or Concept|Hospital Course|5059,5069|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|Hospital Course|5059,5074|false|false|false|C0332290|Consistent with|consistent with
Disorder|Disease or Syndrome|Hospital Course|5075,5079|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|5075,5079|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|5075,5079|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|5075,5079|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|Hospital Course|5081,5093|false|false|false|||exacerbation
Finding|Finding|Hospital Course|5081,5093|false|false|false|C4086268|Exacerbation|exacerbation
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Hospital Course|5098,5101|true|false|false|C0600500|Peptide Nucleic Acids|PNA
Event|Event|Hospital Course|5098,5101|true|false|false|||PNA
Event|Event|Hospital Course|5105,5108|true|false|false|||CXR
Procedure|Diagnostic Procedure|Hospital Course|5105,5108|true|false|false|C0039985|Plain chest X-ray|CXR
Finding|Functional Concept|Hospital Course|5113,5121|true|false|false|C0475224|Ischemic|ischemic
Event|Event|Hospital Course|5122,5125|true|false|false|||EKG
Finding|Intellectual Product|Hospital Course|5122,5125|true|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|Hospital Course|5122,5125|true|false|false|C1623258|Electrocardiography|EKG
Event|Event|Hospital Course|5126,5133|true|false|false|||changes
Finding|Functional Concept|Hospital Course|5126,5133|true|false|false|C0392747|Changing|changes
Event|Event|Hospital Course|5135,5143|false|false|false|||Symptoms
Finding|Functional Concept|Hospital Course|5135,5143|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|Symptoms
Finding|Sign or Symptom|Hospital Course|5135,5143|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|Symptoms
Event|Event|Hospital Course|5145,5153|false|false|false|||improved
Drug|Hormone|Hospital Course|5168,5178|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|Hospital Course|5168,5178|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|Hospital Course|5168,5178|false|false|false|C0032952|prednisone|prednisone
Event|Event|Hospital Course|5168,5178|false|false|false|||prednisone
Drug|Antibiotic|Hospital Course|5183,5194|false|false|false|C0013090|doxycycline|doxycycline
Drug|Organic Chemical|Hospital Course|5183,5194|false|false|false|C0013090|doxycycline|doxycycline
Event|Event|Hospital Course|5183,5194|false|false|false|||doxycycline
Event|Event|Hospital Course|5196,5205|false|false|false|||Evaluated
Event|Event|Hospital Course|5218,5228|false|false|false|||discharged
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5232,5237|false|false|false|C0034991|Rehabilitation therapy|rehab
Event|Event|Hospital Course|5238,5246|false|false|false|||facility
Finding|Intellectual Product|Hospital Course|5238,5246|false|false|false|C4695111|ADMIN.FACILITY|facility
Finding|Finding|Hospital Course|5251,5259|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Finding|Functional Concept|Hospital Course|5251,5259|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Procedure|Health Care Activity|Hospital Course|5251,5259|false|false|false|C0031809|Physical Examination|physical
Event|Event|Hospital Course|5260,5273|false|false|false|||strengthening
Attribute|Clinical Attribute|Hospital Course|5279,5290|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|Hospital Course|5279,5290|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|Hospital Course|5279,5290|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|Hospital Course|5279,5290|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Event|Event|Hospital Course|5291,5296|false|false|false|||rehab
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5291,5296|false|false|false|C0034991|Rehabilitation therapy|rehab
Event|Event|Hospital Course|5298,5308|false|false|false|||Discharged
Finding|Idea or Concept|Hospital Course|5312,5316|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|5312,5316|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|5312,5316|false|false|false|C1553498|home health encounter|home
Disorder|Disease or Syndrome|Hospital Course|5317,5321|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|5317,5321|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|5317,5321|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|5317,5321|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|Hospital Course|5322,5326|false|false|false|C3280240|MICROCEPHALY, EPILEPSY, AND DIABETES SYNDROME 1|meds
Event|Event|Hospital Course|5322,5326|false|false|false|||meds
Finding|Intellectual Product|Hospital Course|5322,5326|false|false|false|C4284232|Medications|meds
Drug|Organic Chemical|Hospital Course|5331,5338|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Drug|Pharmacologic Substance|Hospital Course|5331,5338|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Event|Event|Hospital Course|5331,5338|false|false|false|||steroid
Event|Event|Hospital Course|5340,5345|false|false|false|||taper
Procedure|Health Care Activity|Hospital Course|5340,5345|false|false|false|C0441640||taper
Event|Event|Hospital Course|5354,5360|false|false|false|||course
Event|Activity|Hospital Course|5382,5386|false|false|false|C0871208|Rating (action)|rate
Event|Event|Hospital Course|5382,5386|false|false|false|||rate
Finding|Idea or Concept|Hospital Course|5382,5386|false|false|false|C1549480|Amount type - Rate|rate
Finding|Finding|Hospital Course|5387,5391|false|false|false|C5575035|Well (answer to question)|well
Event|Event|Hospital Course|5392,5402|false|false|false|||controlled
Drug|Organic Chemical|Hospital Course|5407,5415|false|false|false|C1831808|apixaban|apixaban
Drug|Pharmacologic Substance|Hospital Course|5407,5415|false|false|false|C1831808|apixaban|apixaban
Event|Event|Hospital Course|5407,5415|false|false|false|||apixaban
Event|Event|Hospital Course|5419,5428|false|false|false|||continued
Event|Event|Hospital Course|5429,5438|false|false|false|||diltiazam
Event|Event|Hospital Course|5441,5450|false|false|false|||continued
Drug|Organic Chemical|Hospital Course|5451,5459|false|false|false|C1831808|apixaban|apixaban
Drug|Pharmacologic Substance|Hospital Course|5451,5459|false|false|false|C1831808|apixaban|apixaban
Event|Event|Hospital Course|5451,5459|false|false|false|||apixaban
Event|Event|Hospital Course|5462,5471|false|false|false|||continued
Drug|Organic Chemical|Hospital Course|5472,5482|false|false|false|C0002598|amiodarone|amiodarone
Drug|Pharmacologic Substance|Hospital Course|5472,5482|false|false|false|C0002598|amiodarone|amiodarone
Event|Event|Hospital Course|5472,5482|false|false|false|||amiodarone
Procedure|Laboratory Procedure|Hospital Course|5472,5482|false|false|false|C5399868|Drug assay amiodarone|amiodarone
Disorder|Disease or Syndrome|Hospital Course|5486,5492|false|false|false|C0002871|Anemia|Anemia
Event|Event|Hospital Course|5486,5492|false|false|false|||Anemia
Drug|Hazardous or Poisonous Substance|Hospital Course|5497,5500|false|false|false|C0054282|butyl phosphorotrithioate|def
Drug|Organic Chemical|Hospital Course|5497,5500|false|false|false|C0054282|butyl phosphorotrithioate|def
Finding|Gene or Genome|Hospital Course|5497,5500|false|false|false|C1823727|UTP25 gene|def
Disorder|Disease or Syndrome|Hospital Course|5501,5507|false|false|false|C0002871|Anemia|anemia
Event|Event|Hospital Course|5501,5507|false|false|false|||anemia
Event|Event|Hospital Course|5518,5527|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|5518,5527|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|Hospital Course|5529,5539|false|false|false|||discharged
Event|Event|Hospital Course|5548,5557|false|false|false|||continued
Drug|Biologically Active Substance|Hospital Course|5558,5562|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|Hospital Course|5558,5562|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|Hospital Course|5558,5562|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Procedure|Laboratory Procedure|Hospital Course|5558,5562|false|false|false|C0337439|Iron measurement|iron
Drug|Inorganic Chemical|Hospital Course|5558,5573|false|false|false|C0721124;C2825025|Iron Supplement;Iron Supplement [EPC]|iron supplement
Drug|Pharmacologic Substance|Hospital Course|5558,5573|false|false|false|C0721124;C2825025|Iron Supplement;Iron Supplement [EPC]|iron supplement
Drug|Food|Hospital Course|5563,5573|false|false|false|C0242295|Dietary Supplements|supplement
Event|Event|Hospital Course|5563,5573|false|false|false|||supplement
Finding|Functional Concept|Hospital Course|5563,5573|false|false|false|C1549514;C1947943;C2348609|Supplement;Supplement (document);Supplement - Diet Code Specification Type|supplement
Finding|Idea or Concept|Hospital Course|5563,5573|false|false|false|C1549514;C1947943;C2348609|Supplement;Supplement (document);Supplement - Diet Code Specification Type|supplement
Finding|Intellectual Product|Hospital Course|5563,5573|false|false|false|C1549514;C1947943;C2348609|Supplement;Supplement (document);Supplement - Diet Code Specification Type|supplement
Disorder|Disease or Syndrome|Hospital Course|5577,5580|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5577,5580|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|5577,5580|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Hospital Course|5577,5580|false|false|false|||CAD
Finding|Gene or Genome|Hospital Course|5577,5580|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|5577,5580|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|5577,5580|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5577,5580|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|Hospital Course|5582,5590|false|false|false|||continue
Drug|Organic Chemical|Hospital Course|5591,5598|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|Hospital Course|5591,5598|false|false|false|C0004057|aspirin|aspirin
Event|Event|Hospital Course|5591,5598|false|false|false|||aspirin
Drug|Organic Chemical|Hospital Course|5600,5612|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|Hospital Course|5600,5612|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|Hospital Course|5600,5612|false|false|false|||atorvastatin
Event|Event|Hospital Course|5615,5627|false|false|false|||Constipation
Finding|Sign or Symptom|Hospital Course|5615,5627|false|false|false|C0009806|Constipation|Constipation
Event|Event|Hospital Course|5629,5637|false|false|false|||continue
Finding|Idea or Concept|Hospital Course|5638,5642|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|5638,5642|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|5638,5642|false|false|false|C1553498|home health encounter|home
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5643,5648|false|false|false|C0021853|Intestines|bowel
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5649,5652|false|false|false|C0208940|human REG1A protein|reg
Drug|Biologically Active Substance|Hospital Course|5649,5652|false|false|false|C0208940|human REG1A protein|reg
Event|Event|Hospital Course|5649,5652|false|false|false|||reg
Finding|Gene or Genome|Hospital Course|5649,5652|false|false|false|C1419333;C1705631;C4321234|EXTL3 wt Allele;REG1A gene;REG1A wt Allele|reg
Disorder|Mental or Behavioral Dysfunction|Hospital Course|5655,5662|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|Anxiety
Event|Event|Hospital Course|5655,5662|false|false|false|||Anxiety
Finding|Sign or Symptom|Hospital Course|5655,5662|false|false|false|C0860603|Anxiety symptoms|Anxiety
Event|Event|Hospital Course|5664,5673|false|false|false|||continued
Finding|Idea or Concept|Hospital Course|5674,5678|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|5674,5678|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|5674,5678|false|false|false|C1553498|home health encounter|home
Disorder|Disease or Syndrome|Hospital Course|5679,5683|false|false|false|C3280240|MICROCEPHALY, EPILEPSY, AND DIABETES SYNDROME 1|meds
Event|Event|Hospital Course|5679,5683|false|false|false|||meds
Finding|Intellectual Product|Hospital Course|5679,5683|false|false|false|C4284232|Medications|meds
Finding|Idea or Concept|Hospital Course|5685,5697|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Event|Event|Hospital Course|5702,5712|false|false|false|||Discharged
Drug|Organic Chemical|Hospital Course|5716,5723|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Drug|Pharmacologic Substance|Hospital Course|5716,5723|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Event|Event|Hospital Course|5724,5729|false|false|false|||taper
Procedure|Health Care Activity|Hospital Course|5724,5729|false|false|false|C0441640||taper
Event|Activity|Hospital Course|5735,5746|false|false|false|C0024501|Maintenance|maintenance
Event|Event|Hospital Course|5747,5751|false|false|false|||dose
Disorder|Disease or Syndrome|Hospital Course|5782,5785|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|Hospital Course|5782,5785|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|Hospital Course|5782,5785|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5782,5785|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|Hospital Course|5782,5785|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|Hospital Course|5782,5785|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|Hospital Course|5782,5785|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|Hospital Course|5782,5785|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|Hospital Course|5782,5785|false|false|false|||PCP
Finding|Gene or Genome|Hospital Course|5782,5785|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|Hospital Course|5782,5785|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Drug|Antibiotic|Hospital Course|5801,5812|false|false|false|C0013090|doxycycline|Doxycycline
Drug|Organic Chemical|Hospital Course|5801,5812|false|false|false|C0013090|doxycycline|Doxycycline
Disorder|Mental or Behavioral Dysfunction|Hospital Course|5819,5822|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5819,5822|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|5819,5822|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|5819,5822|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|5819,5822|false|false|false|C1332410|BID gene|BID
Attribute|Clinical Attribute|Hospital Course|5832,5843|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|5832,5843|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|5832,5843|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|5832,5843|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|5832,5856|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|5847,5856|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|5847,5856|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|Hospital Course|5875,5885|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Hospital Course|5875,5885|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|Hospital Course|5875,5890|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|Hospital Course|5886,5890|false|false|false|||list
Finding|Intellectual Product|Hospital Course|5886,5890|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|Hospital Course|5894,5902|false|false|false|||accurate
Drug|Organic Chemical|Hospital Course|5907,5915|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Hospital Course|5907,5915|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Hospital Course|5907,5915|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|Hospital Course|5907,5915|false|false|false|||complete
Finding|Functional Concept|Hospital Course|5907,5915|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|5907,5915|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|Hospital Course|5920,5933|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|5920,5933|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Hospital Course|5920,5933|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|5920,5933|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|Hospital Course|5948,5951|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|5952,5956|false|false|false|C2598155||pain
Event|Event|Hospital Course|5952,5956|false|false|false|||pain
Finding|Functional Concept|Hospital Course|5952,5956|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|5952,5956|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|5961,5971|false|false|false|C0002598|amiodarone|Amiodarone
Drug|Pharmacologic Substance|Hospital Course|5961,5971|false|false|false|C0002598|amiodarone|Amiodarone
Event|Event|Hospital Course|5961,5971|false|false|false|||Amiodarone
Procedure|Laboratory Procedure|Hospital Course|5961,5971|false|false|false|C5399868|Drug assay amiodarone|Amiodarone
Drug|Organic Chemical|Hospital Course|5992,6000|false|false|false|C1831808|apixaban|Apixaban
Drug|Pharmacologic Substance|Hospital Course|5992,6000|false|false|false|C1831808|apixaban|Apixaban
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6009,6012|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6009,6012|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|6009,6012|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|6009,6012|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|6009,6012|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|6017,6026|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|Hospital Course|6017,6026|false|false|false|C0001927|albuterol|Albuterol
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6034,6037|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|Hospital Course|6034,6037|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|Hospital Course|6034,6037|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Finding|Cell Function|Hospital Course|6034,6037|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|Hospital Course|6034,6037|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6045,6048|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|Hospital Course|6045,6048|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|Hospital Course|6045,6048|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|Hospital Course|6045,6048|false|false|false|||NEB
Finding|Cell Function|Hospital Course|6045,6048|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|6045,6048|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|6056,6059|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|6060,6063|false|false|false|||SOB
Finding|Sign or Symptom|Hospital Course|6060,6063|false|false|false|C0013404|Dyspnea|SOB
Drug|Pharmacologic Substance|Hospital Course|6068,6084|false|false|false|C0003921;C2608262;C3853661|Artificial Tears;Lubricant Eye Drops;artificial tears (medication)|Artificial Tears
Finding|Body Substance|Hospital Course|6079,6084|false|false|false|C0039409;C1547924;C1611838|Tears (substance);Tears specimen|Tears
Finding|Intellectual Product|Hospital Course|6079,6084|false|false|false|C0039409;C1547924;C1611838|Tears (substance);Tears specimen|Tears
Drug|Biomedical or Dental Material|Hospital Course|6089,6093|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|Hospital Course|6089,6093|false|false|false|C1705648|Dropping|DROP
Event|Event|Hospital Course|6089,6093|false|false|false|||DROP
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6094,6103|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6099,6103|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|Hospital Course|6099,6103|false|false|false|C5848506||EYES
Finding|Gene or Genome|Hospital Course|6104,6107|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|6108,6118|false|false|false|||irritation
Finding|Intellectual Product|Hospital Course|6108,6118|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Finding|Mental Process|Hospital Course|6108,6118|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Finding|Pathologic Function|Hospital Course|6108,6118|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Phenomenon|Phenomenon or Process|Hospital Course|6108,6118|false|false|false|C0441723|Irritation|irritation
Drug|Organic Chemical|Hospital Course|6123,6130|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Hospital Course|6123,6130|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|Hospital Course|6150,6162|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|6150,6162|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|Hospital Course|6180,6189|false|false|false|C0012373|diltiazem|Diltiazem
Drug|Pharmacologic Substance|Hospital Course|6180,6189|false|false|false|C0012373|diltiazem|Diltiazem
Finding|Finding|Hospital Course|6190,6198|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|6190,6198|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Hospital Course|6199,6206|false|false|false|||Release
Finding|Functional Concept|Hospital Course|6199,6206|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|6199,6206|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6199,6206|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6217,6220|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6217,6220|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|6217,6220|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|6217,6220|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|6217,6220|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|6225,6236|false|false|false|C0165590|dorzolamide|Dorzolamide
Drug|Pharmacologic Substance|Hospital Course|6225,6236|false|false|false|C0165590|dorzolamide|Dorzolamide
Finding|Functional Concept|Hospital Course|6240,6245|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|Hospital Course|6255,6259|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|Hospital Course|6255,6259|false|false|false|C1705648|Dropping|DROP
Event|Event|Hospital Course|6255,6259|false|false|false|||DROP
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6260,6269|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6265,6269|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|Hospital Course|6265,6269|false|false|false|C5848506||EYES
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6270,6273|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6270,6273|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|6270,6273|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|6270,6273|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|6270,6273|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|6279,6290|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|6279,6290|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|Hospital Course|6279,6290|false|false|false|||Fluticasone
Drug|Organic Chemical|Hospital Course|6279,6301|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|Hospital Course|6279,6301|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|Hospital Course|6291,6301|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Event|Event|Hospital Course|6291,6301|false|false|false|||Propionate
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6302,6307|false|false|false|C0028429||NASAL
Drug|Biomedical or Dental Material|Hospital Course|6302,6307|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Organic Chemical|Hospital Course|6302,6307|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Pharmacologic Substance|Hospital Course|6302,6307|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Finding|Finding|Hospital Course|6302,6307|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Finding|Functional Concept|Hospital Course|6302,6307|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Event|Event|Hospital Course|6310,6314|false|false|false|||SPRY
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6318,6321|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6318,6321|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|6318,6321|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|6318,6321|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|6318,6321|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|6327,6338|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|6327,6338|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|6327,6349|false|false|false|C0939232|fluticasone / salmeterol|Fluticasone-Salmeterol
Drug|Organic Chemical|Hospital Course|6327,6356|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Pharmacologic Substance|Hospital Course|6327,6356|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Organic Chemical|Hospital Course|6339,6349|false|false|false|C0073992|salmeterol|Salmeterol
Drug|Pharmacologic Substance|Hospital Course|6339,6349|false|false|false|C0073992|salmeterol|Salmeterol
Event|Event|Hospital Course|6350,6356|false|false|false|||Diskus
Drug|Biomedical or Dental Material|Hospital Course|6369,6372|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Organic Chemical|Hospital Course|6369,6372|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Pharmacologic Substance|Hospital Course|6369,6372|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Event|Event|Hospital Course|6369,6372|false|false|false|||INH
Finding|Functional Concept|Hospital Course|6369,6372|false|false|false|C0205535|Inhalation Route of Administration|INH
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6376,6379|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6376,6379|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|6376,6379|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|6376,6379|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|6376,6379|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|6385,6404|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Pharmacologic Substance|Hospital Course|6385,6404|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Organic Chemical|Hospital Course|6425,6435|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|Hospital Course|6425,6435|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|Hospital Course|6425,6447|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|Hospital Course|6425,6447|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Event|Event|Hospital Course|6436,6447|false|false|false|||Mononitrate
Finding|Finding|Hospital Course|6449,6457|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|6449,6457|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Hospital Course|6458,6465|false|false|false|||Release
Finding|Functional Concept|Hospital Course|6458,6465|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|6458,6465|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6458,6465|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Hospital Course|6488,6499|false|false|false|C0090306|latanoprost|Latanoprost
Drug|Pharmacologic Substance|Hospital Course|6488,6499|false|false|false|C0090306|latanoprost|Latanoprost
Finding|Functional Concept|Hospital Course|6507,6512|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|Hospital Course|6522,6526|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|Hospital Course|6522,6526|false|false|false|C1705648|Dropping|DROP
Event|Event|Hospital Course|6527,6531|false|false|false|||LEFT
Finding|Functional Concept|Hospital Course|6527,6531|false|false|false|C1552822|Table Cell Horizontal Align - left|LEFT
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6527,6535|false|false|false|C0229090|Left eye structure|LEFT EYE
Procedure|Diagnostic Procedure|Hospital Course|6527,6535|false|false|false|C2141124|examination of left eye|LEFT EYE
Anatomy|Body Location or Region|Hospital Course|6532,6535|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|EYE
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6532,6535|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|EYE
Disorder|Disease or Syndrome|Hospital Course|6532,6535|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|EYE
Disorder|Neoplastic Process|Hospital Course|6532,6535|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|EYE
Event|Event|Hospital Course|6532,6535|false|false|false|||EYE
Finding|Body Substance|Hospital Course|6532,6535|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Finding|Finding|Hospital Course|6532,6535|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Finding|Intellectual Product|Hospital Course|6532,6535|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Event|Event|Hospital Course|6536,6539|false|false|false|||QHS
Drug|Organic Chemical|Hospital Course|6545,6554|false|false|false|C0024002|lorazepam|Lorazepam
Drug|Pharmacologic Substance|Hospital Course|6545,6554|false|false|false|C0024002|lorazepam|Lorazepam
Event|Event|Hospital Course|6565,6568|false|false|false|||QHS
Finding|Gene or Genome|Hospital Course|6569,6572|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Pharmacologic Substance|Hospital Course|6573,6581|false|false|false|C1950154|Insomnia homeopathic medication|insomnia
Event|Event|Hospital Course|6573,6581|false|false|false|||insomnia
Finding|Sign or Symptom|Hospital Course|6573,6581|false|false|false|C0917801|Sleeplessness|insomnia
Drug|Organic Chemical|Hospital Course|6587,6600|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|Hospital Course|6587,6600|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|Hospital Course|6587,6600|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Event|Event|Hospital Course|6587,6600|false|false|false|||Multivitamins
Drug|Inorganic Chemical|Hospital Course|6603,6611|false|false|false|C0026162|Minerals|minerals
Event|Event|Hospital Course|6603,6611|false|false|false|||minerals
Drug|Biomedical or Dental Material|Hospital Course|6614,6617|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|Hospital Course|6614,6617|false|false|false|||TAB
Drug|Organic Chemical|Hospital Course|6632,6642|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Pharmacologic Substance|Hospital Course|6632,6642|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Organic Chemical|Hospital Course|6664,6674|false|false|false|C0213771|tiotropium|Tiotropium
Drug|Pharmacologic Substance|Hospital Course|6664,6674|false|false|false|C0213771|tiotropium|Tiotropium
Event|Event|Hospital Course|6664,6674|false|false|false|||Tiotropium
Drug|Organic Chemical|Hospital Course|6664,6682|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Pharmacologic Substance|Hospital Course|6664,6682|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Inorganic Chemical|Hospital Course|6675,6682|false|false|false|C0006222|Bromides|Bromide
Event|Event|Hospital Course|6675,6682|false|false|false|||Bromide
Procedure|Laboratory Procedure|Hospital Course|6675,6682|false|false|false|C0202341|Bromides measurement|Bromide
Disorder|Congenital Abnormality|Hospital Course|6685,6688|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|CAP
Drug|Biomedical or Dental Material|Hospital Course|6685,6688|false|false|false|C0006935|capsule (pharmacologic)|CAP
Event|Event|Hospital Course|6685,6688|false|false|false|||CAP
Finding|Gene or Genome|Hospital Course|6685,6688|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|CAP
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6685,6688|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|CAP
Drug|Organic Chemical|Hospital Course|6703,6715|false|false|false|C0039771|theophylline|Theophylline
Drug|Pharmacologic Substance|Hospital Course|6703,6715|false|false|false|C0039771|theophylline|Theophylline
Event|Event|Hospital Course|6703,6715|false|false|false|||Theophylline
Procedure|Laboratory Procedure|Hospital Course|6703,6715|false|false|false|C0039773|Assay of theophylline|Theophylline
Drug|Organic Chemical|Hospital Course|6703,6718|false|false|false|C0939729|Theophylline SR|Theophylline SR
Drug|Pharmacologic Substance|Hospital Course|6703,6718|false|false|false|C0939729|Theophylline SR|Theophylline SR
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6729,6732|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6729,6732|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|6729,6732|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|6729,6732|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|6729,6732|false|false|false|C1332410|BID gene|BID
Drug|Element, Ion, or Isotope|Hospital Course|6738,6745|false|false|false|C2346592|Ferrous|Ferrous
Drug|Inorganic Chemical|Hospital Course|6738,6753|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Pharmacologic Substance|Hospital Course|6738,6753|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Element, Ion, or Isotope|Hospital Course|6746,6753|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Inorganic Chemical|Hospital Course|6746,6753|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Pharmacologic Substance|Hospital Course|6746,6753|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Organic Chemical|Hospital Course|6775,6783|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|6775,6783|false|false|false|C1692318|docusate|Docusate
Drug|Organic Chemical|Hospital Course|6775,6790|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|Hospital Course|6775,6790|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|Hospital Course|6784,6790|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|6784,6790|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|6784,6790|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|6784,6790|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|6784,6790|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|6784,6790|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6801,6804|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6801,6804|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|6801,6804|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|6801,6804|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|6801,6804|false|false|false|C1332410|BID gene|BID
Drug|Biomedical or Dental Material|Hospital Course|6810,6822|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Drug|Organic Chemical|Hospital Course|6810,6822|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Event|Event|Hospital Course|6810,6822|false|false|false|||Polyethylene
Drug|Organic Chemical|Hospital Course|6810,6829|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Pharmacologic Substance|Hospital Course|6810,6829|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Hazardous or Poisonous Substance|Hospital Course|6823,6829|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Drug|Organic Chemical|Hospital Course|6823,6829|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Event|Event|Hospital Course|6823,6829|false|false|false|||Glycol
Drug|Organic Chemical|Hospital Course|6849,6860|false|false|false|C0027235|ipratropium|Ipratropium
Drug|Pharmacologic Substance|Hospital Course|6849,6860|false|false|false|C0027235|ipratropium|Ipratropium
Event|Event|Hospital Course|6849,6860|false|false|false|||Ipratropium
Drug|Organic Chemical|Hospital Course|6849,6868|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Pharmacologic Substance|Hospital Course|6849,6868|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Inorganic Chemical|Hospital Course|6861,6868|false|false|false|C0006222|Bromides|Bromide
Event|Event|Hospital Course|6861,6868|false|false|false|||Bromide
Procedure|Laboratory Procedure|Hospital Course|6861,6868|false|false|false|C0202341|Bromides measurement|Bromide
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6869,6872|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|Hospital Course|6869,6872|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|Hospital Course|6869,6872|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Event|Event|Hospital Course|6869,6872|false|false|false|||Neb
Finding|Cell Function|Hospital Course|6869,6872|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|Hospital Course|6869,6872|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6875,6878|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|Hospital Course|6875,6878|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|Hospital Course|6875,6878|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|Hospital Course|6875,6878|false|false|false|||NEB
Finding|Cell Function|Hospital Course|6875,6878|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|6875,6878|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Event|Event|Hospital Course|6882,6885|false|false|false|||Q6H
Finding|Gene or Genome|Hospital Course|6886,6889|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|6890,6893|false|false|false|||SOB
Finding|Sign or Symptom|Hospital Course|6890,6893|false|false|false|C0013404|Dyspnea|SOB
Drug|Hormone|Hospital Course|6899,6909|false|false|false|C0032952|prednisone|PredniSONE
Drug|Organic Chemical|Hospital Course|6899,6909|false|false|false|C0032952|prednisone|PredniSONE
Drug|Pharmacologic Substance|Hospital Course|6899,6909|false|false|false|C0032952|prednisone|PredniSONE
Event|Event|Hospital Course|6926,6931|false|false|false|||Start
Finding|Idea or Concept|Hospital Course|6950,6954|false|false|false|C1552851|next - HtmlLinkType|Next
Event|Event|Hospital Course|6955,6962|false|false|false|||Routine
Finding|Idea or Concept|Hospital Course|6955,6962|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Finding|Intellectual Product|Hospital Course|6955,6962|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Procedure|Laboratory Procedure|Hospital Course|6955,6962|false|false|false|C1979801|Routine coag|Routine
Event|Occupational Activity|Hospital Course|6963,6977|false|false|false|C0001554|Administration occupational activities|Administration
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6963,6977|false|false|false|C1533734|Administration (procedure)|Administration
Finding|Finding|Hospital Course|6978,6982|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Finding|Idea or Concept|Hospital Course|6978,6982|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Finding|Intellectual Product|Hospital Course|6978,6982|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Attribute|Clinical Attribute|Hospital Course|6992,6998|false|false|false|C1114758||dose #
Event|Event|Hospital Course|7014,7019|false|false|false|||doses
Drug|Hormone|Hospital Course|7024,7034|false|false|false|C0032952|prednisone|PredniSONE
Drug|Organic Chemical|Hospital Course|7024,7034|false|false|false|C0032952|prednisone|PredniSONE
Drug|Pharmacologic Substance|Hospital Course|7024,7034|false|false|false|C0032952|prednisone|PredniSONE
Event|Event|Hospital Course|7051,7056|false|false|false|||Start
Event|Event|Hospital Course|7084,7088|false|false|false|||dose
Attribute|Clinical Attribute|Hospital Course|7098,7104|false|false|false|C1114758||dose #
Event|Event|Hospital Course|7120,7125|false|false|false|||doses
Drug|Hormone|Hospital Course|7130,7140|false|false|false|C0032952|prednisone|PredniSONE
Drug|Organic Chemical|Hospital Course|7130,7140|false|false|false|C0032952|prednisone|PredniSONE
Drug|Pharmacologic Substance|Hospital Course|7130,7140|false|false|false|C0032952|prednisone|PredniSONE
Event|Event|Hospital Course|7157,7162|false|false|false|||Start
Event|Event|Hospital Course|7188,7197|false|false|false|||completes
Event|Activity|Hospital Course|7211,7222|false|false|false|C0024501|Maintenance|maintenance
Event|Event|Hospital Course|7223,7227|false|false|false|||dose
Event|Event|Hospital Course|7231,7237|false|false|false|||follow
Event|Event|Hospital Course|7255,7259|false|false|false|||dose
Event|Event|Hospital Course|7263,7272|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|7263,7272|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|7263,7272|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|7263,7272|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|7263,7272|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|7263,7284|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|7273,7284|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|7273,7284|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|7273,7284|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|7273,7284|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|7289,7302|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|7289,7302|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Hospital Course|7289,7302|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|7289,7302|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|Hospital Course|7317,7320|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|7321,7325|false|false|false|C2598155||pain
Event|Event|Hospital Course|7321,7325|false|false|false|||pain
Finding|Functional Concept|Hospital Course|7321,7325|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|7321,7325|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|7330,7340|false|false|false|C0002598|amiodarone|Amiodarone
Drug|Pharmacologic Substance|Hospital Course|7330,7340|false|false|false|C0002598|amiodarone|Amiodarone
Event|Event|Hospital Course|7330,7340|false|false|false|||Amiodarone
Procedure|Laboratory Procedure|Hospital Course|7330,7340|false|false|false|C5399868|Drug assay amiodarone|Amiodarone
Drug|Organic Chemical|Hospital Course|7361,7369|false|false|false|C1831808|apixaban|Apixaban
Drug|Pharmacologic Substance|Hospital Course|7361,7369|false|false|false|C1831808|apixaban|Apixaban
Disorder|Mental or Behavioral Dysfunction|Hospital Course|7378,7381|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7378,7381|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|7378,7381|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|7378,7381|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|7378,7381|false|false|false|C1332410|BID gene|BID
Drug|Pharmacologic Substance|Hospital Course|7386,7402|false|false|false|C0003921;C2608262;C3853661|Artificial Tears;Lubricant Eye Drops;artificial tears (medication)|Artificial Tears
Finding|Body Substance|Hospital Course|7397,7402|false|false|false|C0039409;C1547924;C1611838|Tears (substance);Tears specimen|Tears
Finding|Intellectual Product|Hospital Course|7397,7402|false|false|false|C0039409;C1547924;C1611838|Tears (substance);Tears specimen|Tears
Drug|Biomedical or Dental Material|Hospital Course|7407,7411|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|Hospital Course|7407,7411|false|false|false|C1705648|Dropping|DROP
Event|Event|Hospital Course|7407,7411|false|false|false|||DROP
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7412,7421|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7417,7421|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|Hospital Course|7417,7421|false|false|false|C5848506||EYES
Finding|Gene or Genome|Hospital Course|7422,7425|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|7426,7436|false|false|false|||irritation
Finding|Intellectual Product|Hospital Course|7426,7436|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Finding|Mental Process|Hospital Course|7426,7436|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Finding|Pathologic Function|Hospital Course|7426,7436|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Phenomenon|Phenomenon or Process|Hospital Course|7426,7436|false|false|false|C0441723|Irritation|irritation
Drug|Organic Chemical|Hospital Course|7441,7448|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Hospital Course|7441,7448|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|Hospital Course|7468,7480|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|7468,7480|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|Hospital Course|7498,7507|false|false|false|C0012373|diltiazem|Diltiazem
Drug|Pharmacologic Substance|Hospital Course|7498,7507|false|false|false|C0012373|diltiazem|Diltiazem
Finding|Finding|Hospital Course|7508,7516|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|7508,7516|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Hospital Course|7517,7524|false|false|false|||Release
Finding|Functional Concept|Hospital Course|7517,7524|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|7517,7524|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7517,7524|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Disorder|Mental or Behavioral Dysfunction|Hospital Course|7535,7538|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7535,7538|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|7535,7538|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|7535,7538|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|7535,7538|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|7543,7551|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|7543,7551|false|false|false|C1692318|docusate|Docusate
Event|Event|Hospital Course|7543,7551|false|false|false|||Docusate
Drug|Organic Chemical|Hospital Course|7543,7558|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|Hospital Course|7543,7558|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|Hospital Course|7552,7558|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|7552,7558|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|7552,7558|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|7552,7558|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|7552,7558|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|7552,7558|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|Hospital Course|7569,7572|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7569,7572|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|7569,7572|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|7569,7572|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|7569,7572|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|7577,7588|false|false|false|C0165590|dorzolamide|Dorzolamide
Drug|Pharmacologic Substance|Hospital Course|7577,7588|false|false|false|C0165590|dorzolamide|Dorzolamide
Finding|Functional Concept|Hospital Course|7592,7597|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|Hospital Course|7607,7611|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|Hospital Course|7607,7611|false|false|false|C1705648|Dropping|DROP
Event|Event|Hospital Course|7607,7611|false|false|false|||DROP
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7612,7621|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7617,7621|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|Hospital Course|7617,7621|false|false|false|C5848506||EYES
Disorder|Mental or Behavioral Dysfunction|Hospital Course|7622,7625|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7622,7625|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|7622,7625|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|7622,7625|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|7622,7625|false|false|false|C1332410|BID gene|BID
Drug|Element, Ion, or Isotope|Hospital Course|7631,7638|false|false|false|C2346592|Ferrous|Ferrous
Drug|Inorganic Chemical|Hospital Course|7631,7646|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Pharmacologic Substance|Hospital Course|7631,7646|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Element, Ion, or Isotope|Hospital Course|7639,7646|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Inorganic Chemical|Hospital Course|7639,7646|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Pharmacologic Substance|Hospital Course|7639,7646|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Event|Event|Hospital Course|7639,7646|false|false|false|||Sulfate
Drug|Organic Chemical|Hospital Course|7668,7679|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|7668,7679|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|Hospital Course|7668,7679|false|false|false|||Fluticasone
Drug|Organic Chemical|Hospital Course|7668,7690|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|Hospital Course|7668,7690|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|Hospital Course|7680,7690|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Event|Event|Hospital Course|7680,7690|false|false|false|||Propionate
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7691,7696|false|false|false|C0028429||NASAL
Drug|Biomedical or Dental Material|Hospital Course|7691,7696|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Organic Chemical|Hospital Course|7691,7696|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Pharmacologic Substance|Hospital Course|7691,7696|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Finding|Finding|Hospital Course|7691,7696|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Finding|Functional Concept|Hospital Course|7691,7696|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Event|Event|Hospital Course|7699,7703|false|false|false|||SPRY
Disorder|Mental or Behavioral Dysfunction|Hospital Course|7707,7710|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7707,7710|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|7707,7710|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|7707,7710|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|7707,7710|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|7716,7727|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|7716,7727|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|7716,7738|false|false|false|C0939232|fluticasone / salmeterol|Fluticasone-Salmeterol
Drug|Organic Chemical|Hospital Course|7716,7745|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Pharmacologic Substance|Hospital Course|7716,7745|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Organic Chemical|Hospital Course|7728,7738|false|false|false|C0073992|salmeterol|Salmeterol
Drug|Pharmacologic Substance|Hospital Course|7728,7738|false|false|false|C0073992|salmeterol|Salmeterol
Event|Event|Hospital Course|7739,7745|false|false|false|||Diskus
Drug|Biomedical or Dental Material|Hospital Course|7758,7761|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Organic Chemical|Hospital Course|7758,7761|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Pharmacologic Substance|Hospital Course|7758,7761|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Event|Event|Hospital Course|7758,7761|false|false|false|||INH
Finding|Functional Concept|Hospital Course|7758,7761|false|false|false|C0205535|Inhalation Route of Administration|INH
Disorder|Mental or Behavioral Dysfunction|Hospital Course|7765,7768|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7765,7768|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|7765,7768|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|7765,7768|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|7765,7768|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|7774,7793|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Pharmacologic Substance|Hospital Course|7774,7793|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Organic Chemical|Hospital Course|7814,7824|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|Hospital Course|7814,7824|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|Hospital Course|7814,7836|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|Hospital Course|7814,7836|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Event|Event|Hospital Course|7825,7836|false|false|false|||Mononitrate
Finding|Finding|Hospital Course|7838,7846|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|7838,7846|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Hospital Course|7847,7854|false|false|false|||Release
Finding|Functional Concept|Hospital Course|7847,7854|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|7847,7854|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7847,7854|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Hospital Course|7877,7888|false|false|false|C0090306|latanoprost|Latanoprost
Drug|Pharmacologic Substance|Hospital Course|7877,7888|false|false|false|C0090306|latanoprost|Latanoprost
Finding|Functional Concept|Hospital Course|7896,7901|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|Hospital Course|7911,7915|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|Hospital Course|7911,7915|false|false|false|C1705648|Dropping|DROP
Event|Event|Hospital Course|7916,7920|false|false|false|||LEFT
Finding|Functional Concept|Hospital Course|7916,7920|false|false|false|C1552822|Table Cell Horizontal Align - left|LEFT
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7916,7924|false|false|false|C0229090|Left eye structure|LEFT EYE
Procedure|Diagnostic Procedure|Hospital Course|7916,7924|false|false|false|C2141124|examination of left eye|LEFT EYE
Anatomy|Body Location or Region|Hospital Course|7921,7924|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|EYE
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7921,7924|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|EYE
Disorder|Disease or Syndrome|Hospital Course|7921,7924|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|EYE
Disorder|Neoplastic Process|Hospital Course|7921,7924|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|EYE
Event|Event|Hospital Course|7921,7924|false|false|false|||EYE
Finding|Body Substance|Hospital Course|7921,7924|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Finding|Finding|Hospital Course|7921,7924|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Finding|Intellectual Product|Hospital Course|7921,7924|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Event|Event|Hospital Course|7925,7928|false|false|false|||QHS
Drug|Organic Chemical|Hospital Course|7934,7943|false|false|false|C0024002|lorazepam|Lorazepam
Drug|Pharmacologic Substance|Hospital Course|7934,7943|false|false|false|C0024002|lorazepam|Lorazepam
Event|Event|Hospital Course|7954,7957|false|false|false|||QHS
Finding|Gene or Genome|Hospital Course|7958,7961|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Pharmacologic Substance|Hospital Course|7962,7970|false|false|false|C1950154|Insomnia homeopathic medication|insomnia
Event|Event|Hospital Course|7962,7970|false|false|false|||insomnia
Finding|Sign or Symptom|Hospital Course|7962,7970|false|false|false|C0917801|Sleeplessness|insomnia
Drug|Organic Chemical|Hospital Course|7976,7989|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|Hospital Course|7976,7989|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|Hospital Course|7976,7989|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Event|Event|Hospital Course|7976,7989|false|false|false|||Multivitamins
Drug|Inorganic Chemical|Hospital Course|7992,8000|false|false|false|C0026162|Minerals|minerals
Event|Event|Hospital Course|7992,8000|false|false|false|||minerals
Drug|Biomedical or Dental Material|Hospital Course|8003,8006|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|Hospital Course|8003,8006|false|false|false|||TAB
Drug|Biomedical or Dental Material|Hospital Course|8021,8033|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Drug|Organic Chemical|Hospital Course|8021,8033|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Event|Event|Hospital Course|8021,8033|false|false|false|||Polyethylene
Drug|Organic Chemical|Hospital Course|8021,8040|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Pharmacologic Substance|Hospital Course|8021,8040|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Hazardous or Poisonous Substance|Hospital Course|8034,8040|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Drug|Organic Chemical|Hospital Course|8034,8040|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Event|Event|Hospital Course|8034,8040|false|false|false|||Glycol
Drug|Organic Chemical|Hospital Course|8060,8070|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Pharmacologic Substance|Hospital Course|8060,8070|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Organic Chemical|Hospital Course|8092,8104|false|false|false|C0039771|theophylline|Theophylline
Drug|Pharmacologic Substance|Hospital Course|8092,8104|false|false|false|C0039771|theophylline|Theophylline
Event|Event|Hospital Course|8092,8104|false|false|false|||Theophylline
Procedure|Laboratory Procedure|Hospital Course|8092,8104|false|false|false|C0039773|Assay of theophylline|Theophylline
Drug|Organic Chemical|Hospital Course|8092,8107|false|false|false|C0939729|Theophylline SR|Theophylline SR
Drug|Pharmacologic Substance|Hospital Course|8092,8107|false|false|false|C0939729|Theophylline SR|Theophylline SR
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8118,8121|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8118,8121|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8118,8121|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|8118,8121|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|8118,8121|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|8127,8137|false|false|false|C0213771|tiotropium|Tiotropium
Drug|Pharmacologic Substance|Hospital Course|8127,8137|false|false|false|C0213771|tiotropium|Tiotropium
Event|Event|Hospital Course|8127,8137|false|false|false|||Tiotropium
Drug|Organic Chemical|Hospital Course|8127,8145|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Pharmacologic Substance|Hospital Course|8127,8145|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Inorganic Chemical|Hospital Course|8138,8145|false|false|false|C0006222|Bromides|Bromide
Event|Event|Hospital Course|8138,8145|false|false|false|||Bromide
Procedure|Laboratory Procedure|Hospital Course|8138,8145|false|false|false|C0202341|Bromides measurement|Bromide
Disorder|Congenital Abnormality|Hospital Course|8148,8151|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|CAP
Drug|Biomedical or Dental Material|Hospital Course|8148,8151|false|false|false|C0006935|capsule (pharmacologic)|CAP
Event|Event|Hospital Course|8148,8151|false|false|false|||CAP
Finding|Gene or Genome|Hospital Course|8148,8151|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|CAP
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8148,8151|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|CAP
Drug|Organic Chemical|Hospital Course|8166,8175|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|Hospital Course|8166,8175|false|false|false|C0001927|albuterol|Albuterol
Finding|Functional Concept|Hospital Course|8176,8183|false|false|false|C4319647|Inhaler (unit of presentation)|Inhaler
Finding|Gene or Genome|Hospital Course|8200,8203|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|8204,8207|false|false|false|||SOB
Finding|Sign or Symptom|Hospital Course|8204,8207|false|false|false|C0013404|Dyspnea|SOB
Drug|Organic Chemical|Hospital Course|8213,8224|false|false|false|C0027235|ipratropium|Ipratropium
Drug|Pharmacologic Substance|Hospital Course|8213,8224|false|false|false|C0027235|ipratropium|Ipratropium
Event|Event|Hospital Course|8213,8224|false|false|false|||Ipratropium
Drug|Organic Chemical|Hospital Course|8213,8232|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Pharmacologic Substance|Hospital Course|8213,8232|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Inorganic Chemical|Hospital Course|8225,8232|false|false|false|C0006222|Bromides|Bromide
Event|Event|Hospital Course|8225,8232|false|false|false|||Bromide
Procedure|Laboratory Procedure|Hospital Course|8225,8232|false|false|false|C0202341|Bromides measurement|Bromide
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8233,8236|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|Hospital Course|8233,8236|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|Hospital Course|8233,8236|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Event|Event|Hospital Course|8233,8236|false|false|false|||Neb
Finding|Cell Function|Hospital Course|8233,8236|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|Hospital Course|8233,8236|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8239,8242|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|Hospital Course|8239,8242|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|Hospital Course|8239,8242|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|Hospital Course|8239,8242|false|false|false|||NEB
Finding|Cell Function|Hospital Course|8239,8242|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|8239,8242|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Event|Event|Hospital Course|8246,8249|false|false|false|||Q6H
Finding|Gene or Genome|Hospital Course|8250,8253|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|8254,8257|false|false|false|||SOB
Finding|Sign or Symptom|Hospital Course|8254,8257|false|false|false|C0013404|Dyspnea|SOB
Drug|Organic Chemical|Hospital Course|8263,8272|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|Hospital Course|8263,8272|false|false|false|C0001927|albuterol|Albuterol
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8280,8283|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|Hospital Course|8280,8283|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|Hospital Course|8280,8283|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Finding|Cell Function|Hospital Course|8280,8283|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|Hospital Course|8280,8283|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8291,8294|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|Hospital Course|8291,8294|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|Hospital Course|8291,8294|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|Hospital Course|8291,8294|false|false|false|||NEB
Finding|Cell Function|Hospital Course|8291,8294|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|8291,8294|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|8302,8305|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|8306,8309|false|false|false|||SOB
Finding|Sign or Symptom|Hospital Course|8306,8309|false|false|false|C0013404|Dyspnea|SOB
Drug|Antibiotic|Hospital Course|8315,8326|false|false|false|C0013090|doxycycline|Doxycycline
Drug|Organic Chemical|Hospital Course|8315,8326|false|false|false|C0013090|doxycycline|Doxycycline
Drug|Antibiotic|Hospital Course|8315,8334|false|false|false|C0058731|doxycycline hyclate|Doxycycline Hyclate
Drug|Organic Chemical|Hospital Course|8315,8334|false|false|false|C0058731|doxycycline hyclate|Doxycycline Hyclate
Drug|Pharmacologic Substance|Hospital Course|8350,8358|false|false|false|C0720099|Duration brand of oxymetazoline|Duration
Event|Event|Hospital Course|8350,8358|false|false|false|||Duration
Event|Event|Hospital Course|8362,8366|false|false|false|||Days
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8371,8374|false|false|false|C0082420|Endoglin, human|end
Drug|Immunologic Factor|Hospital Course|8371,8374|false|false|false|C0082420|Endoglin, human|end
Finding|Functional Concept|Hospital Course|8371,8374|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Finding|Gene or Genome|Hospital Course|8371,8374|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Drug|Hormone|Hospital Course|8384,8394|false|false|false|C0032952|prednisone|PredniSONE
Drug|Organic Chemical|Hospital Course|8384,8394|false|false|false|C0032952|prednisone|PredniSONE
Drug|Pharmacologic Substance|Hospital Course|8384,8394|false|false|false|C0032952|prednisone|PredniSONE
Event|Event|Hospital Course|8411,8415|false|false|false|||Take
Procedure|Health Care Activity|Hospital Course|8422,8429|false|false|false|C0441640||Tapered
Event|Event|Hospital Course|8437,8441|false|false|false|||DOWN
Event|Event|Hospital Course|8446,8455|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|8446,8455|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|8446,8455|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|8446,8455|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|8446,8455|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|8446,8467|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|8446,8467|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|8456,8467|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|8456,8467|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|8456,8467|false|false|false|C0184758|Patient disposition|Disposition
Finding|Finding|Hospital Course|8469,8477|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|8469,8477|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Procedure|Health Care Activity|Hospital Course|8469,8482|false|false|false|C0023977|long-term care|Extended Care
Event|Activity|Hospital Course|8478,8482|false|false|false|C1947933|care activity|Care
Event|Event|Hospital Course|8478,8482|false|false|false|||Care
Finding|Finding|Hospital Course|8478,8482|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Hospital Course|8478,8482|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Event|Event|Hospital Course|8485,8493|false|false|false|||Facility
Finding|Intellectual Product|Hospital Course|8485,8493|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|Hospital Course|8501,8510|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|8501,8510|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|8501,8510|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|8501,8510|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|8501,8510|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|8501,8520|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|8511,8520|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|8511,8520|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|8511,8520|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|8511,8520|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|8511,8520|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Disease or Syndrome|Hospital Course|8531,8535|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|8531,8535|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|8531,8535|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|8531,8535|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|Hospital Course|8531,8548|false|false|false|C0740304|COPD exacerbation|COPD exacerbation
Event|Event|Hospital Course|8536,8548|false|false|false|||exacerbation
Finding|Finding|Hospital Course|8536,8548|false|false|false|C4086268|Exacerbation|exacerbation
Disorder|Neoplastic Process|Hospital Course|8550,8559|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Event|Event|Hospital Course|8550,8559|false|false|false|||Secondary
Finding|Functional Concept|Hospital Course|8550,8559|false|false|false|C1522484|metastatic qualifier|Secondary
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8562,8570|false|false|false|C0018787|Heart|CORONARY
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8562,8577|false|false|false|C0205042|Coronary artery|CORONARY ARTERY
Disorder|Disease or Syndrome|Hospital Course|8562,8585|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|CORONARY ARTERY DISEASE
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8571,8577|false|false|false|C0003842;C0226004|Arterial system;Arteries|ARTERY
Anatomy|Body System|Hospital Course|8571,8577|false|false|false|C0003842;C0226004|Arterial system;Arteries|ARTERY
Disorder|Disease or Syndrome|Hospital Course|8571,8585|false|false|false|C0852949|Arteriopathic disease|ARTERY DISEASE
Disorder|Disease or Syndrome|Hospital Course|8578,8585|false|false|false|C0012634|Disease|DISEASE
Event|Event|Hospital Course|8578,8585|false|false|false|||DISEASE
Disorder|Disease or Syndrome|Hospital Course|8589,8603|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|HYPERLIPIDEMIA
Event|Event|Hospital Course|8589,8603|false|false|false|||HYPERLIPIDEMIA
Finding|Finding|Hospital Course|8589,8603|false|false|false|C0428465|Serum lipids high (finding)|HYPERLIPIDEMIA
Disorder|Disease or Syndrome|Hospital Course|8607,8619|false|false|false|C0020538|Hypertensive disease|HYPERTENSION
Event|Event|Hospital Course|8607,8619|false|false|false|||HYPERTENSION
Disorder|Disease or Syndrome|Hospital Course|8623,8637|false|false|false|C0029408|Degenerative polyarthritis|OSTEOARTHRITIS
Event|Event|Hospital Course|8623,8637|false|false|false|||OSTEOARTHRITIS
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8641,8647|false|false|false|C0018792|Heart Atrium|ATRIAL
Attribute|Clinical Attribute|Hospital Course|8641,8660|false|false|false|C2926591||ATRIAL FIBRILLATION
Disorder|Disease or Syndrome|Hospital Course|8641,8660|false|false|false|C0004238|Atrial Fibrillation|ATRIAL FIBRILLATION
Lab|Laboratory or Test Result|Hospital Course|8641,8660|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|ATRIAL FIBRILLATION
Disorder|Disease or Syndrome|Hospital Course|8648,8660|false|false|false|C0232197|Fibrillation|FIBRILLATION
Event|Event|Hospital Course|8648,8660|false|false|false|||FIBRILLATION
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8664,8671|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|ANXIETY
Event|Event|Hospital Course|8664,8671|false|false|false|||ANXIETY
Finding|Sign or Symptom|Hospital Course|8664,8671|false|false|false|C0860603|Anxiety symptoms|ANXIETY
Finding|Intellectual Product|Hospital Course|8675,8691|false|false|false|C1314977|Gastrointestinal attachment|GASTROINTESTINAL
Finding|Pathologic Function|Hospital Course|8675,8700|false|false|false|C0017181|Gastrointestinal Hemorrhage|GASTROINTESTINAL BLEEDING
Finding|Pathologic Function|Hospital Course|8692,8700|false|false|false|C0019080|Hemorrhage|BLEEDING
Disorder|Disease or Syndrome|Hospital Course|8704,8718|false|false|false|C0029408|Degenerative polyarthritis|OSTEOARTHRITIS
Event|Event|Hospital Course|8704,8718|false|false|false|||OSTEOARTHRITIS
Finding|Mental Process|Discharge Condition|8745,8751|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|8745,8758|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|8745,8758|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|8752,8758|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|8752,8758|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|8760,8765|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|8760,8765|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|8770,8778|false|false|false|||coherent
Finding|Finding|Discharge Condition|8770,8778|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|8780,8785|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|8780,8802|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|8780,8802|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|8789,8802|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|8789,8802|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|8789,8802|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|8804,8809|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|8804,8809|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|8804,8809|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|8804,8809|false|false|false|||Alert
Finding|Finding|Discharge Condition|8804,8809|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|8804,8809|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|8804,8809|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|8814,8825|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|8814,8825|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|8827,8835|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|8827,8835|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|8827,8835|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|8836,8842|false|false|false|C5889824||Status
Event|Event|Discharge Condition|8836,8842|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|8836,8842|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|Discharge Condition|8844,8854|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|8844,8854|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|8844,8854|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|8844,8854|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|8857,8865|false|false|false|||requires
Event|Event|Discharge Condition|8866,8876|false|false|false|||assistance
Finding|Social Behavior|Discharge Condition|8866,8876|false|false|false|C0018896|Helping Behavior|assistance
Drug|Amino Acid, Peptide, or Protein|Discharge Condition|8880,8883|false|false|false|C1454018|AICDA protein, human|aid
Drug|Enzyme|Discharge Condition|8880,8883|false|false|false|C1454018|AICDA protein, human|aid
Event|Event|Discharge Condition|8880,8883|false|false|false|||aid
Finding|Gene or Genome|Discharge Condition|8880,8883|false|false|false|C1421876;C3540469|AICDA gene;AICDA wt Allele|aid
Procedure|Therapeutic or Preventive Procedure|Discharge Condition|8880,8883|false|false|false|C0021588;C0280108|AID - Artificial insemination by donor;dacarbazine/doxorubicin/ifosfamide protocol|aid
Event|Event|Discharge Condition|8885,8891|false|false|false|||walker
Finding|Gene or Genome|Discharge Instructions|8930,8934|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|Discharge Instructions|8954,8962|false|false|false|||admitted
Event|Event|Discharge Instructions|8968,8980|false|false|false|||exacerbation
Finding|Finding|Discharge Instructions|8968,8980|false|false|false|C4086268|Exacerbation|exacerbation
Disorder|Disease or Syndrome|Discharge Instructions|8989,8993|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Discharge Instructions|8989,8993|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Discharge Instructions|8989,8993|false|false|false|||COPD
Finding|Gene or Genome|Discharge Instructions|8989,8993|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|Discharge Instructions|8998,9002|false|false|false|||gave
Event|Event|Discharge Instructions|9013,9023|false|false|false|||treatments
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|9013,9023|false|false|false|C0087111|Therapeutic procedure|treatments
Event|Event|Discharge Instructions|9051,9060|false|false|false|||evaluated
Finding|Finding|Discharge Instructions|9069,9077|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Finding|Functional Concept|Discharge Instructions|9069,9077|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Procedure|Health Care Activity|Discharge Instructions|9069,9077|false|false|false|C0031809|Physical Examination|physical
Finding|Intellectual Product|Discharge Instructions|9069,9085|false|false|false|C1547999|Diagnostic Service Section ID - Physical Therapy|physical therapy
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|9069,9085|false|false|false|C0949766|Physical therapy|physical therapy
Event|Event|Discharge Instructions|9078,9085|false|false|false|||therapy
Finding|Finding|Discharge Instructions|9078,9085|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|Discharge Instructions|9078,9085|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|9078,9085|false|false|false|C0087111|Therapeutic procedure|therapy
Event|Event|Discharge Instructions|9095,9106|false|false|false|||recommended
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|9109,9114|false|false|false|C0034991|Rehabilitation therapy|rehab
Event|Event|Discharge Instructions|9125,9138|false|false|false|||strengthening
Event|Event|Discharge Instructions|9143,9150|false|false|false|||improve
Attribute|Clinical Attribute|Discharge Instructions|9156,9165|false|false|false|C5885990||breathing
Event|Event|Discharge Instructions|9156,9165|false|false|false|||breathing
Finding|Finding|Discharge Instructions|9156,9165|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|Discharge Instructions|9156,9165|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|Discharge Instructions|9156,9165|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|Discharge Instructions|9156,9165|false|false|false|C1160636|respiratory system process|breathing
Attribute|Clinical Attribute|Discharge Instructions|9185,9196|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|9185,9196|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|9185,9196|false|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|9185,9196|false|false|false|C4284232|Medications|medications
Event|Event|Discharge Instructions|9200,9210|false|false|false|||prescribed
Event|Event|Discharge Instructions|9215,9221|false|false|false|||follow
Event|Event|Discharge Instructions|9235,9244|false|false|false|||providers
Finding|Functional Concept|Discharge Instructions|9235,9244|false|false|false|C1138603|Provider|providers
Finding|Functional Concept|Discharge Instructions|9262,9269|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|Discharge Instructions|9262,9269|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|Discharge Instructions|9262,9269|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|Discharge Instructions|9262,9269|false|false|false|C0199168|Medical service|medical
Procedure|Health Care Activity|Discharge Instructions|9277,9285|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|9286,9298|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|9286,9298|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|9286,9298|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

