 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|48,57|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|48,57|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|48,62|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|82,91|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|82,91|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|82,91|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|82,91|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|82,91|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|82,96|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|114,119|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|114,119|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|114,119|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|138,141|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|138,141|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|138,141|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|138,141|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|138,141|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|149,156|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|149,156|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|SIMPLE_SEGMENT|158,170|false|false|false|||NEUROSURGERY
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|158,170|false|false|false|C0524850|Neurosurgical Procedures|NEUROSURGERY
Attribute|Clinical Attribute|SIMPLE_SEGMENT|173,182|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|173,182|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|173,182|false|false|false|C0020517|Hypersensitivity|Allergies
Attribute|Clinical Attribute|SIMPLE_SEGMENT|194,203|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|194,203|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|194,203|false|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|206,228|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|214,218|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|SIMPLE_SEGMENT|214,218|false|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|SIMPLE_SEGMENT|214,228|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Event|Event|SIMPLE_SEGMENT|219,228|false|false|false|||Reactions
Event|Event|SIMPLE_SEGMENT|231,240|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|231,240|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|249,264|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|255,264|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|255,264|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|255,264|false|false|false|C5441521|Complaint (finding)|Complaint
Event|Event|SIMPLE_SEGMENT|266,275|false|false|false|||Headaches
Finding|Sign or Symptom|SIMPLE_SEGMENT|266,275|false|false|false|C0018681|Headache|Headaches
Finding|Classification|SIMPLE_SEGMENT|278,283|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|284,292|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|284,292|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|296,314|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|305,314|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|305,314|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|305,314|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|305,314|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|305,314|false|false|false|C0184661|Interventional procedure|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|322,345|false|false|false|C2066670|suboccipital craniotomy|Suboccipital craniotomy
Event|Event|SIMPLE_SEGMENT|335,345|false|false|false|||craniotomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|335,345|false|false|false|C0010280|Craniotomy|craniotomy
Event|Event|SIMPLE_SEGMENT|350,359|false|false|false|||resection
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|350,359|false|false|false|C0015252;C0728940|Excision;removal technique|resection
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|363,373|false|false|false|C0007765|Cerebellum|cerebellar
Event|Event|SIMPLE_SEGMENT|375,381|false|false|false|||lesion
Finding|Finding|SIMPLE_SEGMENT|375,381|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|SIMPLE_SEGMENT|375,381|false|false|false|C0221198;C1546698|Lesion|lesion
Event|Event|SIMPLE_SEGMENT|385,392|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|385,392|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|385,392|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|385,392|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|385,395|false|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|385,411|false|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|385,411|false|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|396,403|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|396,403|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|396,411|false|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|404,411|false|false|false|C0221423|Illness (finding)|Illness
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|441,449|false|false|false|C0006104;C0228174|Brain;Cerebral hemisphere structure (body structure)|cerebral
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|441,458|false|false|false|C0917996|Cerebral Aneurysm|cerebral aneurysm
Event|Event|SIMPLE_SEGMENT|450,458|false|false|false|||aneurysm
Finding|Pathologic Function|SIMPLE_SEGMENT|450,458|false|false|false|C0002940|Aneurysm|aneurysm
Event|Event|SIMPLE_SEGMENT|460,468|false|false|false|||clipping
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|460,468|false|false|false|C0185010|Closure by clip (procedure)|clipping
Event|Event|SIMPLE_SEGMENT|480,488|false|false|false|||presents
Event|Event|SIMPLE_SEGMENT|494,497|false|false|false|||OSH
Finding|Functional Concept|SIMPLE_SEGMENT|503,507|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|508,518|false|false|false|C0007765|Cerebellum|cerebellar
Event|Event|SIMPLE_SEGMENT|520,531|false|false|false|||hypodensity
Event|Event|SIMPLE_SEGMENT|558,564|false|false|false|||lesion
Finding|Finding|SIMPLE_SEGMENT|558,564|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|SIMPLE_SEGMENT|558,564|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Body Substance|SIMPLE_SEGMENT|566,573|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|566,573|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|566,573|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|566,581|false|false|false|C0747307|Patient-Reported|Patient reports
Event|Event|SIMPLE_SEGMENT|574,581|false|false|false|||reports
Finding|Intellectual Product|SIMPLE_SEGMENT|574,581|false|false|false|C0684224|Report (document)|reports
Procedure|Health Care Activity|SIMPLE_SEGMENT|574,581|false|false|false|C0700287|Reporting|reports
Finding|Gene or Genome|SIMPLE_SEGMENT|600,603|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|SIMPLE_SEGMENT|608,615|false|false|false|||started
Event|Event|SIMPLE_SEGMENT|623,632|false|false|false|||headaches
Finding|Sign or Symptom|SIMPLE_SEGMENT|623,632|false|false|false|C0018681|Headache|headaches
Event|Event|SIMPLE_SEGMENT|644,652|false|false|false|||abnormal
Finding|Finding|SIMPLE_SEGMENT|644,652|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Finding|Idea or Concept|SIMPLE_SEGMENT|644,652|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Event|Event|SIMPLE_SEGMENT|666,675|false|false|false|||describes
Event|Event|SIMPLE_SEGMENT|680,689|false|false|false|||headaches
Finding|Sign or Symptom|SIMPLE_SEGMENT|680,689|false|false|false|C0018681|Headache|headaches
Event|Event|SIMPLE_SEGMENT|708,715|false|false|false|||resolve
Drug|Organic Chemical|SIMPLE_SEGMENT|721,728|false|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|721,728|false|false|false|C0699142|Tylenol|Tylenol
Event|Event|SIMPLE_SEGMENT|769,776|false|false|false|||reports
Event|Event|SIMPLE_SEGMENT|784,794|false|false|false|||difficulty
Finding|Finding|SIMPLE_SEGMENT|784,794|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Finding|Finding|SIMPLE_SEGMENT|784,802|false|false|false|C0311394|Difficulty walking|difficulty walking
Event|Event|SIMPLE_SEGMENT|795,802|false|false|false|||walking
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|795,802|false|false|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Finding|Finding|SIMPLE_SEGMENT|795,802|false|false|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Finding|Sign or Symptom|SIMPLE_SEGMENT|795,802|false|false|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Event|Event|SIMPLE_SEGMENT|815,822|false|false|false|||started
Finding|Gene or Genome|SIMPLE_SEGMENT|842,845|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|SIMPLE_SEGMENT|851,860|false|false|false|||describes
Event|Event|SIMPLE_SEGMENT|865,872|false|false|false|||walking
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|865,872|false|false|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Finding|Finding|SIMPLE_SEGMENT|865,872|false|false|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Finding|Sign or Symptom|SIMPLE_SEGMENT|865,872|false|false|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|877,887|false|false|false|C0344191|Cerebellar decompression injury|staggering
Finding|Sign or Symptom|SIMPLE_SEGMENT|877,887|false|false|false|C0701824|Staggering gait|staggering
Finding|Finding|SIMPLE_SEGMENT|894,901|false|false|false|C0516750|side to side|to side
Event|Event|SIMPLE_SEGMENT|908,914|false|false|false|||denies
Attribute|Clinical Attribute|SIMPLE_SEGMENT|919,925|false|false|false|C2707266||vision
Finding|Organism Function|SIMPLE_SEGMENT|919,925|false|false|false|C0042789|Vision|vision
Event|Event|SIMPLE_SEGMENT|926,933|false|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|926,933|true|false|false|C0392747|Changing|changes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|935,941|true|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|935,941|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|935,941|true|false|false|C0027497|Nausea|nausea
Event|Event|SIMPLE_SEGMENT|943,951|false|false|false|||vomiting
Finding|Sign or Symptom|SIMPLE_SEGMENT|943,951|true|false|false|C0042963|Vomiting|vomiting
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|954,963|false|false|false|C0009676|Confusion|confusion
Event|Event|SIMPLE_SEGMENT|954,963|false|false|false|||confusion
Finding|Finding|SIMPLE_SEGMENT|954,963|false|false|false|C0683369|Clouded consciousness|confusion
Finding|Idea or Concept|SIMPLE_SEGMENT|968,972|false|false|false|C1705313|Term (lexical)|word
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|968,991|false|false|false|C0454643|Word finding difficulty (disorder)|word finding difficulty
Finding|Finding|SIMPLE_SEGMENT|973,980|false|false|false|C0037088;C0243095;C2825141|Experimental Finding;Finding;Signs and Symptoms|finding
Finding|Sign or Symptom|SIMPLE_SEGMENT|973,980|false|false|false|C0037088;C0243095;C2825141|Experimental Finding;Finding;Signs and Symptoms|finding
Event|Event|SIMPLE_SEGMENT|981,991|false|false|false|||difficulty
Finding|Finding|SIMPLE_SEGMENT|981,991|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Event|Event|SIMPLE_SEGMENT|997,1000|false|false|false|||saw
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1005,1008|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1005,1008|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1005,1008|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1005,1008|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Finding|Body Substance|SIMPLE_SEGMENT|1005,1008|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Finding|SIMPLE_SEGMENT|1005,1008|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Intellectual Product|SIMPLE_SEGMENT|1005,1008|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Event|Event|SIMPLE_SEGMENT|1009,1015|false|false|false|||doctor
Finding|Intellectual Product|SIMPLE_SEGMENT|1009,1015|false|false|false|C2348314|Doctor - Title|doctor
Finding|Idea or Concept|SIMPLE_SEGMENT|1034,1041|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|routine
Finding|Intellectual Product|SIMPLE_SEGMENT|1034,1041|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|routine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1034,1041|false|false|false|C1979801|Routine coag|routine
Event|Event|SIMPLE_SEGMENT|1042,1047|false|false|false|||visit
Finding|Social Behavior|SIMPLE_SEGMENT|1042,1047|false|false|false|C0545082|Visit|visit
Event|Event|SIMPLE_SEGMENT|1053,1061|false|false|false|||referred
Event|Event|SIMPLE_SEGMENT|1081,1091|false|false|false|||evaluation
Finding|Idea or Concept|SIMPLE_SEGMENT|1081,1091|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|SIMPLE_SEGMENT|1081,1091|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Event|Event|SIMPLE_SEGMENT|1101,1109|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|1101,1109|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|1101,1109|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|SIMPLE_SEGMENT|1118,1124|false|false|false|||showed
Event|Event|SIMPLE_SEGMENT|1128,1132|false|false|false|||area
Event|Governmental or Regulatory Activity|SIMPLE_SEGMENT|1128,1132|false|false|false|C1510751|Academic Research Enhancement Awards|area
Event|Event|SIMPLE_SEGMENT|1137,1148|false|false|false|||hypodensity
Finding|Functional Concept|SIMPLE_SEGMENT|1156,1160|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1161,1171|false|false|false|C0007765|Cerebellum|cerebellum
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1161,1171|false|false|false|C0153640|Malignant neoplasm of cerebellum|cerebellum
Event|Event|SIMPLE_SEGMENT|1188,1198|false|false|false|||underlying
Finding|Finding|SIMPLE_SEGMENT|1188,1198|false|false|false|C4722602|Underlying|underlying
Event|Event|SIMPLE_SEGMENT|1200,1206|false|false|false|||lesion
Finding|Finding|SIMPLE_SEGMENT|1200,1206|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|SIMPLE_SEGMENT|1200,1206|false|false|false|C0221198;C1546698|Lesion|lesion
Event|Event|SIMPLE_SEGMENT|1229,1240|false|false|false|||transferred
Finding|Body Substance|SIMPLE_SEGMENT|1260,1267|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1260,1267|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1260,1267|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|1268,1275|false|false|false|||reports
Finding|Pathologic Function|SIMPLE_SEGMENT|1280,1288|false|false|false|C0002940|Aneurysm|aneurysm
Event|Event|SIMPLE_SEGMENT|1289,1293|false|false|false|||clip
Finding|Gene or Genome|SIMPLE_SEGMENT|1289,1293|false|false|false|C1337111;C1413237;C1561603;C1704793;C1824746;C1824747;C2827463|CD74 gene;CLIP - Codes for radiology reports;CLIP1 gene;CLIP1 wt Allele;CLIP2 gene;POMC gene;POMC wt Allele|clip
Finding|Intellectual Product|SIMPLE_SEGMENT|1289,1293|false|false|false|C1337111;C1413237;C1561603;C1704793;C1824746;C1824747;C2827463|CD74 gene;CLIP - Codes for radiology reports;CLIP1 gene;CLIP1 wt Allele;CLIP2 gene;POMC gene;POMC wt Allele|clip
Procedure|Health Care Activity|SIMPLE_SEGMENT|1289,1293|false|false|false|C5552742|Comprehensive Lifestyle Intervention Program|clip
Event|Event|SIMPLE_SEGMENT|1301,1304|false|false|false|||MRI
Finding|Gene or Genome|SIMPLE_SEGMENT|1301,1304|true|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1301,1304|true|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|SIMPLE_SEGMENT|1301,1304|true|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Event|Event|SIMPLE_SEGMENT|1306,1316|false|false|false|||compatible
Finding|Idea or Concept|SIMPLE_SEGMENT|1306,1316|false|false|false|C0332290|Consistent with|compatible
Finding|Finding|SIMPLE_SEGMENT|1321,1341|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|1326,1333|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|1326,1333|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|1326,1333|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|1326,1333|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1326,1333|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|1326,1341|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1334,1341|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1334,1341|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1334,1341|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1352,1364|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|SIMPLE_SEGMENT|1352,1364|false|false|false|||Hypertension
Finding|Pathologic Function|SIMPLE_SEGMENT|1372,1380|false|false|false|C0002940|Aneurysm|aneurysm
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1372,1389|false|false|false|C0189711|Clipping arterial aneurysm|aneurysm clipping
Event|Event|SIMPLE_SEGMENT|1381,1389|false|false|false|||clipping
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1381,1389|false|false|false|C0185010|Closure by clip (procedure)|clipping
Finding|Functional Concept|SIMPLE_SEGMENT|1414,1420|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|1414,1428|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|1421,1428|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1421,1428|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1421,1428|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1421,1428|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|1434,1440|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|1434,1440|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|1434,1440|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|1434,1440|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|1434,1448|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|1441,1448|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1441,1448|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1441,1448|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1441,1448|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Event|Event|SIMPLE_SEGMENT|1459,1466|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|1459,1466|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|1459,1466|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|1459,1466|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|1459,1469|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1470,1476|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|SIMPLE_SEGMENT|1470,1476|false|false|false|||stroke
Finding|Finding|SIMPLE_SEGMENT|1470,1476|false|false|false|C5977286|Stroke (heart beat)|stroke
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1478,1484|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|SIMPLE_SEGMENT|1478,1484|false|false|false|||cancer
Event|Event|SIMPLE_SEGMENT|1486,1494|false|false|false|||aneurysm
Finding|Pathologic Function|SIMPLE_SEGMENT|1486,1494|true|false|false|C0002940|Aneurysm|aneurysm
Event|Event|SIMPLE_SEGMENT|1500,1508|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|1500,1508|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|1500,1508|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1500,1508|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|1500,1513|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1500,1513|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|1509,1513|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|1509,1513|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1509,1513|false|false|false|C0582103|Medical Examination|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1518,1527|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|SIMPLE_SEGMENT|1588,1591|false|false|false|||Gen
Finding|Classification|SIMPLE_SEGMENT|1588,1591|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Finding|Gene or Genome|SIMPLE_SEGMENT|1588,1591|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Event|Event|SIMPLE_SEGMENT|1600,1611|false|false|false|||comfortable
Finding|Finding|SIMPLE_SEGMENT|1600,1611|false|false|false|C5546696|Feeling comfortable|comfortable
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1613,1616|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1613,1616|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1613,1616|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|1613,1616|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1613,1616|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|1613,1616|false|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|1613,1616|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1618,1623|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1625,1631|false|false|false|C0034121|Pupil|Pupils
Finding|Functional Concept|SIMPLE_SEGMENT|1653,1657|false|false|false|C0241886|Extraocular|EOMs
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1663,1667|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|SIMPLE_SEGMENT|1663,1667|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|SIMPLE_SEGMENT|1663,1667|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|SIMPLE_SEGMENT|1669,1675|false|false|false|||Supple
Finding|Functional Concept|SIMPLE_SEGMENT|1669,1675|false|false|false|C0332254|Supple|Supple
Event|Event|SIMPLE_SEGMENT|1685,1689|false|false|false|||Warm
Finding|Finding|SIMPLE_SEGMENT|1685,1689|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|1685,1689|false|false|false|C0687712|warming process|Warm
Finding|Finding|SIMPLE_SEGMENT|1694,1698|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|1699,1707|false|false|false|||perfused
Finding|Mental Process|SIMPLE_SEGMENT|1717,1723|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1717,1730|false|false|false|C0488568;C0488569||Mental status
Finding|Finding|SIMPLE_SEGMENT|1717,1730|false|false|false|C0278060|Mental state|Mental status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1724,1730|false|false|false|C5889824||status
Event|Event|SIMPLE_SEGMENT|1724,1730|false|false|false|||status
Finding|Idea or Concept|SIMPLE_SEGMENT|1724,1730|false|false|false|C1546481|What subject filter - Status|status
Event|Event|SIMPLE_SEGMENT|1732,1737|false|false|false|||Awake
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1742,1747|false|false|false|C5890168||alert
Drug|Organic Chemical|SIMPLE_SEGMENT|1742,1747|false|false|false|C0718338|Alert brand of caffeine|alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1742,1747|false|false|false|C0718338|Alert brand of caffeine|alert
Event|Event|SIMPLE_SEGMENT|1742,1747|false|false|false|||alert
Finding|Finding|SIMPLE_SEGMENT|1742,1747|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Functional Concept|SIMPLE_SEGMENT|1742,1747|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Intellectual Product|SIMPLE_SEGMENT|1742,1747|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Event|Event|SIMPLE_SEGMENT|1749,1760|false|false|false|||cooperative
Event|Event|SIMPLE_SEGMENT|1766,1770|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|1766,1770|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1766,1770|false|false|false|C0582103|Medical Examination|exam
Event|Event|SIMPLE_SEGMENT|1772,1778|false|false|false|||normal
Event|Event|SIMPLE_SEGMENT|1779,1785|false|false|false|||affect
Finding|Mental Process|SIMPLE_SEGMENT|1779,1785|false|false|false|C0001721|Affect (mental function)|affect
Procedure|Health Care Activity|SIMPLE_SEGMENT|1779,1785|false|false|false|C2237113|assessment of affect|affect
Event|Event|SIMPLE_SEGMENT|1787,1798|false|false|false|||Orientation
Finding|Mental Process|SIMPLE_SEGMENT|1787,1798|false|false|false|C0029266|Mental Orientation|Orientation
Event|Event|SIMPLE_SEGMENT|1800,1808|false|false|false|||Oriented
Finding|Finding|SIMPLE_SEGMENT|1800,1808|false|false|false|C1961028|Oriented to place|Oriented
Finding|Finding|SIMPLE_SEGMENT|1800,1818|false|false|false|C1961030|Oriented to person|Oriented to person
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1812,1818|false|false|false|C5890614||person
Event|Event|SIMPLE_SEGMENT|1812,1818|false|false|false|||person
Finding|Intellectual Product|SIMPLE_SEGMENT|1812,1818|false|false|false|C1522390|Person Info|person
Event|Activity|SIMPLE_SEGMENT|1820,1825|false|false|false|C1882509|put - instruction imperative|place
Event|Event|SIMPLE_SEGMENT|1820,1825|false|false|false|||place
Finding|Functional Concept|SIMPLE_SEGMENT|1820,1825|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|SIMPLE_SEGMENT|1820,1825|false|false|false|C1533810||place
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1837,1845|false|false|false|C2706915||Language
Event|Event|SIMPLE_SEGMENT|1837,1845|false|false|false|||Language
Finding|Intellectual Product|SIMPLE_SEGMENT|1837,1845|false|false|false|C0033348|Programming Languages|Language
Event|Event|SIMPLE_SEGMENT|1847,1853|false|false|false|||Speech
Finding|Organism Function|SIMPLE_SEGMENT|1847,1853|false|false|false|C0037817|Speech|Speech
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1847,1853|false|false|false|C0846595|Speech assessment|Speech
Finding|Idea or Concept|SIMPLE_SEGMENT|1866,1870|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Event|Event|SIMPLE_SEGMENT|1871,1884|false|false|false|||comprehension
Finding|Mental Process|SIMPLE_SEGMENT|1871,1884|false|false|false|C0162340|Comprehension|comprehension
Event|Event|SIMPLE_SEGMENT|1889,1899|false|false|false|||repetition
Finding|Finding|SIMPLE_SEGMENT|1889,1899|false|false|false|C0205341;C2018025|Repeat;speech fluency repetition (physical finding)|repetition
Finding|Functional Concept|SIMPLE_SEGMENT|1889,1899|false|false|false|C0205341;C2018025|Repeat;speech fluency repetition (physical finding)|repetition
Event|Event|SIMPLE_SEGMENT|1901,1907|false|false|false|||Naming
Finding|Mental Process|SIMPLE_SEGMENT|1901,1907|false|false|false|C0233735|Naming (function)|Naming
Event|Event|SIMPLE_SEGMENT|1908,1914|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|1908,1914|false|false|false|C1554187|Gender Status - Intact|intact
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1919,1929|true|false|false|C0013362|Dysarthria|dysarthria
Event|Event|SIMPLE_SEGMENT|1919,1929|false|false|false|||dysarthria
Event|Event|SIMPLE_SEGMENT|1944,1950|false|false|false|||errors
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1953,1960|false|false|false|C0037303|Bone structure of cranium|Cranial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1953,1967|false|false|false|C0010268|Cranial Nerves|Cranial Nerves
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1953,1967|false|false|false|C0004992;C0496937|Benign neoplasm of cranial nerves;Neoplasm of uncertain or unknown behavior of cranial nerves|Cranial Nerves
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1961,1967|false|false|false|C0027740|Nerve|Nerves
Event|Event|SIMPLE_SEGMENT|1976,1982|false|false|false|||tested
Finding|Functional Concept|SIMPLE_SEGMENT|1987,1991|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1987,1997|false|false|false|C0229187|Structure of pupil of left eye|Left pupil
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1992,1997|false|false|false|C0034121;C1305618|Pupil|pupil
Finding|Functional Concept|SIMPLE_SEGMENT|2005,2010|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Event|Event|SIMPLE_SEGMENT|2031,2039|false|false|false|||reactive
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2031,2039|false|false|false|C4722408|Reactive Therapy|reactive
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2043,2048|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2043,2048|false|false|false|C1570446|TNFSF14 protein, human|light
Event|Event|SIMPLE_SEGMENT|2043,2048|false|false|false|||light
Finding|Finding|SIMPLE_SEGMENT|2043,2048|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|SIMPLE_SEGMENT|2043,2048|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|SIMPLE_SEGMENT|2043,2048|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2043,2048|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2043,2048|false|false|false|C0031765|Phototherapy|light
Finding|Functional Concept|SIMPLE_SEGMENT|2064,2075|false|false|false|C0241886|Extraocular|Extraocular
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2064,2085|false|false|false|C2228439|examination of extraocular movements|Extraocular movements
Event|Event|SIMPLE_SEGMENT|2076,2085|false|false|false|||movements
Finding|Organism Function|SIMPLE_SEGMENT|2076,2085|false|false|false|C0026649|Movement|movements
Event|Event|SIMPLE_SEGMENT|2086,2092|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|2086,2092|false|false|false|C1554187|Gender Status - Intact|intact
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2113,2122|false|false|false|C0028738|Nystagmus|nystagmus
Event|Event|SIMPLE_SEGMENT|2113,2122|false|false|false|||nystagmus
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2127,2130|false|false|false|C2338708;C3496273;C3496274|Lamina VII of gray matter of spinal cord;layer VII (Cajal);lobule VII|VII
Finding|Intellectual Product|SIMPLE_SEGMENT|2127,2130|false|false|false|C0445385|Roman numeral VII|VII
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2132,2138|false|false|false|C0015450|Face|Facial
Event|Event|SIMPLE_SEGMENT|2139,2147|false|false|false|||strength
Finding|Idea or Concept|SIMPLE_SEGMENT|2139,2147|false|false|false|C0808080|Strength (attribute)|strength
Event|Event|SIMPLE_SEGMENT|2152,2161|false|false|false|||sensation
Finding|Finding|SIMPLE_SEGMENT|2152,2161|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|2152,2161|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|SIMPLE_SEGMENT|2152,2161|false|false|false|C2229507|sensory exam|sensation
Event|Event|SIMPLE_SEGMENT|2162,2168|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|2162,2168|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|SIMPLE_SEGMENT|2173,2182|false|false|false|||symmetric
Finding|Conceptual Entity|SIMPLE_SEGMENT|2173,2182|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|SIMPLE_SEGMENT|2173,2182|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2188,2207|false|false|false|C0224153|Structure of sternocleidomastoid muscle|Sternocleidomastoid
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2212,2221|false|false|false|C0224361|Structure of trapezius muscle|trapezius
Event|Event|SIMPLE_SEGMENT|2222,2228|false|false|false|||normal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2247,2253|false|false|false|C0040408|Tongue|Tongue
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2247,2253|false|false|false|C0153933|Benign neoplasm of tongue|Tongue
Procedure|Health Care Activity|SIMPLE_SEGMENT|2247,2253|false|false|false|C0872394|Procedure on tongue|Tongue
Finding|Finding|SIMPLE_SEGMENT|2247,2261|false|false|false|C3693372|tongue midline|Tongue midline
Anatomy|Cell Component|SIMPLE_SEGMENT|2254,2261|false|false|false|C1660780|midline cell component|midline
Event|Event|SIMPLE_SEGMENT|2270,2284|false|false|false|||fasciculations
Finding|Sign or Symptom|SIMPLE_SEGMENT|2270,2284|true|false|false|C0015644|Muscular fasciculation|fasciculations
Event|Event|SIMPLE_SEGMENT|2287,2292|false|false|false|||Motor
Finding|Functional Concept|SIMPLE_SEGMENT|2287,2292|false|false|false|C1513492|motor movement|Motor
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2301,2305|false|false|false|C0012173;C1337615|Bulk (conceptual);Dietary Fiber|bulk
Drug|Food|SIMPLE_SEGMENT|2301,2305|false|false|false|C0012173;C1337615|Bulk (conceptual);Dietary Fiber|bulk
Event|Event|SIMPLE_SEGMENT|2301,2305|false|false|false|||bulk
Event|Event|SIMPLE_SEGMENT|2310,2314|false|false|false|||tone
Finding|Finding|SIMPLE_SEGMENT|2331,2339|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Finding|Idea or Concept|SIMPLE_SEGMENT|2331,2339|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2331,2349|true|false|false|C0013384|Dyskinetic syndrome|abnormal movements
Finding|Finding|SIMPLE_SEGMENT|2331,2349|true|false|false|C0558189|Abnormal movement|abnormal movements
Event|Event|SIMPLE_SEGMENT|2340,2349|false|false|false|||movements
Finding|Organism Function|SIMPLE_SEGMENT|2340,2349|true|false|false|C0026649|Movement|movements
Event|Event|SIMPLE_SEGMENT|2351,2358|false|false|false|||tremors
Finding|Sign or Symptom|SIMPLE_SEGMENT|2351,2358|false|false|false|C0040822|Tremor|tremors
Finding|Idea or Concept|SIMPLE_SEGMENT|2360,2368|false|false|false|C0808080|Strength (attribute)|Strength
Finding|Social Behavior|SIMPLE_SEGMENT|2374,2379|false|false|false|C0032863|Power (Psychology)|power
Finding|Finding|SIMPLE_SEGMENT|2396,2402|false|false|false|C5202796|Intensity and Distress 1|Slight
Finding|Functional Concept|SIMPLE_SEGMENT|2403,2407|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Event|Event|SIMPLE_SEGMENT|2423,2432|false|false|false|||Sensation
Finding|Finding|SIMPLE_SEGMENT|2423,2432|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|2423,2432|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Procedure|Health Care Activity|SIMPLE_SEGMENT|2423,2432|false|false|false|C2229507|sensory exam|Sensation
Event|Event|SIMPLE_SEGMENT|2434,2440|false|false|false|||Intact
Finding|Finding|SIMPLE_SEGMENT|2434,2440|false|false|false|C1554187|Gender Status - Intact|Intact
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2444,2449|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2444,2449|false|false|false|C1570446|TNFSF14 protein, human|light
Event|Event|SIMPLE_SEGMENT|2444,2449|false|false|false|||light
Finding|Finding|SIMPLE_SEGMENT|2444,2449|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|SIMPLE_SEGMENT|2444,2449|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|SIMPLE_SEGMENT|2444,2449|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2444,2449|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2444,2449|false|false|false|C0031765|Phototherapy|light
Finding|Physiologic Function|SIMPLE_SEGMENT|2444,2455|false|false|false|C0423553|Light touch|light touch
Event|Event|SIMPLE_SEGMENT|2450,2455|false|false|false|||touch
Finding|Mental Process|SIMPLE_SEGMENT|2450,2455|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|2450,2455|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2450,2455|false|false|false|C0152054|Therapeutic Touch|touch
Event|Event|SIMPLE_SEGMENT|2457,2469|false|false|false|||Coordination
Finding|Functional Concept|SIMPLE_SEGMENT|2457,2469|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Finding|Idea or Concept|SIMPLE_SEGMENT|2457,2469|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Finding|Physiologic Function|SIMPLE_SEGMENT|2457,2469|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Event|Event|SIMPLE_SEGMENT|2471,2477|false|false|false|||normal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2481,2487|false|false|false|C0016129;C0851278;C4299059|Fingers;Fingers not including thumb;Upper extremity>Finger|finger
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2493,2499|false|false|false|C0016129;C0851278;C4299059|Fingers;Fingers not including thumb;Upper extremity>Finger|finger
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2504,2508|false|false|false|C0018870|Heel|heel
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2512,2516|false|false|false|C0230444|Shin|shin
Finding|Body Substance|SIMPLE_SEGMENT|2577,2586|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|2577,2586|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|2577,2586|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|2577,2586|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|SIMPLE_SEGMENT|2589,2593|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|2589,2593|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2589,2593|false|false|false|C0582103|Medical Examination|Exam
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2602,2606|false|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2602,2606|false|false|false|C5848506||eyes
Event|Event|SIMPLE_SEGMENT|2611,2622|false|false|false|||Spontaneous
Event|Event|SIMPLE_SEGMENT|2650,2661|false|false|false|||Orientation
Finding|Mental Process|SIMPLE_SEGMENT|2650,2661|false|false|false|C0029266|Mental Orientation|Orientation
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2666,2672|false|false|false|C5890614||Person
Finding|Intellectual Product|SIMPLE_SEGMENT|2666,2672|false|false|false|C1522390|Person Info|Person
Event|Activity|SIMPLE_SEGMENT|2676,2681|false|false|false|C1882509|put - instruction imperative|Place
Event|Event|SIMPLE_SEGMENT|2676,2681|false|false|false|||Place
Finding|Functional Concept|SIMPLE_SEGMENT|2676,2681|false|false|false|C1704765|Place - dosing instruction imperative|Place
Procedure|Health Care Activity|SIMPLE_SEGMENT|2676,2681|false|false|false|C1533810||Place
Finding|Finding|SIMPLE_SEGMENT|2685,2689|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Finding|Idea or Concept|SIMPLE_SEGMENT|2685,2689|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Finding|Intellectual Product|SIMPLE_SEGMENT|2685,2689|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Event|Event|SIMPLE_SEGMENT|2699,2707|false|false|false|||commands
Finding|Gene or Genome|SIMPLE_SEGMENT|2712,2718|false|false|false|C1424587|LITAF gene|Simple
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|2722,2729|false|false|false|C1704241|complex (molecular entity)|Complex
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2739,2745|false|false|false|C0034121|Pupil|Pupils
Finding|Functional Concept|SIMPLE_SEGMENT|2748,2753|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Finding|Functional Concept|SIMPLE_SEGMENT|2766,2770|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Event|Event|SIMPLE_SEGMENT|2779,2786|false|false|false|||chronic
Finding|Intellectual Product|SIMPLE_SEGMENT|2779,2786|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|2779,2786|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2788,2791|false|false|false|C0028863|Muscle of orbit|EOM
Finding|Functional Concept|SIMPLE_SEGMENT|2788,2791|false|false|false|C0241886|Extraocular|EOM
Event|Event|SIMPLE_SEGMENT|2817,2824|false|false|false|||chronic
Finding|Intellectual Product|SIMPLE_SEGMENT|2817,2824|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|2817,2824|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Finding|Functional Concept|SIMPLE_SEGMENT|2841,2845|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2856,2860|false|false|false|C0015450;C4266571|Face;Head>Face|Face
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2856,2860|false|false|false|C3160739|FANCONI ANEMIA, COMPLEMENTATION GROUP E|Face
Event|Event|SIMPLE_SEGMENT|2856,2860|false|false|false|||Face
Finding|Gene or Genome|SIMPLE_SEGMENT|2856,2860|false|false|false|C1414531;C1423759;C2828055|ELOVL6 gene;FANCE gene;FANCE wt Allele|Face
Finding|Conceptual Entity|SIMPLE_SEGMENT|2861,2870|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|Symmetric
Finding|Finding|SIMPLE_SEGMENT|2861,2870|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|Symmetric
Finding|Finding|SIMPLE_SEGMENT|2875,2878|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Gene or Genome|SIMPLE_SEGMENT|2875,2878|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Idea or Concept|SIMPLE_SEGMENT|2875,2878|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Intellectual Product|SIMPLE_SEGMENT|2875,2878|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Anatomy|Cell Component|SIMPLE_SEGMENT|2891,2898|false|false|false|C1660780|midline cell component|Midline
Finding|Finding|SIMPLE_SEGMENT|2903,2906|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Gene or Genome|SIMPLE_SEGMENT|2903,2906|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Idea or Concept|SIMPLE_SEGMENT|2903,2906|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Intellectual Product|SIMPLE_SEGMENT|2903,2906|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Pathologic Function|SIMPLE_SEGMENT|2914,2928|false|false|false|C1504476|Pronator drift|Pronator Drift
Event|Event|SIMPLE_SEGMENT|2923,2928|false|false|false|||Drift
Finding|Finding|SIMPLE_SEGMENT|2933,2936|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Gene or Genome|SIMPLE_SEGMENT|2933,2936|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Idea or Concept|SIMPLE_SEGMENT|2933,2936|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Intellectual Product|SIMPLE_SEGMENT|2933,2936|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Event|Event|SIMPLE_SEGMENT|2946,2952|false|false|false|||Speech
Finding|Organism Function|SIMPLE_SEGMENT|2946,2952|true|false|false|C0037817|Speech|Speech
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2946,2952|true|false|false|C0846595|Speech assessment|Speech
Finding|Finding|SIMPLE_SEGMENT|2964,2967|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Gene or Genome|SIMPLE_SEGMENT|2964,2967|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Idea or Concept|SIMPLE_SEGMENT|2964,2967|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Intellectual Product|SIMPLE_SEGMENT|2964,2967|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Mental Process|SIMPLE_SEGMENT|2975,2988|false|false|false|C0162340|Comprehension|Comprehension
Event|Event|SIMPLE_SEGMENT|2989,2995|false|false|false|||Intact
Finding|Finding|SIMPLE_SEGMENT|2989,2995|false|false|false|C1554187|Gender Status - Intact|Intact
Finding|Finding|SIMPLE_SEGMENT|3000,3003|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Gene or Genome|SIMPLE_SEGMENT|3000,3003|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Idea or Concept|SIMPLE_SEGMENT|3000,3003|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Intellectual Product|SIMPLE_SEGMENT|3000,3003|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Event|Event|SIMPLE_SEGMENT|3011,3016|false|false|false|||Motor
Finding|Functional Concept|SIMPLE_SEGMENT|3011,3016|false|false|false|C1513492|motor movement|Motor
Finding|Functional Concept|SIMPLE_SEGMENT|3047,3052|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Finding|Functional Concept|SIMPLE_SEGMENT|3088,3092|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Event|Event|SIMPLE_SEGMENT|3249,3258|false|false|false|||Sensation
Finding|Finding|SIMPLE_SEGMENT|3249,3258|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3249,3258|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Procedure|Health Care Activity|SIMPLE_SEGMENT|3249,3258|false|false|false|C2229507|sensory exam|Sensation
Event|Event|SIMPLE_SEGMENT|3259,3265|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|3259,3265|false|false|false|C1554187|Gender Status - Intact|intact
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3269,3274|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3269,3274|false|false|false|C1570446|TNFSF14 protein, human|light
Finding|Finding|SIMPLE_SEGMENT|3269,3274|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|SIMPLE_SEGMENT|3269,3274|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|SIMPLE_SEGMENT|3269,3274|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3269,3274|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3269,3274|false|false|false|C0031765|Phototherapy|light
Finding|Physiologic Function|SIMPLE_SEGMENT|3269,3280|false|false|false|C0423553|Light touch|light touch
Event|Event|SIMPLE_SEGMENT|3275,3280|false|false|false|||touch
Finding|Mental Process|SIMPLE_SEGMENT|3275,3280|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3275,3280|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3275,3280|false|false|false|C0152054|Therapeutic Touch|touch
Event|Event|SIMPLE_SEGMENT|3310,3313|false|false|false|||see
Event|Event|SIMPLE_SEGMENT|3314,3317|false|false|false|||OMR
Finding|Gene or Genome|SIMPLE_SEGMENT|3314,3317|false|false|false|C1412647|ATP5F1A gene|OMR
Event|Event|SIMPLE_SEGMENT|3332,3335|false|false|false|||lab
Finding|Gene or Genome|SIMPLE_SEGMENT|3332,3335|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|lab
Finding|Intellectual Product|SIMPLE_SEGMENT|3332,3335|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|lab
Finding|Finding|SIMPLE_SEGMENT|3340,3347|false|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3340,3347|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Event|Event|SIMPLE_SEGMENT|3348,3355|false|false|false|||results
Finding|Intellectual Product|SIMPLE_SEGMENT|3359,3364|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|3365,3373|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3365,3380|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|3365,3380|false|false|false|C0489547|Hospital course|Hospital Course
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3383,3388|false|false|false|C0006104;C4266577|Brain;Head>Brain|Brain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3383,3388|false|false|false|C0006111|Brain Diseases|Brain
Finding|Finding|SIMPLE_SEGMENT|3383,3395|false|false|false|C0221505|Lesion of brain|Brain lesion
Event|Event|SIMPLE_SEGMENT|3389,3395|false|false|false|||lesion
Finding|Finding|SIMPLE_SEGMENT|3389,3395|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|SIMPLE_SEGMENT|3389,3395|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Body Substance|SIMPLE_SEGMENT|3396,3403|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|3396,3403|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|3396,3403|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|3408,3413|false|false|false|||found
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3422,3432|false|false|false|C0007765|Cerebellum|cerebellar
Event|Event|SIMPLE_SEGMENT|3433,3444|false|false|false|||hypodensity
Event|Event|SIMPLE_SEGMENT|3460,3463|false|false|false|||OSH
Event|Event|SIMPLE_SEGMENT|3465,3467|false|false|false|||CT
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|3473,3481|false|false|false|C0009924|Contrast Media|contrast
Event|Event|SIMPLE_SEGMENT|3473,3481|false|false|false|||contrast
Event|Event|SIMPLE_SEGMENT|3486,3494|false|false|false|||obtained
Event|Event|SIMPLE_SEGMENT|3529,3539|false|false|false|||concerning
Event|Event|SIMPLE_SEGMENT|3544,3554|false|false|false|||underlying
Finding|Finding|SIMPLE_SEGMENT|3555,3559|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|SIMPLE_SEGMENT|3555,3559|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|SIMPLE_SEGMENT|3555,3559|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3555,3566|false|false|false|C0746408|mass lesion|mass lesion
Event|Event|SIMPLE_SEGMENT|3560,3566|false|false|false|||lesion
Finding|Finding|SIMPLE_SEGMENT|3560,3566|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|SIMPLE_SEGMENT|3560,3566|false|false|false|C0221198;C1546698|Lesion|lesion
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3572,3585|false|false|false|C0020255|Hydrocephalus|hydrocephalus
Event|Event|SIMPLE_SEGMENT|3572,3585|false|false|false|||hydrocephalus
Event|Event|SIMPLE_SEGMENT|3605,3611|false|false|false|||unable
Finding|Finding|SIMPLE_SEGMENT|3605,3611|false|false|false|C1299582|Unable|unable
Event|Event|SIMPLE_SEGMENT|3619,3622|false|false|false|||MRI
Finding|Gene or Genome|SIMPLE_SEGMENT|3619,3622|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3619,3622|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|SIMPLE_SEGMENT|3619,3622|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Finding|Pathologic Function|SIMPLE_SEGMENT|3666,3674|false|false|false|C0002940|Aneurysm|aneurysm
Event|Event|SIMPLE_SEGMENT|3675,3679|false|false|false|||clip
Finding|Gene or Genome|SIMPLE_SEGMENT|3675,3679|false|false|false|C1337111;C1413237;C1561603;C1704793;C1824746;C1824747;C2827463|CD74 gene;CLIP - Codes for radiology reports;CLIP1 gene;CLIP1 wt Allele;CLIP2 gene;POMC gene;POMC wt Allele|clip
Finding|Intellectual Product|SIMPLE_SEGMENT|3675,3679|false|false|false|C1337111;C1413237;C1561603;C1704793;C1824746;C1824747;C2827463|CD74 gene;CLIP - Codes for radiology reports;CLIP1 gene;CLIP1 wt Allele;CLIP2 gene;POMC gene;POMC wt Allele|clip
Procedure|Health Care Activity|SIMPLE_SEGMENT|3675,3679|false|false|false|C5552742|Comprehensive Lifestyle Intervention Program|clip
Event|Event|SIMPLE_SEGMENT|3689,3695|false|false|false|||placed
Finding|Body Substance|SIMPLE_SEGMENT|3712,3719|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|3712,3719|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|3712,3719|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|3724,3732|false|false|false|||admitted
Event|Event|SIMPLE_SEGMENT|3748,3753|false|false|false|||close
Finding|Finding|SIMPLE_SEGMENT|3748,3753|false|false|false|C0587267;C3810854|Close;Closed|close
Finding|Functional Concept|SIMPLE_SEGMENT|3748,3753|false|false|false|C0587267;C3810854|Close;Closed|close
Event|Activity|SIMPLE_SEGMENT|3755,3765|false|false|false|C1283169||monitoring
Event|Event|SIMPLE_SEGMENT|3755,3765|false|false|false|||monitoring
Procedure|Health Care Activity|SIMPLE_SEGMENT|3755,3765|false|false|false|C0150369|Preventive monitoring|monitoring
Procedure|Health Care Activity|SIMPLE_SEGMENT|3770,3778|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3770,3778|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Event|Event|SIMPLE_SEGMENT|3779,3787|false|false|false|||planning
Finding|Functional Concept|SIMPLE_SEGMENT|3779,3787|false|false|false|C0032074;C1301732|Planned|planning
Finding|Mental Process|SIMPLE_SEGMENT|3779,3787|false|false|false|C0032074;C1301732|Planned|planning
Event|Event|SIMPLE_SEGMENT|3797,3804|false|false|false|||started
Drug|Organic Chemical|SIMPLE_SEGMENT|3809,3822|false|false|false|C0011777|dexamethasone|dexamethasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3809,3822|false|false|false|C0011777|dexamethasone|dexamethasone
Finding|Finding|SIMPLE_SEGMENT|3836,3840|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|SIMPLE_SEGMENT|3836,3840|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|SIMPLE_SEGMENT|3836,3840|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Finding|SIMPLE_SEGMENT|3836,3847|false|false|false|C4086564|Mass Effect|mass effect
Event|Event|SIMPLE_SEGMENT|3841,3847|false|false|false|||effect
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3852,3857|false|false|false|C0460005|Trunk structure|torso
Event|Event|SIMPLE_SEGMENT|3862,3870|false|false|false|||obtained
Event|Event|SIMPLE_SEGMENT|3878,3884|false|false|false|||showed
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3889,3893|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3889,3893|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3889,3893|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|3889,3893|false|false|false|C0740941|Lung Problem|lung
Finding|Finding|SIMPLE_SEGMENT|3889,3901|false|false|false|C0034079||lung nodules
Event|Event|SIMPLE_SEGMENT|3894,3901|false|false|false|||nodules
Event|Event|SIMPLE_SEGMENT|3903,3906|false|false|false|||see
Event|Event|SIMPLE_SEGMENT|3922,3933|false|false|false|||information
Finding|Idea or Concept|SIMPLE_SEGMENT|3922,3933|false|false|false|C0870705;C1533716;C1561527;C1561528|Acknowledgement Detail Type - Information;Error severity - Information;Information;control act - information|information
Finding|Intellectual Product|SIMPLE_SEGMENT|3922,3933|false|false|false|C0870705;C1533716;C1561527;C1561528|Acknowledgement Detail Type - Information;Error severity - Information;Information;control act - information|information
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3946,3955|false|false|false|C0034519;C0851346|Electromagnetic Radiation;Radiation|radiation
Procedure|Research Activity|SIMPLE_SEGMENT|3946,3955|false|false|false|C1522449;C1524020;C1524021|Radiation Ionizing Radiotherapy;Radiation therapy (procedure);Radiotherapy Research|radiation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3946,3955|false|false|false|C1522449;C1524020;C1524021|Radiation Ionizing Radiotherapy;Radiation therapy (procedure);Radiotherapy Research|radiation
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3946,3964|false|false|false|C2183259|diagnostic service sources radiology labs radiation oncology|radiation oncology
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3956,3964|false|false|false|C0027651|Neoplasms|oncology
Event|Event|SIMPLE_SEGMENT|3956,3964|false|false|false|||oncology
Procedure|Health Care Activity|SIMPLE_SEGMENT|3956,3964|false|false|false|C1555459|oncology services|oncology
Event|Event|SIMPLE_SEGMENT|3970,3979|false|false|false|||consulted
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3981,3985|false|false|false|C0270724|Infantile Neuroaxonal Dystrophy|Plan
Event|Event|SIMPLE_SEGMENT|3981,3985|false|false|false|||Plan
Finding|Functional Concept|SIMPLE_SEGMENT|3981,3985|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|Plan
Finding|Intellectual Product|SIMPLE_SEGMENT|3981,3985|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|Plan
Finding|Mental Process|SIMPLE_SEGMENT|3981,3985|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|Plan
Procedure|Health Care Activity|SIMPLE_SEGMENT|4000,4008|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4000,4008|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4000,4018|false|false|false|C0015252;C0728940|Excision;removal technique|surgical resection
Event|Event|SIMPLE_SEGMENT|4009,4018|false|false|false|||resection
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4009,4018|false|false|false|C0015252;C0728940|Excision;removal technique|resection
Event|Event|SIMPLE_SEGMENT|4026,4032|false|false|false|||lesion
Finding|Finding|SIMPLE_SEGMENT|4026,4032|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|SIMPLE_SEGMENT|4026,4032|false|false|false|C0221198;C1546698|Lesion|lesion
Event|Event|SIMPLE_SEGMENT|4049,4059|false|false|false|||determined
Finding|Pathologic Function|SIMPLE_SEGMENT|4070,4078|false|false|false|C0002940|Aneurysm|aneurysm
Event|Event|SIMPLE_SEGMENT|4079,4083|false|false|false|||clip
Finding|Gene or Genome|SIMPLE_SEGMENT|4079,4083|false|false|false|C1337111;C1413237;C1561603;C1704793;C1824746;C1824747;C2827463|CD74 gene;CLIP - Codes for radiology reports;CLIP1 gene;CLIP1 wt Allele;CLIP2 gene;POMC gene;POMC wt Allele|clip
Finding|Intellectual Product|SIMPLE_SEGMENT|4079,4083|false|false|false|C1337111;C1413237;C1561603;C1704793;C1824746;C1824747;C2827463|CD74 gene;CLIP - Codes for radiology reports;CLIP1 gene;CLIP1 wt Allele;CLIP2 gene;POMC gene;POMC wt Allele|clip
Procedure|Health Care Activity|SIMPLE_SEGMENT|4079,4083|false|false|false|C5552742|Comprehensive Lifestyle Intervention Program|clip
Event|Event|SIMPLE_SEGMENT|4088,4091|false|false|false|||MRI
Finding|Gene or Genome|SIMPLE_SEGMENT|4088,4091|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4088,4091|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|SIMPLE_SEGMENT|4088,4091|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Event|Event|SIMPLE_SEGMENT|4092,4102|false|false|false|||compatible
Finding|Idea or Concept|SIMPLE_SEGMENT|4092,4102|false|false|false|C0332290|Consistent with|compatible
Event|Event|SIMPLE_SEGMENT|4115,4119|false|false|false|||able
Finding|Finding|SIMPLE_SEGMENT|4115,4119|false|false|false|C1299581|Able (qualifier value)|able
Event|Event|SIMPLE_SEGMENT|4131,4134|false|false|false|||MRI
Finding|Gene or Genome|SIMPLE_SEGMENT|4131,4134|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4131,4134|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|SIMPLE_SEGMENT|4131,4134|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4131,4140|false|false|false|C4028269|Nuclear magnetic resonance imaging brain|MRI Brain
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4135,4140|false|false|false|C0006104;C4266577|Brain;Head>Brain|Brain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4135,4140|false|false|false|C0006111|Brain Diseases|Brain
Event|Event|SIMPLE_SEGMENT|4135,4140|false|false|false|||Brain
Procedure|Health Care Activity|SIMPLE_SEGMENT|4145,4153|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4145,4153|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Event|Event|SIMPLE_SEGMENT|4154,4162|false|false|false|||planning
Finding|Functional Concept|SIMPLE_SEGMENT|4154,4162|false|false|false|C0032074;C1301732|Planned|planning
Finding|Mental Process|SIMPLE_SEGMENT|4154,4162|false|false|false|C0032074;C1301732|Planned|planning
Event|Event|SIMPLE_SEGMENT|4168,4172|false|false|false|||went
Event|Event|SIMPLE_SEGMENT|4188,4195|false|false|false|||evening
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4209,4232|false|false|false|C2066670|suboccipital craniotomy|suboccipital craniotomy
Event|Event|SIMPLE_SEGMENT|4222,4232|false|false|false|||craniotomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4222,4232|false|false|false|C0010280|Craniotomy|craniotomy
Event|Event|SIMPLE_SEGMENT|4237,4246|false|false|false|||resection
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4237,4246|false|false|false|C0015252;C0728940|Excision;removal technique|resection
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4255,4265|false|false|false|C0007765|Cerebellum|cerebellar
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4255,4272|false|false|false|C0742035||cerebellar lesion
Event|Event|SIMPLE_SEGMENT|4266,4272|false|false|false|||lesion
Finding|Finding|SIMPLE_SEGMENT|4266,4272|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|SIMPLE_SEGMENT|4266,4272|false|false|false|C0221198;C1546698|Lesion|lesion
Event|Event|SIMPLE_SEGMENT|4298,4307|false|false|false|||monitored
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4318,4321|false|false|false|C0228479|Structure of intraculminate fissure|ICU
Event|Event|SIMPLE_SEGMENT|4318,4321|false|false|false|||ICU
Finding|Intellectual Product|SIMPLE_SEGMENT|4318,4321|false|false|false|C4554035|Inventory of Callous-Unemotional Traits|ICU
Event|Event|SIMPLE_SEGMENT|4333,4341|false|false|false|||remained
Event|Event|SIMPLE_SEGMENT|4378,4384|false|false|false|||stable
Finding|Intellectual Product|SIMPLE_SEGMENT|4378,4384|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|SIMPLE_SEGMENT|4394,4405|false|false|false|||transferred
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|4435,4440|false|false|false|C3714591|Floor (anatomic)|floor
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4442,4448|false|false|false|C5889824||status
Event|Event|SIMPLE_SEGMENT|4442,4448|false|false|false|||status
Finding|Idea or Concept|SIMPLE_SEGMENT|4442,4448|false|false|false|C1546481|What subject filter - Status|status
Drug|Organic Chemical|SIMPLE_SEGMENT|4454,4467|false|false|false|C0011777|dexamethasone|Dexamethasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4454,4467|false|false|false|C0011777|dexamethasone|Dexamethasone
Event|Event|SIMPLE_SEGMENT|4454,4467|false|false|false|||Dexamethasone
Event|Event|SIMPLE_SEGMENT|4472,4479|false|false|false|||ordered
Event|Event|SIMPLE_SEGMENT|4483,4488|false|false|false|||taper
Event|Activity|SIMPLE_SEGMENT|4500,4511|false|false|false|C0024501|Maintenance|maintenance
Event|Event|SIMPLE_SEGMENT|4512,4516|false|false|false|||dose
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|4524,4527|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4524,4527|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4524,4527|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|4524,4527|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|4524,4527|false|false|false|C1332410|BID gene|BID
Finding|Intellectual Product|SIMPLE_SEGMENT|4551,4555|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|SIMPLE_SEGMENT|4562,4571|false|false|false|||pathology
Finding|Functional Concept|SIMPLE_SEGMENT|4562,4571|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Finding|Pathologic Function|SIMPLE_SEGMENT|4562,4571|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4562,4571|false|false|false|C0919386|Pathology procedure|pathology
Event|Event|SIMPLE_SEGMENT|4572,4581|false|false|false|||finalized
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4585,4610|false|false|false|C0149925|Small cell carcinoma of lung|small cell lung carcinoma
Anatomy|Cell|SIMPLE_SEGMENT|4591,4595|false|false|false|C0007634|Cells|cell
Finding|Gene or Genome|SIMPLE_SEGMENT|4591,4595|false|false|false|C1413336;C1413337|CEL gene;CELP gene|cell
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4596,4600|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4596,4600|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4596,4600|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|4596,4600|false|false|false|C0740941|Lung Problem|lung
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4596,4610|false|false|false|C0684249|Carcinoma of lung|lung carcinoma
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4601,4610|false|false|false|C0007097|Carcinoma|carcinoma
Event|Event|SIMPLE_SEGMENT|4601,4610|false|false|false|||carcinoma
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4615,4619|false|false|false|C0024109;C4037972|Chest>Lung;Lung|Lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4615,4619|false|false|false|C0024109;C4037972|Chest>Lung;Lung|Lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4615,4619|false|false|false|C0024115|Lung diseases|Lung
Finding|Finding|SIMPLE_SEGMENT|4615,4619|false|false|false|C0740941|Lung Problem|Lung
Event|Event|SIMPLE_SEGMENT|4620,4627|false|false|false|||lesions
Finding|Finding|SIMPLE_SEGMENT|4620,4627|false|false|false|C0221198|Lesion|lesions
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4631,4636|false|false|false|C0460005|Trunk structure|torso
Event|Event|SIMPLE_SEGMENT|4641,4649|false|false|false|||obtained
Event|Event|SIMPLE_SEGMENT|4656,4662|false|false|false|||showed
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4667,4671|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4667,4671|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4667,4671|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|4667,4671|false|false|false|C0740941|Lung Problem|lung
Finding|Finding|SIMPLE_SEGMENT|4667,4679|false|false|false|C0034079||lung nodules
Event|Event|SIMPLE_SEGMENT|4672,4679|false|false|false|||nodules
Finding|Functional Concept|SIMPLE_SEGMENT|4693,4697|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4722,4728|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4722,4733|false|false|false|C0003489;C4037976|Aortic arch structure;Chest>Aortic arch|aortic arch
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|4722,4733|false|false|false|C4759703|Aortic arch malformation|aortic arch
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4729,4733|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4729,4733|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4729,4733|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Finding|Finding|SIMPLE_SEGMENT|4729,4733|false|false|false|C1538146;C4722404|Age-Related Clonal Hematopoiesis;ZBTB8OS gene|arch
Finding|Gene or Genome|SIMPLE_SEGMENT|4729,4733|false|false|false|C1538146;C4722404|Age-Related Clonal Hematopoiesis;ZBTB8OS gene|arch
Finding|Functional Concept|SIMPLE_SEGMENT|4756,4761|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4756,4772|false|false|false|C1261074|Structure of right upper lobe of lung|right upper lobe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4762,4772|false|false|false|C0225756|Structure of upper lobe of lung|upper lobe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4768,4772|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|SIMPLE_SEGMENT|4768,4772|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4774,4783|false|false|false|C0024109|Lung|Pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4774,4783|false|false|false|C2707265||Pulmonary
Finding|Finding|SIMPLE_SEGMENT|4774,4783|false|false|false|C4522268|Pulmonary (intended site)|Pulmonary
Event|Event|SIMPLE_SEGMENT|4788,4797|false|false|false|||consulted
Event|Event|SIMPLE_SEGMENT|4802,4808|false|false|false|||stated
Event|Event|SIMPLE_SEGMENT|4826,4838|false|false|false|||intervention
Procedure|Health Care Activity|SIMPLE_SEGMENT|4826,4838|false|false|false|C0184661;C0886296;C1273869|Intervention regimes;Interventional procedure;Nursing interventions|intervention
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4826,4838|false|false|false|C0184661;C0886296;C1273869|Intervention regimes;Interventional procedure;Nursing interventions|intervention
Event|Event|SIMPLE_SEGMENT|4843,4852|false|false|false|||indicated
Finding|Idea or Concept|SIMPLE_SEGMENT|4859,4864|false|false|false|C1546485|Diagnosis Type - Final|final
Event|Event|SIMPLE_SEGMENT|4865,4874|false|false|false|||pathology
Finding|Functional Concept|SIMPLE_SEGMENT|4865,4874|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Finding|Pathologic Function|SIMPLE_SEGMENT|4865,4874|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4865,4874|false|false|false|C0919386|Pathology procedure|pathology
Event|Event|SIMPLE_SEGMENT|4880,4884|false|false|false|||back
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4886,4890|false|false|false|C0018966|Heme|Heme
Drug|Organic Chemical|SIMPLE_SEGMENT|4886,4890|false|false|false|C0018966|Heme|Heme
Event|Event|SIMPLE_SEGMENT|4904,4913|false|false|false|||consulted
Event|Event|SIMPLE_SEGMENT|4924,4939|false|false|false|||recommendations
Finding|Idea or Concept|SIMPLE_SEGMENT|4924,4939|false|false|false|C0034866|Recommendation|recommendations
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4957,4961|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4957,4961|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4957,4961|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|4957,4961|false|false|false|C0740941|Lung Problem|lung
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4957,4969|true|false|false|C0203683|Radioisotope scan of lung|lung imaging
Event|Event|SIMPLE_SEGMENT|4962,4969|false|false|false|||imaging
Finding|Finding|SIMPLE_SEGMENT|4962,4969|true|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4962,4969|true|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4982,4986|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4982,4986|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4982,4986|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|4982,4986|false|false|false|C0740941|Lung Problem|lung
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4982,4993|false|false|false|C0189485|Biopsy of lung|lung biopsy
Event|Event|SIMPLE_SEGMENT|4987,4993|false|false|false|||biopsy
Finding|Finding|SIMPLE_SEGMENT|4987,4993|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Finding|Intellectual Product|SIMPLE_SEGMENT|4987,4993|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4987,4993|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Procedure|Health Care Activity|SIMPLE_SEGMENT|4987,4993|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Event|Event|SIMPLE_SEGMENT|4998,5004|false|false|false|||needed
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5012,5021|false|false|false|C0024109|Lung|Pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5012,5021|false|false|false|C2707265||Pulmonary
Finding|Finding|SIMPLE_SEGMENT|5012,5021|false|false|false|C4522268|Pulmonary (intended site)|Pulmonary
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5026,5030|false|false|false|C0018966|Heme|Heme
Drug|Organic Chemical|SIMPLE_SEGMENT|5026,5030|false|false|false|C0018966|Heme|Heme
Event|Event|SIMPLE_SEGMENT|5035,5041|false|false|false|||stated
Event|Event|SIMPLE_SEGMENT|5047,5054|false|false|false|||staging
Finding|Functional Concept|SIMPLE_SEGMENT|5047,5054|false|false|false|C0332305|With staging|staging
Event|Event|SIMPLE_SEGMENT|5059,5068|false|false|false|||treatment
Finding|Conceptual Entity|SIMPLE_SEGMENT|5059,5068|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|SIMPLE_SEGMENT|5059,5068|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|SIMPLE_SEGMENT|5059,5068|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5059,5068|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Event|Event|SIMPLE_SEGMENT|5079,5089|false|false|false|||determined
Anatomy|Tissue|SIMPLE_SEGMENT|5103,5109|false|false|false|C0040300|Body tissue|tissue
Finding|Intellectual Product|SIMPLE_SEGMENT|5103,5109|false|false|false|C1547928|Tissue Specimen Code|tissue
Event|Event|SIMPLE_SEGMENT|5110,5119|false|false|false|||pathology
Finding|Functional Concept|SIMPLE_SEGMENT|5110,5119|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Finding|Pathologic Function|SIMPLE_SEGMENT|5110,5119|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5110,5119|false|false|false|C0919386|Pathology procedure|pathology
Event|Event|SIMPLE_SEGMENT|5125,5134|false|false|false|||resection
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5125,5134|false|false|false|C0015252;C0728940|Excision;removal technique|resection
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5143,5148|false|false|false|C0006104;C4266577|Brain;Head>Brain|brain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5143,5148|false|false|false|C0006111|Brain Diseases|brain
Finding|Finding|SIMPLE_SEGMENT|5143,5155|false|false|false|C0221505|Lesion of brain|brain lesion
Event|Event|SIMPLE_SEGMENT|5149,5155|false|false|false|||lesion
Finding|Finding|SIMPLE_SEGMENT|5149,5155|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|SIMPLE_SEGMENT|5149,5155|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Idea or Concept|SIMPLE_SEGMENT|5161,5166|false|false|false|C1546485|Diagnosis Type - Final|final
Event|Event|SIMPLE_SEGMENT|5167,5176|false|false|false|||pathology
Finding|Functional Concept|SIMPLE_SEGMENT|5167,5176|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Finding|Pathologic Function|SIMPLE_SEGMENT|5167,5176|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5167,5176|false|false|false|C0919386|Pathology procedure|pathology
Event|Event|SIMPLE_SEGMENT|5177,5181|false|false|false|||came
Anatomy|Cell|SIMPLE_SEGMENT|5196,5200|false|false|false|C0007634|Cells|cell
Finding|Gene or Genome|SIMPLE_SEGMENT|5196,5200|false|false|false|C1413336;C1413337|CEL gene;CELP gene|cell
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5202,5206|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5202,5206|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5202,5206|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|5202,5206|false|false|false|C0740941|Lung Problem|lung
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5202,5216|false|false|false|C0684249|Carcinoma of lung|lung carcinoma
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5207,5216|false|false|false|C0007097|Carcinoma|carcinoma
Event|Event|SIMPLE_SEGMENT|5207,5216|false|false|false|||carcinoma
Event|Event|SIMPLE_SEGMENT|5227,5233|false|false|false|||follow
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5246,5254|false|false|false|C0817096|Chest|thoracic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5246,5254|false|false|false|C5779551|Dissecting Thoracic Aortic Aneurysm|thoracic
Drug|Organic Chemical|SIMPLE_SEGMENT|5278,5285|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|Steroid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5278,5285|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|Steroid
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5278,5307|false|false|false|C0745098|Hyperglycemia steroid-induced|Steroid-induced hyperglycemia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5294,5307|false|false|false|C0020456|Hyperglycemia|hyperglycemia
Event|Event|SIMPLE_SEGMENT|5294,5307|false|false|false|||hyperglycemia
Finding|Finding|SIMPLE_SEGMENT|5294,5307|false|false|false|C2919432|Glucose in blood specimen above reference range|hyperglycemia
Event|Event|SIMPLE_SEGMENT|5323,5332|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|5323,5332|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Body Substance|SIMPLE_SEGMENT|5338,5345|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|5338,5345|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|5338,5345|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|5361,5369|false|false|false|||required
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5379,5384|false|false|false|C0222045|Integumentary scale|scale
Event|Activity|SIMPLE_SEGMENT|5379,5384|false|false|false|C1947916|Scaling|scale
Finding|Conceptual Entity|SIMPLE_SEGMENT|5379,5384|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Finding|Intellectual Product|SIMPLE_SEGMENT|5379,5384|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5385,5392|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Hormone|SIMPLE_SEGMENT|5385,5392|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5385,5392|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Event|Event|SIMPLE_SEGMENT|5385,5392|false|false|false|||Insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|5385,5392|false|false|false|C1337112|INS gene|Insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5385,5392|false|false|false|C0202098|Insulin measurement|Insulin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5406,5411|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|5406,5411|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|5406,5411|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Organic Chemical|SIMPLE_SEGMENT|5406,5418|false|false|false|C0005802|Blood Glucose|blood sugars
Drug|Organic Chemical|SIMPLE_SEGMENT|5412,5418|false|false|false|C0242209|Sugars|sugars
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5412,5418|false|false|false|C0242209|Sugars|sugars
Event|Event|SIMPLE_SEGMENT|5412,5418|false|false|false|||sugars
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5412,5418|false|false|false|C2239291|sugars (lab test)|sugars
Drug|Organic Chemical|SIMPLE_SEGMENT|5429,5442|false|false|false|C0011777|dexamethasone|Dexamethasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5429,5442|false|false|false|C0011777|dexamethasone|Dexamethasone
Event|Event|SIMPLE_SEGMENT|5429,5442|false|false|false|||Dexamethasone
Event|Event|SIMPLE_SEGMENT|5452,5461|false|false|false|||evaluated
Event|Event|SIMPLE_SEGMENT|5473,5482|false|false|false|||inpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|5473,5482|false|false|false|C1548438;C1549404|Patient Class - Inpatient;Referral category - Inpatient|inpatient
Procedure|Health Care Activity|SIMPLE_SEGMENT|5473,5482|false|false|false|C1555324|inpatient encounter|inpatient
Event|Event|SIMPLE_SEGMENT|5501,5508|false|false|false|||decided
Event|Event|SIMPLE_SEGMENT|5526,5530|false|false|false|||need
Event|Event|SIMPLE_SEGMENT|5537,5541|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|5537,5541|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|5537,5541|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|5537,5541|false|false|false|C1553498|home health encounter|home
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5545,5552|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Hormone|SIMPLE_SEGMENT|5545,5552|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5545,5552|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Event|Event|SIMPLE_SEGMENT|5545,5552|false|false|false|||Insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|5545,5552|false|false|false|C1337112|INS gene|Insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5545,5552|false|false|false|C0202098|Insulin measurement|Insulin
Event|Event|SIMPLE_SEGMENT|5560,5571|false|false|false|||recommended
Event|Event|SIMPLE_SEGMENT|5572,5583|false|false|false|||discharging
Event|Event|SIMPLE_SEGMENT|5595,5605|false|false|false|||glucometer
Event|Event|SIMPLE_SEGMENT|5625,5630|false|false|false|||check
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5635,5640|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|5635,5640|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|5635,5640|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Organic Chemical|SIMPLE_SEGMENT|5635,5647|false|false|false|C0005802|Blood Glucose|blood sugars
Drug|Organic Chemical|SIMPLE_SEGMENT|5641,5647|false|false|false|C0242209|Sugars|sugars
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5641,5647|false|false|false|C0242209|Sugars|sugars
Event|Event|SIMPLE_SEGMENT|5641,5647|false|false|false|||sugars
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5641,5647|false|false|false|C2239291|sugars (lab test)|sugars
Finding|Idea or Concept|SIMPLE_SEGMENT|5661,5665|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Finding|Intellectual Product|SIMPLE_SEGMENT|5661,5665|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5666,5671|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|5666,5671|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|5666,5671|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Organic Chemical|SIMPLE_SEGMENT|5666,5677|false|false|false|C0005802|Blood Glucose|blood sugar
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5666,5677|false|false|false|C0392201|Blood glucose measurement|blood sugar
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5672,5677|false|false|false|C0007004;C0242209;C3665462|Carbohydrates;Sugars;raw sugar|sugar
Drug|Organic Chemical|SIMPLE_SEGMENT|5672,5677|false|false|false|C0007004;C0242209;C3665462|Carbohydrates;Sugars;raw sugar|sugar
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5672,5677|false|false|false|C0007004;C0242209;C3665462|Carbohydrates;Sugars;raw sugar|sugar
Event|Event|SIMPLE_SEGMENT|5678,5682|false|false|false|||less
Event|Event|SIMPLE_SEGMENT|5702,5709|false|false|false|||advised
Event|Event|SIMPLE_SEGMENT|5713,5719|false|false|false|||record
Event|Event|SIMPLE_SEGMENT|5724,5732|false|false|false|||readings
Event|Event|SIMPLE_SEGMENT|5737,5743|false|false|false|||follow
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5757,5760|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|5757,5760|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5757,5760|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5757,5760|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|5757,5760|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|5757,5760|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|5757,5760|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5757,5760|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|5757,5760|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|5757,5760|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|5757,5760|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|SIMPLE_SEGMENT|5773,5784|false|false|false|||Bradycardia
Finding|Finding|SIMPLE_SEGMENT|5773,5784|false|false|false|C0428977;C3812171|Bradycardia;Bradycardia by ECG Finding|Bradycardia
Event|Event|SIMPLE_SEGMENT|5800,5808|false|false|false|||transfer
Finding|Functional Concept|SIMPLE_SEGMENT|5800,5808|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|SIMPLE_SEGMENT|5800,5808|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|SIMPLE_SEGMENT|5800,5808|false|false|false|C4706767|Transfer (immobility management)|transfer
Finding|Gene or Genome|SIMPLE_SEGMENT|5827,5831|false|false|false|C1420638;C1539127;C1710283|CORO7 gene;TCF21 gene;TCF21 wt Allele|POD1
Event|Event|SIMPLE_SEGMENT|5846,5850|false|false|false|||kept
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5858,5861|false|false|false|C0228479|Structure of intraculminate fissure|ICU
Finding|Intellectual Product|SIMPLE_SEGMENT|5858,5861|false|false|false|C4554035|Inventory of Callous-Unemotional Traits|ICU
Finding|Finding|SIMPLE_SEGMENT|5866,5878|false|false|false|C0231221;C0332151|Asymptomatic (finding);Asymptomatic diagnosis of|asymptomatic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5866,5890|false|false|false|C0741624|Asymptomatic bradycardia|asymptomatic bradycardia
Event|Event|SIMPLE_SEGMENT|5879,5890|false|false|false|||bradycardia
Finding|Finding|SIMPLE_SEGMENT|5879,5890|false|false|false|C0428977;C3812171|Bradycardia;Bradycardia by ECG Finding|bradycardia
Event|Event|SIMPLE_SEGMENT|5908,5916|false|false|false|||remained
Event|Event|SIMPLE_SEGMENT|5917,5929|false|false|false|||asymptomatic
Finding|Finding|SIMPLE_SEGMENT|5917,5929|false|false|false|C0231221;C0332151|Asymptomatic (finding);Asymptomatic diagnosis of|asymptomatic
Event|Event|SIMPLE_SEGMENT|5939,5948|false|false|false|||heartrate
Event|Event|SIMPLE_SEGMENT|5949,5957|false|false|false|||improved
Drug|Substance|SIMPLE_SEGMENT|5963,5969|false|false|false|C0302908|Liquid substance|fluids
Event|Event|SIMPLE_SEGMENT|5963,5969|false|false|false|||fluids
Finding|Body Substance|SIMPLE_SEGMENT|5963,5969|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5963,5969|false|false|false|C0016286|Fluid Therapy|fluids
Event|Event|SIMPLE_SEGMENT|5976,5990|false|false|false|||administration
Event|Occupational Activity|SIMPLE_SEGMENT|5976,5990|false|false|false|C0001554|Administration occupational activities|administration
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5976,5990|false|false|false|C1533734|Administration (procedure)|administration
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5998,6011|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Hormone|SIMPLE_SEGMENT|5998,6011|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Organic Chemical|SIMPLE_SEGMENT|5998,6011|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5998,6011|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Event|Event|SIMPLE_SEGMENT|5998,6011|false|false|false|||levothyroxine
Event|Event|SIMPLE_SEGMENT|6033,6039|false|false|false|||dipped
Event|Event|SIMPLE_SEGMENT|6060,6068|false|false|false|||remained
Event|Event|SIMPLE_SEGMENT|6069,6081|false|false|false|||asymptomatic
Finding|Finding|SIMPLE_SEGMENT|6069,6081|false|false|false|C0231221;C0332151|Asymptomatic (finding);Asymptomatic diagnosis of|asymptomatic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6085,6097|false|false|false|C0015469;C0376175|Bell Palsy;Facial paralysis|Bell's palsy
Event|Event|SIMPLE_SEGMENT|6092,6097|false|false|false|||palsy
Finding|Finding|SIMPLE_SEGMENT|6092,6097|false|false|false|C0522224;C3887651|Palsy;Paralysed|palsy
Finding|Body Substance|SIMPLE_SEGMENT|6102,6109|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6102,6109|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6102,6109|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|6114,6121|false|false|false|||resumed
Finding|Idea or Concept|SIMPLE_SEGMENT|6129,6133|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|6129,6133|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|6129,6133|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|6134,6146|false|false|false|C0249458|valacyclovir|Valacyclovir
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6134,6146|false|false|false|C0249458|valacyclovir|Valacyclovir
Event|Event|SIMPLE_SEGMENT|6134,6146|false|false|false|||Valacyclovir
Event|Event|SIMPLE_SEGMENT|6151,6162|false|false|false|||Prenisolone
Event|Event|SIMPLE_SEGMENT|6164,6168|false|false|false|||gtts
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6164,6168|false|false|false|C0017741|Glucose tolerance test|gtts
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6173,6180|false|false|false|C0042027|Urinary tract|Urinary
Finding|Sign or Symptom|SIMPLE_SEGMENT|6173,6188|false|false|false|C0085606|Urgency of micturition|Urinary urgency
Event|Event|SIMPLE_SEGMENT|6181,6188|false|false|false|||urgency
Finding|Body Substance|SIMPLE_SEGMENT|6203,6210|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6203,6210|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6203,6210|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|6211,6221|false|false|false|||complained
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6225,6232|false|false|false|C0042027|Urinary tract|urinary
Finding|Sign or Symptom|SIMPLE_SEGMENT|6225,6240|false|false|false|C0085606|Urgency of micturition|urinary urgency
Event|Event|SIMPLE_SEGMENT|6246,6255|false|false|false|||increased
Event|Event|SIMPLE_SEGMENT|6256,6265|false|false|false|||frequency
Finding|Intellectual Product|SIMPLE_SEGMENT|6256,6265|false|false|false|C3898838;C4321352|Frequency;How Often|frequency
Event|Event|SIMPLE_SEGMENT|6275,6283|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|6275,6283|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|6275,6283|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6275,6283|false|false|false|C5237010|Expression Negative|negative
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6288,6295|false|false|false|C1706355|Culture Dose Form|culture
Event|Event|SIMPLE_SEGMENT|6288,6295|false|false|false|||culture
Finding|Functional Concept|SIMPLE_SEGMENT|6288,6295|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Finding|Idea or Concept|SIMPLE_SEGMENT|6288,6295|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6288,6295|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|culture
Event|Event|SIMPLE_SEGMENT|6300,6308|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|6300,6308|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|6300,6308|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6300,6308|false|false|false|C5237010|Expression Negative|negative
Event|Event|SIMPLE_SEGMENT|6315,6323|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|6315,6323|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|6315,6323|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|SIMPLE_SEGMENT|6328,6336|false|false|false|||resolved
Finding|Finding|SIMPLE_SEGMENT|6344,6348|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|6344,6348|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|6344,6348|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|SIMPLE_SEGMENT|6352,6361|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|6352,6361|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6352,6361|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6352,6361|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6352,6361|false|false|false|C0030685|Patient Discharge|discharge
Finding|Body Substance|SIMPLE_SEGMENT|6376,6383|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6376,6383|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6376,6383|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|6388,6397|false|false|false|||evaluated
Event|Event|SIMPLE_SEGMENT|6416,6423|false|false|false|||cleared
Event|Event|SIMPLE_SEGMENT|6432,6436|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|6432,6436|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|6432,6436|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|6432,6436|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|6443,6451|false|false|false|||services
Event|Occupational Activity|SIMPLE_SEGMENT|6443,6451|false|false|false|C0557854|Services|services
Procedure|Health Care Activity|SIMPLE_SEGMENT|6443,6451|false|false|false|C1704289|Clinical Service|services
Event|Event|SIMPLE_SEGMENT|6461,6471|false|false|false|||discharged
Finding|Intellectual Product|SIMPLE_SEGMENT|6482,6488|false|false|false|C1547311|Patient Condition Code - Stable|stable
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6489,6498|false|false|false|C3864998||condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6489,6498|false|false|false|C0012634|Disease|condition
Event|Event|SIMPLE_SEGMENT|6489,6498|false|false|false|||condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|6489,6498|false|false|false|C1705253|Logical Condition|condition
Event|Event|SIMPLE_SEGMENT|6510,6516|false|false|false|||follow
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6538,6549|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6538,6549|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|6538,6549|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|6538,6549|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|6538,6562|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|SIMPLE_SEGMENT|6553,6562|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|6553,6562|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6566,6569|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Enzyme|SIMPLE_SEGMENT|6566,6569|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Organic Chemical|SIMPLE_SEGMENT|6566,6569|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6566,6569|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Event|Event|SIMPLE_SEGMENT|6566,6569|false|false|false|||ASA
Finding|Gene or Genome|SIMPLE_SEGMENT|6566,6569|false|false|false|C1412553|ARSA gene|ASA
Drug|Organic Chemical|SIMPLE_SEGMENT|6577,6588|false|false|false|C0102118|alendronate|Alendronate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6577,6588|false|false|false|C0102118|alendronate|Alendronate
Drug|Organic Chemical|SIMPLE_SEGMENT|6603,6610|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6603,6610|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|SIMPLE_SEGMENT|6603,6610|false|false|false|C0042890|Vitamins|Vitamin
Drug|Organic Chemical|SIMPLE_SEGMENT|6603,6613|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|Vitamin D3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6603,6613|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|Vitamin D3
Drug|Vitamin|SIMPLE_SEGMENT|6603,6613|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|Vitamin D3
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6632,6645|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Hormone|SIMPLE_SEGMENT|6632,6645|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Organic Chemical|SIMPLE_SEGMENT|6632,6645|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6632,6645|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6660,6670|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6660,6670|false|false|false|C0065374|lisinopril|Lisinopril
Event|Event|SIMPLE_SEGMENT|6685,6694|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|6685,6694|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6685,6694|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6685,6694|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6685,6694|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|6685,6706|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6695,6706|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6695,6706|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|6695,6706|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|6695,6706|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|6712,6725|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6712,6725|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|SIMPLE_SEGMENT|6712,6725|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6712,6725|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|SIMPLE_SEGMENT|6740,6743|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6744,6748|false|false|false|C2598155||Pain
Event|Event|SIMPLE_SEGMENT|6744,6748|false|false|false|||Pain
Finding|Functional Concept|SIMPLE_SEGMENT|6744,6748|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6744,6748|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Intellectual Product|SIMPLE_SEGMENT|6751,6755|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Finding|Finding|SIMPLE_SEGMENT|6756,6761|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|6756,6761|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Drug|Organic Chemical|SIMPLE_SEGMENT|6768,6777|false|false|false|C0005632|bisacodyl|Bisacodyl
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6768,6777|false|false|false|C0005632|bisacodyl|Bisacodyl
Drug|Organic Chemical|SIMPLE_SEGMENT|6802,6815|false|false|false|C0011777|dexamethasone|Dexamethasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6802,6815|false|false|false|C0011777|dexamethasone|Dexamethasone
Event|Event|SIMPLE_SEGMENT|6802,6815|false|false|false|||Dexamethasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6828,6836|false|false|false|C0720099|Duration brand of oxymetazoline|Duration
Event|Event|SIMPLE_SEGMENT|6828,6836|false|false|false|||Duration
Event|Event|SIMPLE_SEGMENT|6847,6852|false|false|false|||start
Event|Event|SIMPLE_SEGMENT|6873,6883|false|false|false|||2tabsq8hrs
Event|Event|SIMPLE_SEGMENT|6888,6899|false|false|false|||2tabsq12hrs
Event|Activity|SIMPLE_SEGMENT|6901,6912|false|false|false|C0024501|Maintenance|maintenance
Event|Event|SIMPLE_SEGMENT|6913,6917|false|false|false|||dose
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6929,6935|false|false|false|C1114758||dose #
Event|Event|SIMPLE_SEGMENT|6951,6956|false|false|false|||doses
Event|Event|SIMPLE_SEGMENT|6957,6959|false|false|false|||RX
Drug|Organic Chemical|SIMPLE_SEGMENT|6961,6974|false|false|false|C0011777|dexamethasone|dexamethasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6961,6974|false|false|false|C0011777|dexamethasone|dexamethasone
Event|Event|SIMPLE_SEGMENT|6961,6974|false|false|false|||dexamethasone
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6982,6988|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|SIMPLE_SEGMENT|6992,7000|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6995,7000|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6995,7000|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7035,7041|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|7042,7049|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|7042,7049|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|7058,7066|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7058,7066|false|false|false|C1692318|docusate|Docusate
Event|Event|SIMPLE_SEGMENT|7058,7066|false|false|false|||Docusate
Drug|Organic Chemical|SIMPLE_SEGMENT|7058,7073|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7058,7073|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7067,7073|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7067,7073|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7067,7073|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|7067,7073|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|7067,7073|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7067,7073|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7084,7087|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7084,7087|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7084,7087|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|7084,7087|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|7084,7087|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|7094,7104|false|false|false|C0015620|famotidine|Famotidine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7094,7104|false|false|false|C0015620|famotidine|Famotidine
Drug|Organic Chemical|SIMPLE_SEGMENT|7124,7134|false|false|false|C0015620|famotidine|famotidine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7124,7134|false|false|false|C0015620|famotidine|famotidine
Event|Event|SIMPLE_SEGMENT|7124,7134|false|false|false|||famotidine
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7143,7149|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|SIMPLE_SEGMENT|7153,7161|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7156,7161|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|7156,7161|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|SIMPLE_SEGMENT|7170,7173|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|7170,7173|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7185,7191|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|7192,7199|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|7192,7199|false|false|false|C0807726|refill|Refills
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7208,7220|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Drug|Organic Chemical|SIMPLE_SEGMENT|7208,7220|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Event|Event|SIMPLE_SEGMENT|7208,7220|false|false|false|||Polyethylene
Drug|Organic Chemical|SIMPLE_SEGMENT|7208,7227|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7208,7227|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|7221,7227|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Drug|Organic Chemical|SIMPLE_SEGMENT|7221,7227|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Event|Event|SIMPLE_SEGMENT|7221,7227|false|false|false|||Glycol
Finding|Gene or Genome|SIMPLE_SEGMENT|7242,7245|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|7246,7258|false|false|false|||Constipation
Finding|Sign or Symptom|SIMPLE_SEGMENT|7246,7258|false|false|false|C0009806|Constipation|Constipation
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7268,7272|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|7268,7272|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Drug|Substance|SIMPLE_SEGMENT|7268,7272|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Finding|Intellectual Product|SIMPLE_SEGMENT|7268,7272|false|false|false|C1546701|line source specimen code|Line
Drug|Organic Chemical|SIMPLE_SEGMENT|7279,7284|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7279,7284|false|false|false|C3489575|sennosides, USP|Senna
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7305,7318|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Hormone|SIMPLE_SEGMENT|7305,7318|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Organic Chemical|SIMPLE_SEGMENT|7305,7318|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7305,7318|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7305,7325|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Hormone|SIMPLE_SEGMENT|7305,7325|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7305,7325|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7319,7325|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7319,7325|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7319,7325|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|7319,7325|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|7319,7325|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7319,7325|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7348,7358|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7348,7358|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Organic Chemical|SIMPLE_SEGMENT|7381,7393|false|false|false|C0032950|prednisolone|PrednisoLONE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7381,7393|false|false|false|C0032950|prednisolone|PrednisoLONE
Drug|Organic Chemical|SIMPLE_SEGMENT|7381,7401|false|false|false|C0071839|prednisolone acetate|PrednisoLONE Acetate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7381,7401|false|false|false|C0071839|prednisolone acetate|PrednisoLONE Acetate
Drug|Organic Chemical|SIMPLE_SEGMENT|7394,7401|false|false|false|C0000975|acetate|Acetate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7394,7401|false|false|false|C0000975|acetate|Acetate
Finding|Functional Concept|SIMPLE_SEGMENT|7405,7410|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7420,7424|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|SIMPLE_SEGMENT|7420,7424|false|false|false|C1705648|Dropping|DROP
Event|Event|SIMPLE_SEGMENT|7425,7429|false|false|false|||LEFT
Finding|Functional Concept|SIMPLE_SEGMENT|7425,7429|false|false|false|C1552822|Table Cell Horizontal Align - left|LEFT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7425,7433|false|false|false|C0229090|Left eye structure|LEFT EYE
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7425,7433|false|false|false|C2141124|examination of left eye|LEFT EYE
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7430,7433|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|EYE
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7430,7433|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|EYE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7430,7433|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|EYE
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7430,7433|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|EYE
Event|Event|SIMPLE_SEGMENT|7430,7433|false|false|false|||EYE
Finding|Body Substance|SIMPLE_SEGMENT|7430,7433|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Finding|Finding|SIMPLE_SEGMENT|7430,7433|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Finding|Intellectual Product|SIMPLE_SEGMENT|7430,7433|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Drug|Organic Chemical|SIMPLE_SEGMENT|7445,7457|false|false|false|C0249458|valacyclovir|ValACYclovir
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7445,7457|false|false|false|C0249458|valacyclovir|ValACYclovir
Drug|Organic Chemical|SIMPLE_SEGMENT|7480,7487|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7480,7487|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|SIMPLE_SEGMENT|7480,7487|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|SIMPLE_SEGMENT|7480,7489|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|SIMPLE_SEGMENT|7480,7489|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7480,7489|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|SIMPLE_SEGMENT|7480,7489|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7480,7489|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|SIMPLE_SEGMENT|7488,7489|false|false|false|||D
Event|Event|SIMPLE_SEGMENT|7494,7498|false|false|false|||UNIT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7514,7518|false|false|false|C0675390|ARID1A protein, human|HELD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7514,7518|false|false|false|C0675390|ARID1A protein, human|HELD
Event|Event|SIMPLE_SEGMENT|7514,7518|false|false|false|||HELD
Finding|Gene or Genome|SIMPLE_SEGMENT|7514,7518|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|HELD
Finding|Idea or Concept|SIMPLE_SEGMENT|7514,7518|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|HELD
Drug|Organic Chemical|SIMPLE_SEGMENT|7520,7531|false|false|false|C0102118|alendronate|Alendronate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7520,7531|false|false|false|C0102118|alendronate|Alendronate
Drug|Organic Chemical|SIMPLE_SEGMENT|7520,7538|false|false|false|C0700482|alendronate sodium|Alendronate Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7520,7538|false|false|false|C0700482|alendronate sodium|Alendronate Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7532,7538|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7532,7538|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7532,7538|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|7532,7538|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|7532,7538|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7532,7538|false|false|false|C0337443|Sodium measurement|Sodium
Finding|Intellectual Product|SIMPLE_SEGMENT|7551,7555|false|false|false|C1561540|Transaction counts and value totals - week|WEEK
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7569,7579|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|7569,7579|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|7569,7579|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|7584,7588|false|false|false|||held
Event|Event|SIMPLE_SEGMENT|7597,7604|false|false|false|||restart
Drug|Organic Chemical|SIMPLE_SEGMENT|7605,7616|false|false|false|C0102118|alendronate|Alendronate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7605,7616|false|false|false|C0102118|alendronate|Alendronate
Drug|Organic Chemical|SIMPLE_SEGMENT|7605,7623|false|false|false|C0700482|alendronate sodium|Alendronate Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7605,7623|false|false|false|C0700482|alendronate sodium|Alendronate Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7617,7623|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7617,7623|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7617,7623|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|7617,7623|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|7617,7623|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7617,7623|false|false|false|C0337443|Sodium measurement|Sodium
Event|Event|SIMPLE_SEGMENT|7630,7633|false|false|false|||POD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7649,7653|false|false|false|C0675390|ARID1A protein, human|HELD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7649,7653|false|false|false|C0675390|ARID1A protein, human|HELD
Event|Event|SIMPLE_SEGMENT|7649,7653|false|false|false|||HELD
Finding|Gene or Genome|SIMPLE_SEGMENT|7649,7653|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|HELD
Finding|Idea or Concept|SIMPLE_SEGMENT|7649,7653|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|HELD
Drug|Organic Chemical|SIMPLE_SEGMENT|7655,7662|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7655,7662|false|false|false|C0004057|aspirin|Aspirin
Event|Event|SIMPLE_SEGMENT|7655,7662|false|false|false|||Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7684,7694|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|7684,7694|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|7684,7694|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|7699,7703|false|false|false|||held
Event|Event|SIMPLE_SEGMENT|7713,7720|false|false|false|||restart
Drug|Organic Chemical|SIMPLE_SEGMENT|7721,7728|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7721,7728|false|false|false|C0004057|aspirin|Aspirin
Event|Event|SIMPLE_SEGMENT|7721,7728|false|false|false|||Aspirin
Event|Event|SIMPLE_SEGMENT|7735,7738|false|false|false|||POD
Event|Event|SIMPLE_SEGMENT|7752,7762|false|false|false|||glucometer
Event|Event|SIMPLE_SEGMENT|7789,7794|false|false|false|||Check
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7795,7800|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|7795,7800|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|7795,7800|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Organic Chemical|SIMPLE_SEGMENT|7795,7807|false|false|false|C0005802|Blood Glucose|blood sugars
Drug|Organic Chemical|SIMPLE_SEGMENT|7801,7807|false|false|false|C0242209|Sugars|sugars
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7801,7807|false|false|false|C0242209|Sugars|sugars
Event|Event|SIMPLE_SEGMENT|7801,7807|false|false|false|||sugars
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7801,7807|false|false|false|C2239291|sugars (lab test)|sugars
Event|Event|SIMPLE_SEGMENT|7809,7810|false|false|false|||_
Event|Event|SIMPLE_SEGMENT|7835,7839|false|false|false|||meal
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|7835,7839|false|false|false|C1998602|Meal (occasion for eating)|meal
Finding|Intellectual Product|SIMPLE_SEGMENT|7841,7847|false|false|false|C0034869|Records|Record
Event|Event|SIMPLE_SEGMENT|7860,7864|false|false|false|||show
Event|Event|SIMPLE_SEGMENT|7873,7883|false|false|false|||Oncologist
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7890,7894|false|false|false|C4318744|Test - temporal region|test
Finding|Functional Concept|SIMPLE_SEGMENT|7890,7894|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|SIMPLE_SEGMENT|7890,7894|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7890,7894|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7890,7894|false|false|false|C0022885|Laboratory Procedures|test
Event|Event|SIMPLE_SEGMENT|7895,7901|false|false|false|||strips
Event|Event|SIMPLE_SEGMENT|7907,7912|false|false|false|||Check
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7913,7918|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|7913,7918|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|7913,7918|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Organic Chemical|SIMPLE_SEGMENT|7913,7925|false|false|false|C0005802|Blood Glucose|blood sugars
Drug|Organic Chemical|SIMPLE_SEGMENT|7919,7925|false|false|false|C0242209|Sugars|sugars
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7919,7925|false|false|false|C0242209|Sugars|sugars
Event|Event|SIMPLE_SEGMENT|7919,7925|false|false|false|||sugars
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7919,7925|false|false|false|C2239291|sugars (lab test)|sugars
Event|Event|SIMPLE_SEGMENT|7932,7939|false|false|false|||refills
Finding|Idea or Concept|SIMPLE_SEGMENT|7932,7939|false|false|false|C0807726|refill|refills
Event|Event|SIMPLE_SEGMENT|7960,7965|false|false|false|||Check
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7966,7971|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|7966,7971|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|7966,7971|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Organic Chemical|SIMPLE_SEGMENT|7966,7978|false|false|false|C0005802|Blood Glucose|blood sugars
Drug|Organic Chemical|SIMPLE_SEGMENT|7972,7978|false|false|false|C0242209|Sugars|sugars
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7972,7978|false|false|false|C0242209|Sugars|sugars
Event|Event|SIMPLE_SEGMENT|7972,7978|false|false|false|||sugars
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7972,7978|false|false|false|C2239291|sugars (lab test)|sugars
Event|Event|SIMPLE_SEGMENT|7985,7992|false|false|false|||refills
Finding|Idea or Concept|SIMPLE_SEGMENT|7985,7992|false|false|false|C0807726|refill|refills
Event|Event|SIMPLE_SEGMENT|7998,8007|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|7998,8007|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|7998,8007|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|7998,8007|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|7998,8007|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7998,8019|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|7998,8019|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8008,8019|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|8008,8019|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|8008,8019|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|SIMPLE_SEGMENT|8021,8025|false|false|false|||Home
Finding|Idea or Concept|SIMPLE_SEGMENT|8021,8025|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|8021,8025|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|8021,8025|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|SIMPLE_SEGMENT|8031,8038|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|8031,8038|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|SIMPLE_SEGMENT|8041,8049|false|false|false|||Facility
Finding|Intellectual Product|SIMPLE_SEGMENT|8041,8049|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|SIMPLE_SEGMENT|8057,8066|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|8057,8066|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8057,8066|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8057,8066|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8057,8066|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|8057,8076|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8067,8076|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|8067,8076|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|8067,8076|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|8067,8076|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8067,8076|false|false|false|C0011900|Diagnosis|Diagnosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8078,8083|false|false|false|C0006104;C4266577|Brain;Head>Brain|Brain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8078,8083|false|false|false|C0006111|Brain Diseases|Brain
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8078,8089|false|false|false|C0006118|Brain Neoplasms|Brain tumor
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8084,8089|false|false|false|C0027651|Neoplasms|tumor
Event|Event|SIMPLE_SEGMENT|8084,8089|false|false|false|||tumor
Finding|Finding|SIMPLE_SEGMENT|8084,8089|false|false|false|C1578706;C3273930|Tumor Mass|tumor
Finding|Intellectual Product|SIMPLE_SEGMENT|8084,8089|false|false|false|C1578706;C3273930|Tumor Mass|tumor
Event|Event|SIMPLE_SEGMENT|8093,8102|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|8093,8102|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8093,8102|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8093,8102|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8093,8102|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8103,8112|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8103,8112|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|8103,8112|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|8103,8112|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|8114,8120|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8114,8127|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|8114,8127|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8121,8127|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|8121,8127|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|8129,8134|false|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|8129,8134|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|8139,8147|false|false|false|||coherent
Finding|Finding|SIMPLE_SEGMENT|8139,8147|false|false|false|C4068804|Coherent|coherent
Event|Event|SIMPLE_SEGMENT|8149,8154|false|false|false|||Level
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8149,8171|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|8149,8171|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|SIMPLE_SEGMENT|8158,8171|false|false|false|||Consciousness
Finding|Finding|SIMPLE_SEGMENT|8158,8171|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|8158,8171|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8173,8178|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|8173,8178|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8173,8178|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|8173,8178|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|8173,8178|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|8173,8178|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|8173,8178|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|8183,8194|false|false|false|||interactive
Finding|Functional Concept|SIMPLE_SEGMENT|8183,8194|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|8196,8204|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|8196,8204|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|8196,8204|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8205,8211|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|8205,8211|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|8205,8211|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|SIMPLE_SEGMENT|8213,8223|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|8213,8223|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|8213,8223|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|8213,8223|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|SIMPLE_SEGMENT|8226,8234|false|false|false|||requires
Event|Event|SIMPLE_SEGMENT|8235,8245|false|false|false|||assistance
Finding|Social Behavior|SIMPLE_SEGMENT|8235,8245|false|false|false|C0018896|Helping Behavior|assistance
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8249,8252|false|false|false|C1454018|AICDA protein, human|aid
Drug|Enzyme|SIMPLE_SEGMENT|8249,8252|false|false|false|C1454018|AICDA protein, human|aid
Event|Event|SIMPLE_SEGMENT|8249,8252|false|false|false|||aid
Finding|Gene or Genome|SIMPLE_SEGMENT|8249,8252|false|false|false|C1421876;C3540469|AICDA gene;AICDA wt Allele|aid
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8249,8252|false|false|false|C0021588;C0280108|AID - Artificial insemination by donor;dacarbazine/doxorubicin/ifosfamide protocol|aid
Event|Event|SIMPLE_SEGMENT|8257,8266|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|8257,8266|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8257,8266|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8257,8266|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8257,8266|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8257,8279|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|8257,8279|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|8257,8279|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8267,8279|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|8267,8279|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|8267,8279|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Finding|Finding|SIMPLE_SEGMENT|8281,8288|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Finding|Functional Concept|SIMPLE_SEGMENT|8281,8288|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|8281,8288|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8281,8288|false|false|false|C0543467|Operative Surgical Procedures|Surgery
Event|Event|SIMPLE_SEGMENT|8307,8314|false|false|false|||surgery
Finding|Finding|SIMPLE_SEGMENT|8307,8314|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|8307,8314|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|8307,8314|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8307,8314|false|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Event|SIMPLE_SEGMENT|8318,8324|false|false|false|||remove
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8327,8332|false|false|false|C0006104;C4266577|Brain;Head>Brain|brain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8327,8332|false|false|false|C0006111|Brain Diseases|brain
Finding|Finding|SIMPLE_SEGMENT|8327,8339|false|false|false|C0221505|Lesion of brain|brain lesion
Event|Event|SIMPLE_SEGMENT|8333,8339|false|false|false|||lesion
Finding|Finding|SIMPLE_SEGMENT|8333,8339|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|SIMPLE_SEGMENT|8333,8339|false|false|false|C0221198;C1546698|Lesion|lesion
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8351,8356|false|false|false|C0006104;C4266577|Brain;Head>Brain|brain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8351,8356|false|false|false|C0006111|Brain Diseases|brain
Event|Event|SIMPLE_SEGMENT|8351,8356|false|false|false|||brain
Drug|Substance|SIMPLE_SEGMENT|8364,8370|false|false|false|C0370003|Specimen|sample
Event|Event|SIMPLE_SEGMENT|8364,8370|false|false|false|||sample
Finding|Body Substance|SIMPLE_SEGMENT|8364,8370|false|false|false|C2347026;C5551027|Biospecimen;Nucleotide Sequence Sample Name|sample
Finding|Intellectual Product|SIMPLE_SEGMENT|8364,8370|false|false|false|C2347026;C5551027|Biospecimen;Nucleotide Sequence Sample Name|sample
Anatomy|Tissue|SIMPLE_SEGMENT|8374,8380|false|false|false|C0040300|Body tissue|tissue
Finding|Intellectual Product|SIMPLE_SEGMENT|8374,8380|false|false|false|C1547928|Tissue Specimen Code|tissue
Event|Event|SIMPLE_SEGMENT|8390,8396|false|false|false|||lesion
Finding|Finding|SIMPLE_SEGMENT|8390,8396|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|SIMPLE_SEGMENT|8390,8396|false|false|false|C0221198;C1546698|Lesion|lesion
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8405,8410|false|false|false|C0006104;C4266577|Brain;Head>Brain|brain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8405,8410|false|false|false|C0006111|Brain Diseases|brain
Event|Event|SIMPLE_SEGMENT|8415,8419|false|false|false|||sent
Event|Event|SIMPLE_SEGMENT|8424,8433|false|false|false|||pathology
Finding|Functional Concept|SIMPLE_SEGMENT|8424,8433|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Finding|Pathologic Function|SIMPLE_SEGMENT|8424,8433|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8424,8433|false|false|false|C0919386|Pathology procedure|pathology
Event|Event|SIMPLE_SEGMENT|8438,8445|false|false|false|||testing
Finding|Functional Concept|SIMPLE_SEGMENT|8438,8445|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|testing
Finding|Intellectual Product|SIMPLE_SEGMENT|8438,8445|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|testing
Event|Event|SIMPLE_SEGMENT|8458,8462|false|false|false|||keep
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8468,8476|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|8468,8476|false|false|false|C0332803|Surgical wound|incision
Event|Event|SIMPLE_SEGMENT|8468,8476|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8468,8476|false|false|false|C0184898|Surgical incisions|incision
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|8492,8499|false|false|false|C0502420|Suture Joint|sutures
Event|Event|SIMPLE_SEGMENT|8492,8499|false|false|false|||sutures
Event|Event|SIMPLE_SEGMENT|8504,8511|false|false|false|||removed
Event|Event|SIMPLE_SEGMENT|8525,8531|false|false|false|||shower
Finding|Finding|SIMPLE_SEGMENT|8540,8544|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|8540,8544|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|8540,8544|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8559,8567|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|8559,8567|false|false|false|C0332803|Surgical wound|incision
Event|Event|SIMPLE_SEGMENT|8559,8567|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8559,8567|false|false|false|C0184898|Surgical incisions|incision
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8582,8586|false|false|false|C0339510|Vitelliform Macular Dystrophy|best
Event|Event|SIMPLE_SEGMENT|8582,8586|false|false|false|||best
Finding|Gene or Genome|SIMPLE_SEGMENT|8582,8586|false|false|false|C1826421;C5781213|BEST1 gene;BEST1 wt Allele|best
Event|Event|SIMPLE_SEGMENT|8590,8594|false|false|false|||keep
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8600,8608|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|8600,8608|false|false|false|C0332803|Surgical wound|incision
Event|Event|SIMPLE_SEGMENT|8600,8608|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8600,8608|false|false|false|C0184898|Surgical incisions|incision
Event|Event|SIMPLE_SEGMENT|8609,8613|false|false|false|||open
Drug|Inorganic Chemical|SIMPLE_SEGMENT|8617,8620|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8617,8620|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|SIMPLE_SEGMENT|8617,8620|false|false|false|C0001861;C3536832|Air (substance);air|air
Event|Event|SIMPLE_SEGMENT|8617,8620|false|false|false|||air
Finding|Finding|SIMPLE_SEGMENT|8617,8620|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|SIMPLE_SEGMENT|8617,8620|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|SIMPLE_SEGMENT|8617,8620|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Event|Event|SIMPLE_SEGMENT|8638,8643|false|false|false|||cover
Event|Event|SIMPLE_SEGMENT|8665,8669|false|false|false|||Call
Finding|Functional Concept|SIMPLE_SEGMENT|8665,8669|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|Call
Finding|Gene or Genome|SIMPLE_SEGMENT|8665,8669|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|Call
Finding|Intellectual Product|SIMPLE_SEGMENT|8665,8669|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|Call
Finding|Mental Process|SIMPLE_SEGMENT|8665,8669|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|Call
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8675,8682|false|false|false|C5444295||surgeon
Event|Event|SIMPLE_SEGMENT|8700,8705|false|false|false|||signs
Finding|Finding|SIMPLE_SEGMENT|8700,8705|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|8700,8705|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8709,8718|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|8709,8718|false|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|8709,8718|false|false|false|C3714514|Infection|infection
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8725,8732|false|false|false|C0041834|Erythema|redness
Event|Event|SIMPLE_SEGMENT|8725,8732|false|false|false|||redness
Finding|Finding|SIMPLE_SEGMENT|8725,8732|false|false|false|C0332575|Redness|redness
Event|Event|SIMPLE_SEGMENT|8734,8739|false|false|false|||fever
Finding|Finding|SIMPLE_SEGMENT|8734,8739|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|8734,8739|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|SIMPLE_SEGMENT|8744,8752|false|false|false|||drainage
Finding|Body Substance|SIMPLE_SEGMENT|8744,8752|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|SIMPLE_SEGMENT|8744,8752|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8744,8752|false|false|false|C0013103|Drainage procedure|drainage
Event|Activity|SIMPLE_SEGMENT|8756,8764|false|false|false|C0441655|Activities|Activity
Event|Event|SIMPLE_SEGMENT|8756,8764|false|false|false|||Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|8756,8764|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|8756,8764|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Event|Event|SIMPLE_SEGMENT|8772,8781|false|false|false|||recommend
Event|Event|SIMPLE_SEGMENT|8791,8796|false|false|false|||avoid
Event|Activity|SIMPLE_SEGMENT|8803,8810|false|false|false|C0206244|Lifting|lifting
Event|Event|SIMPLE_SEGMENT|8803,8810|false|false|false|||lifting
Event|Event|SIMPLE_SEGMENT|8812,8819|false|false|false|||running
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|8812,8819|false|false|false|C0035953;C2346414;C4722187|Go Jogging or Running Question;Running (physical activity);running (history)|running
Finding|Finding|SIMPLE_SEGMENT|8812,8819|false|false|false|C0035953;C2346414;C4722187|Go Jogging or Running Question;Running (physical activity);running (history)|running
Finding|Intellectual Product|SIMPLE_SEGMENT|8812,8819|false|false|false|C0035953;C2346414;C4722187|Go Jogging or Running Question;Running (physical activity);running (history)|running
Event|Event|SIMPLE_SEGMENT|8821,8829|false|false|false|||climbing
Finding|Finding|SIMPLE_SEGMENT|8821,8829|false|false|false|C0561942;C2362653;C2584300|Climbing;Does climb;climbing (history)|climbing
Finding|Individual Behavior|SIMPLE_SEGMENT|8821,8829|false|false|false|C0561942;C2362653;C2584300|Climbing;Does climb;climbing (history)|climbing
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|8841,8859|false|false|false|C1514989|Strenuous Exercise|strenuous exercise
Event|Event|SIMPLE_SEGMENT|8851,8859|false|false|false|||exercise
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|8851,8859|false|false|false|C0015259|Exercise|exercise
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8851,8859|false|false|false|C1522704|Exercise Pain Management|exercise
Event|Event|SIMPLE_SEGMENT|8871,8877|false|false|false|||follow
Finding|Functional Concept|SIMPLE_SEGMENT|8871,8877|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|8871,8877|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|SIMPLE_SEGMENT|8871,8880|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|SIMPLE_SEGMENT|8871,8880|false|false|false|C1522577|follow-up|follow-up
Event|Activity|SIMPLE_SEGMENT|8881,8892|false|false|false|C0003629|Appointments|appointment
Event|Event|SIMPLE_SEGMENT|8881,8892|false|false|false|||appointment
Event|Event|SIMPLE_SEGMENT|8921,8926|false|false|false|||walks
Finding|Finding|SIMPLE_SEGMENT|8921,8926|false|false|false|C0600108|Does walk|walks
Event|Event|SIMPLE_SEGMENT|8938,8946|false|false|false|||increase
Event|Activity|SIMPLE_SEGMENT|8953,8961|false|false|false|C0441655|Activities|activity
Event|Event|SIMPLE_SEGMENT|8953,8961|false|false|false|||activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|8953,8961|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Finding|Finding|SIMPLE_SEGMENT|8953,8961|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Finding|Finding|SIMPLE_SEGMENT|8970,8973|false|false|false|C5939094|Own|own
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8974,8978|false|false|false|C0281567;C1310542;C4048252|FURIN protein, human;cisplatin/cyclophosphamide/doxorubicin/etoposide;cyclophosphamide/doxorubicin/etoposide/prednisone|pace
Drug|Enzyme|SIMPLE_SEGMENT|8974,8978|false|false|false|C0281567;C1310542;C4048252|FURIN protein, human;cisplatin/cyclophosphamide/doxorubicin/etoposide;cyclophosphamide/doxorubicin/etoposide/prednisone|pace
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8974,8978|false|false|false|C0281567;C1310542;C4048252|FURIN protein, human;cisplatin/cyclophosphamide/doxorubicin/etoposide;cyclophosphamide/doxorubicin/etoposide/prednisone|pace
Event|Event|SIMPLE_SEGMENT|8974,8978|false|false|false|||pace
Finding|Gene or Genome|SIMPLE_SEGMENT|8974,8978|false|false|false|C0919550;C1150256;C5444037|FURIN gene;Patient Assessment of Cancer Communication Experiences;furin activity|pace
Finding|Intellectual Product|SIMPLE_SEGMENT|8974,8978|false|false|false|C0919550;C1150256;C5444037|FURIN gene;Patient Assessment of Cancer Communication Experiences;furin activity|pace
Finding|Molecular Function|SIMPLE_SEGMENT|8974,8978|false|false|false|C0919550;C1150256;C5444037|FURIN gene;Patient Assessment of Cancer Communication Experiences;furin activity|pace
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8974,8978|false|false|false|C0280022|cisplatin/cyclophosphamide/doxorubicin/vindesine protocol|pace
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8992,8999|false|false|false|C3854129||symptom
Event|Event|SIMPLE_SEGMENT|8992,8999|false|false|false|||symptom
Finding|Sign or Symptom|SIMPLE_SEGMENT|8992,8999|false|false|false|C1457887|Symptoms|symptom
Event|Event|SIMPLE_SEGMENT|9000,9004|false|false|false|||free
Finding|Functional Concept|SIMPLE_SEGMENT|9000,9004|false|false|false|C0332296|Free of (attribute)|free
Finding|Functional Concept|SIMPLE_SEGMENT|9005,9012|false|false|false|C0443144|At rest (qualifier value)|at rest
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9008,9012|false|false|false|C1742913|REST protein, human|rest
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9008,9012|false|false|false|C1742913|REST protein, human|rest
Event|Event|SIMPLE_SEGMENT|9008,9012|false|false|false|||rest
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|9008,9012|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Gene or Genome|SIMPLE_SEGMENT|9008,9012|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Molecular Function|SIMPLE_SEGMENT|9008,9012|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Finding|SIMPLE_SEGMENT|9029,9037|false|false|false|C3843660|Too much|too much
Finding|Finding|SIMPLE_SEGMENT|9033,9037|false|false|false|C4281574|Much|much
Finding|Intellectual Product|SIMPLE_SEGMENT|9045,9049|false|false|false|C1720092|Once - dosing instruction fragment|once
Event|Event|SIMPLE_SEGMENT|9057,9064|false|false|false|||driving
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|9057,9064|false|false|false|C0004379|Automobile Driving|driving
Event|Event|SIMPLE_SEGMENT|9071,9077|false|false|false|||taking
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|9082,9090|true|false|false|C0027415|Narcotics|narcotic
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9082,9090|true|false|false|C0027415|Narcotics|narcotic
Event|Event|SIMPLE_SEGMENT|9082,9090|false|false|false|||narcotic
Event|Event|SIMPLE_SEGMENT|9094,9102|false|false|false|||sedating
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9103,9113|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|9103,9113|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|9103,9113|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|9140,9147|false|false|false|||seizure
Finding|Sign or Symptom|SIMPLE_SEGMENT|9140,9147|false|false|false|C0036572|Seizures|seizure
Event|Event|SIMPLE_SEGMENT|9154,9162|false|false|false|||admitted
Event|Event|SIMPLE_SEGMENT|9177,9184|false|false|false|||allowed
Event|Event|SIMPLE_SEGMENT|9188,9193|false|false|false|||drive
Finding|Intellectual Product|SIMPLE_SEGMENT|9197,9200|false|false|false|C1947938|Law (document)|law
Event|Activity|SIMPLE_SEGMENT|9209,9216|false|false|false|C3812666|Personal Contact|contact
Finding|Functional Concept|SIMPLE_SEGMENT|9209,9216|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|contact
Finding|Idea or Concept|SIMPLE_SEGMENT|9209,9216|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|contact
Finding|Intellectual Product|SIMPLE_SEGMENT|9209,9216|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|contact
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|9209,9216|false|false|false|C0392367|Physical contact|contact
Event|Event|SIMPLE_SEGMENT|9217,9223|false|false|false|||sports
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|9217,9223|false|false|false|C0038039|Sports|sports
Event|Event|SIMPLE_SEGMENT|9230,9237|false|false|false|||cleared
Event|Event|SIMPLE_SEGMENT|9246,9258|false|false|false|||neurosurgeon
Event|Activity|SIMPLE_SEGMENT|9278,9285|false|false|false|C3812666|Personal Contact|contact
Event|Event|SIMPLE_SEGMENT|9278,9285|false|false|false|||contact
Finding|Functional Concept|SIMPLE_SEGMENT|9278,9285|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|contact
Finding|Idea or Concept|SIMPLE_SEGMENT|9278,9285|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|contact
Finding|Intellectual Product|SIMPLE_SEGMENT|9278,9285|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|contact
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|9278,9285|false|false|false|C0392367|Physical contact|contact
Event|Event|SIMPLE_SEGMENT|9286,9292|false|false|false|||sports
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|9286,9292|false|false|false|C0038039|Sports|sports
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9309,9320|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9309,9320|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|9309,9320|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|9309,9320|false|false|false|C4284232|Medications|Medications
Event|Event|SIMPLE_SEGMENT|9339,9343|false|false|false|||take
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9348,9353|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|9348,9353|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|9348,9353|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Sign or Symptom|SIMPLE_SEGMENT|9354,9362|false|false|false|C0851184|Thinning Weight Loss|thinning
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9363,9373|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|9363,9373|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|9363,9373|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Drug|Organic Chemical|SIMPLE_SEGMENT|9375,9382|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9375,9382|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|9385,9394|false|false|false|C0020740|ibuprofen|Ibuprofen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9385,9394|false|false|false|C0020740|ibuprofen|Ibuprofen
Event|Event|SIMPLE_SEGMENT|9385,9394|false|false|false|||Ibuprofen
Drug|Organic Chemical|SIMPLE_SEGMENT|9396,9402|false|false|false|C0633084|Plavix|Plavix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9396,9402|false|false|false|C0633084|Plavix|Plavix
Event|Event|SIMPLE_SEGMENT|9396,9402|false|false|false|||Plavix
Drug|Organic Chemical|SIMPLE_SEGMENT|9404,9412|false|false|false|C0699129|Coumadin|Coumadin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9404,9412|false|false|false|C0699129|Coumadin|Coumadin
Event|Event|SIMPLE_SEGMENT|9404,9412|false|false|false|||Coumadin
Event|Event|SIMPLE_SEGMENT|9420,9427|false|false|false|||cleared
Event|Event|SIMPLE_SEGMENT|9453,9457|false|false|false|||held
Drug|Organic Chemical|SIMPLE_SEGMENT|9463,9470|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9463,9470|false|false|false|C0004057|aspirin|Aspirin
Event|Event|SIMPLE_SEGMENT|9491,9498|false|false|false|||cleared
Event|Event|SIMPLE_SEGMENT|9502,9508|false|false|false|||resume
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9515,9525|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|9515,9525|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|9515,9525|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|9529,9532|false|false|false|||POD
Event|Event|SIMPLE_SEGMENT|9550,9554|false|false|false|||held
Finding|Idea or Concept|SIMPLE_SEGMENT|9560,9564|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|9560,9564|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|9560,9564|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|9565,9576|false|false|false|C0102118|alendronate|Alendronate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9565,9576|false|false|false|C0102118|alendronate|Alendronate
Event|Event|SIMPLE_SEGMENT|9565,9576|false|false|false|||Alendronate
Event|Event|SIMPLE_SEGMENT|9589,9598|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|9589,9598|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|9609,9616|false|false|false|||cleared
Event|Event|SIMPLE_SEGMENT|9620,9626|false|false|false|||resume
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9632,9642|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|9632,9642|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|9632,9642|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|9646,9649|false|false|false|||POD
Event|Event|SIMPLE_SEGMENT|9672,9675|false|false|false|||use
Drug|Organic Chemical|SIMPLE_SEGMENT|9676,9689|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9676,9689|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|SIMPLE_SEGMENT|9676,9689|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9676,9689|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Organic Chemical|SIMPLE_SEGMENT|9691,9698|false|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9691,9698|false|false|false|C0699142|Tylenol|Tylenol
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9704,9709|false|false|false|C1446899|minor (disease)|minor
Event|Event|SIMPLE_SEGMENT|9704,9709|false|false|false|||minor
Finding|Gene or Genome|SIMPLE_SEGMENT|9704,9709|false|false|false|C1417837;C3272493|NR4A3 gene;NR4A3 wt Allele|minor
Event|Event|SIMPLE_SEGMENT|9710,9720|false|false|false|||discomfort
Finding|Sign or Symptom|SIMPLE_SEGMENT|9710,9720|false|false|false|C2364135|Discomfort|discomfort
Event|Event|SIMPLE_SEGMENT|9747,9757|false|false|false|||restricted
Event|Event|SIMPLE_SEGMENT|9763,9769|false|false|false|||taking
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9775,9785|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|9775,9785|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|9775,9785|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|9799,9806|false|false|false|||started
Drug|Organic Chemical|SIMPLE_SEGMENT|9810,9823|false|false|false|C0011777|dexamethasone|Dexamethasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9810,9823|false|false|false|C0011777|dexamethasone|Dexamethasone
Event|Event|SIMPLE_SEGMENT|9810,9823|false|false|false|||Dexamethasone
Drug|Organic Chemical|SIMPLE_SEGMENT|9827,9834|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9827,9834|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Event|Event|SIMPLE_SEGMENT|9827,9834|false|false|false|||steroid
Event|Event|SIMPLE_SEGMENT|9840,9846|false|false|false|||treats
Finding|Functional Concept|SIMPLE_SEGMENT|9840,9846|false|false|false|C1292734;C5966192|Intent To Treat;Treats (attribute)|treats
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9848,9860|false|false|false|C0524466|Intracranial|intracranial
Finding|Functional Concept|SIMPLE_SEGMENT|9848,9860|false|false|false|C1522213|Intracranial Route of Administration|intracranial
Finding|Pathologic Function|SIMPLE_SEGMENT|9848,9869|false|false|false|C1527311|Brain Edema|intracranial swelling
Event|Event|SIMPLE_SEGMENT|9861,9869|false|false|false|||swelling
Finding|Finding|SIMPLE_SEGMENT|9861,9869|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|9861,9869|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Drug|Organic Chemical|SIMPLE_SEGMENT|9876,9889|false|false|false|C0011777|dexamethasone|Dexamethasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9876,9889|false|false|false|C0011777|dexamethasone|Dexamethasone
Event|Event|SIMPLE_SEGMENT|9876,9889|false|false|false|||Dexamethasone
Event|Event|SIMPLE_SEGMENT|9899,9906|false|false|false|||tapered
Event|Activity|SIMPLE_SEGMENT|9918,9929|false|false|false|C0024501|Maintenance|maintenance
Event|Event|SIMPLE_SEGMENT|9930,9934|false|false|false|||dose
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9942,9945|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9942,9945|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9942,9945|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|9942,9945|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|9942,9945|false|false|false|C1332410|BID gene|BID
Event|Event|SIMPLE_SEGMENT|9954,9958|false|false|false|||take
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9964,9974|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|9964,9974|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|9964,9974|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|9979,9989|false|false|false|||prescribed
Event|Event|SIMPLE_SEGMENT|10000,10008|false|false|false|||admitted
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10018,10040|false|false|false|C0020456|Hyperglycemia|elevated blood glucose
Finding|Finding|SIMPLE_SEGMENT|10018,10040|false|false|false|C0595877;C2703060|Blood glucose increased;elevated random blood glucose level|elevated blood glucose
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10027,10032|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|10027,10032|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|10027,10032|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Organic Chemical|SIMPLE_SEGMENT|10027,10040|false|false|false|C0005802|Blood Glucose|blood glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|10027,10040|false|false|false|C0428554|Finding of blood glucose level|blood glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10027,10040|false|false|false|C0392201|Blood glucose measurement|blood glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|10027,10047|false|false|false|C0428554|Finding of blood glucose level|blood glucose levels
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10033,10040|false|false|false|C0017725|glucose|glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|10033,10040|false|false|false|C0017725|glucose|glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10033,10040|false|false|false|C0017725|glucose|glucose
Event|Event|SIMPLE_SEGMENT|10033,10040|false|false|false|||glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|10033,10040|false|false|false|C5781949|Glucose^1.5H post dose glucagon|glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10033,10040|false|false|false|C0337438|Glucose measurement|glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|10033,10047|false|false|false|C0428548||glucose levels
Event|Event|SIMPLE_SEGMENT|10041,10047|false|false|false|||levels
Event|Event|SIMPLE_SEGMENT|10054,10060|false|false|false|||needed
Event|Event|SIMPLE_SEGMENT|10067,10074|false|false|false|||treated
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10078,10085|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Hormone|SIMPLE_SEGMENT|10078,10085|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10078,10085|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Event|Event|SIMPLE_SEGMENT|10078,10085|false|false|false|||Insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|10078,10085|false|false|false|C1337112|INS gene|Insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10078,10085|false|false|false|C0202098|Insulin measurement|Insulin
Event|Event|SIMPLE_SEGMENT|10098,10106|false|false|false|||continue
Event|Activity|SIMPLE_SEGMENT|10110,10115|false|false|false|C1283174||check
Event|Event|SIMPLE_SEGMENT|10110,10115|false|false|false|||check
Finding|Functional Concept|SIMPLE_SEGMENT|10110,10115|false|false|false|C4321547|Check|check
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10122,10127|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|10122,10127|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|10122,10127|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Organic Chemical|SIMPLE_SEGMENT|10122,10134|false|false|false|C0005802|Blood Glucose|blood sugars
Drug|Organic Chemical|SIMPLE_SEGMENT|10128,10134|false|false|false|C0242209|Sugars|sugars
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10128,10134|false|false|false|C0242209|Sugars|sugars
Event|Event|SIMPLE_SEGMENT|10128,10134|false|false|false|||sugars
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10128,10134|false|false|false|C2239291|sugars (lab test)|sugars
Finding|Finding|SIMPLE_SEGMENT|10141,10148|false|false|false|C4534363|At home|at home
Event|Event|SIMPLE_SEGMENT|10144,10148|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|10144,10148|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|10144,10148|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|10144,10148|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|10169,10179|false|false|false|||glucometer
Event|Event|SIMPLE_SEGMENT|10208,10213|false|false|false|||teach
Event|Event|SIMPLE_SEGMENT|10225,10228|false|false|false|||use
Event|Event|SIMPLE_SEGMENT|10234,10240|false|false|false|||device
Finding|Functional Concept|SIMPLE_SEGMENT|10234,10240|false|false|false|C1550509|Participation Type - device|device
Event|Event|SIMPLE_SEGMENT|10245,10249|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|10245,10249|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|10245,10249|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|10245,10249|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|10258,10264|false|false|false|||record
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10270,10275|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|10270,10275|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|10270,10275|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Organic Chemical|SIMPLE_SEGMENT|10270,10282|false|false|false|C0005802|Blood Glucose|blood sugars
Drug|Organic Chemical|SIMPLE_SEGMENT|10276,10282|false|false|false|C0242209|Sugars|sugars
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10276,10282|false|false|false|C0242209|Sugars|sugars
Event|Event|SIMPLE_SEGMENT|10276,10282|false|false|false|||sugars
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10276,10282|false|false|false|C2239291|sugars (lab test)|sugars
Event|Event|SIMPLE_SEGMENT|10287,10293|false|false|false|||follow
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10308,10311|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|10308,10311|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|10308,10311|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10308,10311|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|10308,10311|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|10308,10311|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|10308,10311|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10308,10311|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|10308,10311|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|10308,10311|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|10308,10311|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|SIMPLE_SEGMENT|10348,10352|false|false|false|||goal
Finding|Idea or Concept|SIMPLE_SEGMENT|10348,10352|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Finding|Intellectual Product|SIMPLE_SEGMENT|10348,10352|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10353,10358|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|10353,10358|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|10353,10358|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Organic Chemical|SIMPLE_SEGMENT|10353,10364|false|false|false|C0005802|Blood Glucose|blood sugar
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10353,10364|false|false|false|C0392201|Blood glucose measurement|blood sugar
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10359,10364|false|false|false|C0007004;C0242209;C3665462|Carbohydrates;Sugars;raw sugar|sugar
Drug|Organic Chemical|SIMPLE_SEGMENT|10359,10364|false|false|false|C0007004;C0242209;C3665462|Carbohydrates;Sugars;raw sugar|sugar
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10359,10364|false|false|false|C0007004;C0242209;C3665462|Carbohydrates;Sugars;raw sugar|sugar
Event|Event|SIMPLE_SEGMENT|10359,10364|false|false|false|||sugar
Finding|Mental Process|SIMPLE_SEGMENT|10399,10409|false|false|false|C0237607;C0596545|Experience;Experience (Practice)|Experience
Event|Event|SIMPLE_SEGMENT|10433,10442|false|false|false|||headaches
Finding|Sign or Symptom|SIMPLE_SEGMENT|10433,10442|false|false|false|C0018681|Headache|headaches
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10447,10457|false|false|false|C0184898|Surgical incisions|incisional
Finding|Sign or Symptom|SIMPLE_SEGMENT|10447,10462|false|false|false|C1717947|Incisional pain|incisional pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10458,10462|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|10458,10462|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|10458,10462|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|10458,10462|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|10481,10491|false|false|false|||experience
Finding|Finding|SIMPLE_SEGMENT|10512,10520|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|10512,10520|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Event|Event|SIMPLE_SEGMENT|10521,10527|false|false|false|||around
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10534,10538|false|false|false|C0015450;C4266571|Face;Head>Face|face
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10534,10538|false|false|false|C3160739|FANCONI ANEMIA, COMPLEMENTATION GROUP E|face
Event|Event|SIMPLE_SEGMENT|10534,10538|false|false|false|||face
Finding|Gene or Genome|SIMPLE_SEGMENT|10534,10538|false|false|false|C1414531;C1423759;C2828055|ELOVL6 gene;FANCE gene;FANCE wt Allele|face
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10543,10547|false|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10543,10547|false|false|false|C5848506||eyes
Event|Event|SIMPLE_SEGMENT|10557,10563|false|false|false|||normal
Finding|Finding|SIMPLE_SEGMENT|10564,10577|false|false|false|C0241311|post operative (finding)|after surgery
Event|Event|SIMPLE_SEGMENT|10570,10577|false|false|false|||surgery
Finding|Finding|SIMPLE_SEGMENT|10570,10577|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|10570,10577|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|10570,10577|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10570,10577|false|false|false|C0543467|Operative Surgical Procedures|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|10606,10612|false|false|false|C1522484;C1561503;C1705190|Precision - second;Second Suffix;metastatic qualifier|second
Finding|Idea or Concept|SIMPLE_SEGMENT|10606,10612|false|false|false|C1522484;C1561503;C1705190|Precision - second;Second Suffix;metastatic qualifier|second
Finding|Intellectual Product|SIMPLE_SEGMENT|10606,10612|false|false|false|C1522484;C1561503;C1705190|Precision - second;Second Suffix;metastatic qualifier|second
Finding|Idea or Concept|SIMPLE_SEGMENT|10623,10626|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|10623,10626|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|10630,10637|false|false|false|||surgery
Finding|Finding|SIMPLE_SEGMENT|10630,10637|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|10630,10637|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|10630,10637|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10630,10637|false|false|false|C0543467|Operative Surgical Procedures|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|10644,10649|false|false|false|C1632850;C1879355;C4048755;C4521676|Apply;Apply (administration method);Apply (instruction)|apply
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10651,10654|false|false|false|C0228434;C3496566|Structure of inferior central nucleus of pons;intracentral fissure|ice
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|10651,10654|false|false|false|C0228434;C3496566|Structure of inferior central nucleus of pons;intracentral fissure|ice
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10651,10654|false|false|false|C0020746;C0025611;C1873773;C4721557|Caspase-1, human;Ice;Ice Pharmaceutical;methamphetamine|ice
Drug|Enzyme|SIMPLE_SEGMENT|10651,10654|false|false|false|C0020746;C0025611;C1873773;C4721557|Caspase-1, human;Ice;Ice Pharmaceutical;methamphetamine|ice
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|10651,10654|false|false|false|C0020746;C0025611;C1873773;C4721557|Caspase-1, human;Ice;Ice Pharmaceutical;methamphetamine|ice
Drug|Inorganic Chemical|SIMPLE_SEGMENT|10651,10654|false|false|false|C0020746;C0025611;C1873773;C4721557|Caspase-1, human;Ice;Ice Pharmaceutical;methamphetamine|ice
Drug|Organic Chemical|SIMPLE_SEGMENT|10651,10654|false|false|false|C0020746;C0025611;C1873773;C4721557|Caspase-1, human;Ice;Ice Pharmaceutical;methamphetamine|ice
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10651,10654|false|false|false|C0020746;C0025611;C1873773;C4721557|Caspase-1, human;Ice;Ice Pharmaceutical;methamphetamine|ice
Event|Event|SIMPLE_SEGMENT|10651,10654|false|false|false|||ice
Finding|Gene or Genome|SIMPLE_SEGMENT|10651,10654|false|false|false|C1150137;C1366479;C1413348;C1705786;C3889432|CASP1 gene;CASP1 wt Allele;CES2 gene;CES2 wt Allele;caspase-1 activity|ice
Finding|Molecular Function|SIMPLE_SEGMENT|10651,10654|false|false|false|C1150137;C1366479;C1413348;C1705786;C3889432|CASP1 gene;CASP1 wt Allele;CES2 gene;CES2 wt Allele;caspase-1 activity|ice
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10651,10654|false|false|false|C0249492;C0280697;C0556917;C1879508|AIE Regimen;carboplatin/etoposide/ifosfamide;cryotherapy using ice;cytarabine/etoposide/idarubicin|ice
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|10660,10664|false|false|false|C0678568||cool
Event|Event|SIMPLE_SEGMENT|10668,10672|false|false|false|||warm
Finding|Finding|SIMPLE_SEGMENT|10668,10672|false|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|10668,10672|false|false|false|C0687712|warming process|warm
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10691,10695|false|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10691,10695|false|false|false|C5848506||eyes
Event|Event|SIMPLE_SEGMENT|10699,10703|false|false|false|||help
Event|Event|SIMPLE_SEGMENT|10714,10722|false|false|false|||swelling
Finding|Finding|SIMPLE_SEGMENT|10714,10722|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|10714,10722|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Event|Event|SIMPLE_SEGMENT|10728,10736|false|false|false|||swelling
Finding|Finding|SIMPLE_SEGMENT|10728,10736|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|10728,10736|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Event|Event|SIMPLE_SEGMENT|10749,10754|false|false|false|||worse
Finding|Finding|SIMPLE_SEGMENT|10749,10754|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Idea or Concept|SIMPLE_SEGMENT|10749,10754|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Drug|Organic Chemical|SIMPLE_SEGMENT|10762,10775|false|false|false|C4019028|Morning After|morning after
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10762,10775|false|false|false|C4019028|Morning After|morning after
Event|Event|SIMPLE_SEGMENT|10770,10775|false|false|false|||after
Event|Event|SIMPLE_SEGMENT|10777,10783|false|false|false|||laying
Event|Event|SIMPLE_SEGMENT|10794,10802|false|false|false|||sleeping
Event|Event|SIMPLE_SEGMENT|10807,10815|false|false|false|||decrease
Event|Event|SIMPLE_SEGMENT|10837,10847|false|false|false|||experience
Event|Event|SIMPLE_SEGMENT|10848,10856|false|false|false|||soreness
Finding|Sign or Symptom|SIMPLE_SEGMENT|10848,10856|false|false|false|C0234233|Sore to touch|soreness
Event|Event|SIMPLE_SEGMENT|10862,10869|false|false|false|||chewing
Finding|Finding|SIMPLE_SEGMENT|10862,10869|false|false|false|C0024888;C2015927|Chewing;outcomes otolaryngology chewing|chewing
Finding|Organism Function|SIMPLE_SEGMENT|10862,10869|false|false|false|C0024888;C2015927|Chewing;outcomes otolaryngology chewing|chewing
Event|Event|SIMPLE_SEGMENT|10879,10885|false|false|false|||normal
Event|Event|SIMPLE_SEGMENT|10896,10903|false|false|false|||surgery
Finding|Finding|SIMPLE_SEGMENT|10896,10903|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|10896,10903|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|10896,10903|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10896,10903|false|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Event|SIMPLE_SEGMENT|10913,10920|false|false|false|||improve
Finding|Finding|SIMPLE_SEGMENT|10926,10930|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|10926,10930|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|10926,10930|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Drug|Food|SIMPLE_SEGMENT|10939,10944|false|false|false|C0016452|Food|foods
Event|Event|SIMPLE_SEGMENT|10939,10944|false|false|false|||foods
Finding|Finding|SIMPLE_SEGMENT|10972,10976|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|10972,10976|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|10972,10976|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|SIMPLE_SEGMENT|10995,11000|false|false|false|||tired
Finding|Finding|SIMPLE_SEGMENT|10995,11000|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Finding|Intellectual Product|SIMPLE_SEGMENT|10995,11000|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Finding|Sign or Symptom|SIMPLE_SEGMENT|10995,11000|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Event|Event|SIMPLE_SEGMENT|11004,11016|false|false|false|||restlessness
Finding|Finding|SIMPLE_SEGMENT|11004,11016|false|false|false|C0085631;C3887611;C3887612|Agitation;Psychomotor Agitation;Restlessness|restlessness
Finding|Sign or Symptom|SIMPLE_SEGMENT|11004,11016|false|false|false|C0085631;C3887611;C3887612|Agitation;Psychomotor Agitation;Restlessness|restlessness
Event|Event|SIMPLE_SEGMENT|11025,11031|false|false|false|||common
Finding|Functional Concept|SIMPLE_SEGMENT|11025,11031|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Finding|Intellectual Product|SIMPLE_SEGMENT|11025,11031|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Event|Event|SIMPLE_SEGMENT|11036,11048|false|false|false|||Constipation
Finding|Sign or Symptom|SIMPLE_SEGMENT|11036,11048|false|false|false|C0009806|Constipation|Constipation
Event|Event|SIMPLE_SEGMENT|11052,11058|false|false|false|||common
Finding|Functional Concept|SIMPLE_SEGMENT|11052,11058|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Finding|Intellectual Product|SIMPLE_SEGMENT|11052,11058|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Event|Event|SIMPLE_SEGMENT|11063,11067|false|false|false|||sure
Finding|Intellectual Product|SIMPLE_SEGMENT|11063,11067|false|false|false|C4724437|SURE Test|sure
Drug|Food|SIMPLE_SEGMENT|11071,11076|false|false|false|C0452428|Drink (dietary substance)|drink
Event|Event|SIMPLE_SEGMENT|11071,11076|false|false|false|||drink
Event|Event|SIMPLE_SEGMENT|11077,11083|false|false|false|||plenty
Drug|Substance|SIMPLE_SEGMENT|11087,11093|false|false|false|C0302908|Liquid substance|fluids
Event|Event|SIMPLE_SEGMENT|11087,11093|false|false|false|||fluids
Finding|Body Substance|SIMPLE_SEGMENT|11087,11093|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11087,11093|false|false|false|C0016286|Fluid Therapy|fluids
Finding|Finding|SIMPLE_SEGMENT|11105,11109|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|SIMPLE_SEGMENT|11105,11109|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|SIMPLE_SEGMENT|11105,11109|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11105,11120|false|false|false|C0301568|High residue diet|high-fiber diet
Anatomy|Tissue|SIMPLE_SEGMENT|11110,11115|false|false|false|C1304649|Tissue fiber|fiber
Drug|Organic Chemical|SIMPLE_SEGMENT|11110,11115|false|false|false|C0225326;C1321801|Fiber brand of calcium polycarbophil;fiber|fiber
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11110,11115|false|false|false|C0225326;C1321801|Fiber brand of calcium polycarbophil;fiber|fiber
Drug|Food|SIMPLE_SEGMENT|11116,11120|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|SIMPLE_SEGMENT|11116,11120|false|false|false|||diet
Finding|Functional Concept|SIMPLE_SEGMENT|11116,11120|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|SIMPLE_SEGMENT|11116,11120|false|false|false|C0012159|Diet therapy|diet
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|11140,11149|false|false|false|C0027415|Narcotics|narcotics
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11140,11149|false|false|false|C0027415|Narcotics|narcotics
Event|Event|SIMPLE_SEGMENT|11140,11149|false|false|false|||narcotics
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11151,11163|false|false|false|C5886759|Prescription (attribute)|prescription
Event|Event|SIMPLE_SEGMENT|11151,11163|false|false|false|||prescription
Finding|Intellectual Product|SIMPLE_SEGMENT|11151,11163|false|false|false|C1521941|prescription document|prescription
Procedure|Health Care Activity|SIMPLE_SEGMENT|11151,11163|false|false|false|C0033080|Prescription (procedure)|prescription
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11165,11169|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|11165,11169|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|11165,11169|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11170,11181|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11170,11181|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|11170,11181|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|11170,11181|false|false|false|C4284232|Medications|medications
Event|Event|SIMPLE_SEGMENT|11184,11187|false|false|false|||try
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11191,11207|false|false|false|C0013231|Drugs, Non-Prescription|over-the-counter
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|11200,11207|false|false|false|C0702263|Counter brand of Terbufos|counter
Drug|Organic Chemical|SIMPLE_SEGMENT|11200,11207|false|false|false|C0702263|Counter brand of Terbufos|counter
Event|Event|SIMPLE_SEGMENT|11208,11213|false|false|false|||stool
Finding|Body Substance|SIMPLE_SEGMENT|11208,11213|false|false|false|C0015733|Feces|stool
Drug|Organic Chemical|SIMPLE_SEGMENT|11208,11222|false|false|false|C0301470;C1154263|Stool Softener;Stool Softener brand of docusate sodium|stool softener
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11208,11222|false|false|false|C0301470;C1154263|Stool Softener;Stool Softener brand of docusate sodium|stool softener
Event|Event|SIMPLE_SEGMENT|11214,11222|false|false|false|||softener
Event|Event|SIMPLE_SEGMENT|11233,11237|false|false|false|||Call
Event|Event|SIMPLE_SEGMENT|11243,11249|false|false|false|||Doctor
Finding|Intellectual Product|SIMPLE_SEGMENT|11243,11249|false|false|false|C2348314|Doctor - Title|Doctor
Finding|Finding|SIMPLE_SEGMENT|11265,11271|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Finding|Intellectual Product|SIMPLE_SEGMENT|11265,11271|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Finding|Finding|SIMPLE_SEGMENT|11265,11276|false|false|false|C0278140;C4050465;C4521229|Neck Pain Score 6;Severe Extremity Pain;Severe pain|Severe pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11272,11276|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|11272,11276|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|11272,11276|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|11272,11276|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|11278,11286|false|false|false|||swelling
Finding|Finding|SIMPLE_SEGMENT|11278,11286|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|11278,11286|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11288,11295|false|false|false|C0041834|Erythema|redness
Event|Event|SIMPLE_SEGMENT|11288,11295|false|false|false|||redness
Finding|Finding|SIMPLE_SEGMENT|11288,11295|false|false|false|C0332575|Redness|redness
Event|Event|SIMPLE_SEGMENT|11299,11307|false|false|false|||drainage
Finding|Body Substance|SIMPLE_SEGMENT|11299,11307|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|SIMPLE_SEGMENT|11299,11307|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11299,11307|false|false|false|C0013103|Drainage procedure|drainage
Anatomy|Body Location or Region|SIMPLE_SEGMENT|11317,11325|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|11317,11325|false|false|false|C0332803|Surgical wound|incision
Event|Event|SIMPLE_SEGMENT|11317,11325|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11317,11325|false|false|false|C0184898|Surgical incisions|incision
Anatomy|Body Location or Region|SIMPLE_SEGMENT|11327,11331|false|false|false|C1515974|Anatomic Site|site
Finding|Intellectual Product|SIMPLE_SEGMENT|11327,11331|false|false|false|C1546778||site
Finding|Finding|SIMPLE_SEGMENT|11337,11342|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|11337,11342|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Finding|Intellectual Product|SIMPLE_SEGMENT|11362,11369|false|false|false|C0542560|Academic degree|degrees
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11384,11390|false|false|false|C4255480||Nausea
Event|Event|SIMPLE_SEGMENT|11384,11390|false|false|false|||Nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|11384,11390|false|false|false|C0027497|Nausea|Nausea
Event|Event|SIMPLE_SEGMENT|11398,11406|false|false|false|||vomiting
Finding|Sign or Symptom|SIMPLE_SEGMENT|11398,11406|false|false|false|C0042963|Vomiting|vomiting
Finding|Finding|SIMPLE_SEGMENT|11410,11417|false|false|false|C4085555|Extreme Response|Extreme
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|11418,11428|false|false|false|C2830004|Somnolence|sleepiness
Event|Event|SIMPLE_SEGMENT|11418,11428|false|false|false|||sleepiness
Finding|Finding|SIMPLE_SEGMENT|11418,11428|false|false|false|C0013144|Drowsiness|sleepiness
Event|Event|SIMPLE_SEGMENT|11443,11447|false|false|false|||able
Finding|Finding|SIMPLE_SEGMENT|11443,11447|false|true|false|C1299581|Able (qualifier value)|able
Event|Event|SIMPLE_SEGMENT|11451,11455|false|false|false|||stay
Drug|Organic Chemical|SIMPLE_SEGMENT|11451,11461|false|false|false|C0723446|Stay Awake|stay awake
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11451,11461|false|false|false|C0723446|Stay Awake|stay awake
Event|Event|SIMPLE_SEGMENT|11456,11461|false|false|false|||awake
Finding|Finding|SIMPLE_SEGMENT|11456,11461|false|false|false|C0234422|Awake (finding)|awake
Finding|Finding|SIMPLE_SEGMENT|11465,11471|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Finding|Intellectual Product|SIMPLE_SEGMENT|11465,11471|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Event|Event|SIMPLE_SEGMENT|11472,11481|false|false|false|||headaches
Finding|Sign or Symptom|SIMPLE_SEGMENT|11472,11481|false|false|false|C0018681|Headache|headaches
Event|Event|SIMPLE_SEGMENT|11486,11494|false|false|false|||relieved
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11498,11502|false|true|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|11498,11502|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|11498,11502|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|11498,11512|false|false|false|C0002771;C0722425|Analgesics;Pain Relieve brand of acetaminophen|pain relievers
Drug|Organic Chemical|SIMPLE_SEGMENT|11498,11512|false|false|false|C0002771;C0722425|Analgesics;Pain Relieve brand of acetaminophen|pain relievers
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11498,11512|false|false|false|C0002771;C0722425|Analgesics;Pain Relieve brand of acetaminophen|pain relievers
Event|Event|SIMPLE_SEGMENT|11503,11512|false|false|false|||relievers
Event|Event|SIMPLE_SEGMENT|11516,11524|false|false|false|||Seizures
Finding|Sign or Symptom|SIMPLE_SEGMENT|11516,11524|false|false|false|C0036572|Seizures|Seizures
Finding|Finding|SIMPLE_SEGMENT|11532,11535|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|11532,11535|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Event|Event|SIMPLE_SEGMENT|11536,11544|false|false|false|||problems
Finding|Idea or Concept|SIMPLE_SEGMENT|11536,11544|false|false|false|C1546466|Problems - What subject filter|problems
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11555,11561|false|false|false|C2707266||vision
Event|Event|SIMPLE_SEGMENT|11555,11561|false|false|false|||vision
Finding|Organism Function|SIMPLE_SEGMENT|11555,11561|false|false|false|C0042789|Vision|vision
Event|Event|SIMPLE_SEGMENT|11565,11572|false|false|false|||ability
Finding|Functional Concept|SIMPLE_SEGMENT|11565,11572|false|false|false|C5891046|Oral Intake Ability|ability
Finding|Intellectual Product|SIMPLE_SEGMENT|11565,11575|false|false|false|C5420000|Ability Question|ability to
Finding|Finding|SIMPLE_SEGMENT|11565,11581|false|false|false|C0564214|Ability to speak|ability to speak
Event|Event|SIMPLE_SEGMENT|11576,11581|false|false|false|||speak
Finding|Finding|SIMPLE_SEGMENT|11576,11581|false|false|false|C0234856;C0600116;C1547187|Does speak;Speak - language ability;Speaking (function)|speak
Finding|Idea or Concept|SIMPLE_SEGMENT|11576,11581|false|false|false|C0234856;C0600116;C1547187|Does speak;Speak - language ability;Speaking (function)|speak
Finding|Individual Behavior|SIMPLE_SEGMENT|11576,11581|false|false|false|C0234856;C0600116;C1547187|Does speak;Speak - language ability;Speaking (function)|speak
Event|Event|SIMPLE_SEGMENT|11585,11593|false|false|false|||Weakness
Finding|Sign or Symptom|SIMPLE_SEGMENT|11585,11593|false|false|false|C0004093;C3714552|Asthenia;Weakness|Weakness
Event|Event|SIMPLE_SEGMENT|11597,11604|false|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|11597,11604|false|false|false|C0392747|Changing|changes
Event|Event|SIMPLE_SEGMENT|11608,11617|false|false|false|||sensation
Finding|Finding|SIMPLE_SEGMENT|11608,11617|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|11608,11617|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|SIMPLE_SEGMENT|11608,11617|false|false|false|C2229507|sensory exam|sensation
Anatomy|Body Location or Region|SIMPLE_SEGMENT|11626,11630|false|false|false|C0015450;C4266571|Face;Head>Face|face
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11626,11630|false|false|false|C3160739|FANCONI ANEMIA, COMPLEMENTATION GROUP E|face
Finding|Gene or Genome|SIMPLE_SEGMENT|11626,11630|false|false|false|C1414531;C1423759;C2828055|ELOVL6 gene;FANCE gene;FANCE wt Allele|face
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11632,11636|false|false|false|C0446516|Upper arm|arms
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11632,11636|false|false|false|C5782111||arms
Disorder|Neoplastic Process|SIMPLE_SEGMENT|11632,11636|false|false|false|C0206655|Alveolar rhabdomyosarcoma|arms
Event|Event|SIMPLE_SEGMENT|11632,11636|false|false|false|||arms
Finding|Gene or Genome|SIMPLE_SEGMENT|11632,11636|false|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Finding|Intellectual Product|SIMPLE_SEGMENT|11632,11636|false|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11641,11644|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Functional Concept|SIMPLE_SEGMENT|11646,11650|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|Call
Finding|Gene or Genome|SIMPLE_SEGMENT|11646,11650|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|Call
Finding|Intellectual Product|SIMPLE_SEGMENT|11646,11650|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|Call
Finding|Mental Process|SIMPLE_SEGMENT|11646,11650|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|Call
Finding|Finding|SIMPLE_SEGMENT|11677,11686|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Idea or Concept|SIMPLE_SEGMENT|11677,11686|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Intellectual Product|SIMPLE_SEGMENT|11677,11686|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Pathologic Function|SIMPLE_SEGMENT|11677,11686|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|11677,11686|false|false|false|C0013956|Emergency Situation|Emergency
Procedure|Health Care Activity|SIMPLE_SEGMENT|11677,11686|false|false|false|C1553500|emergency encounter|Emergency
Finding|Idea or Concept|SIMPLE_SEGMENT|11677,11691|false|false|false|C1546435|Encounter Referral Source - emergency room|Emergency Room
Finding|Mental Process|SIMPLE_SEGMENT|11699,11709|false|false|false|C0237607;C0596545|Experience;Experience (Practice)|experience
Event|Event|SIMPLE_SEGMENT|11743,11751|false|false|false|||numbness
Finding|Finding|SIMPLE_SEGMENT|11743,11751|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|SIMPLE_SEGMENT|11743,11751|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Event|Event|SIMPLE_SEGMENT|11755,11763|false|false|false|||weakness
Finding|Sign or Symptom|SIMPLE_SEGMENT|11755,11763|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Anatomy|Body Location or Region|SIMPLE_SEGMENT|11771,11775|false|false|false|C0015450;C4266571|Face;Head>Face|face
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11771,11775|false|false|false|C3160739|FANCONI ANEMIA, COMPLEMENTATION GROUP E|face
Finding|Gene or Genome|SIMPLE_SEGMENT|11771,11775|false|false|false|C1414531;C1423759;C2828055|ELOVL6 gene;FANCE gene;FANCE wt Allele|face
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11777,11780|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|11777,11780|false|false|false|C3495676|Anorectal Malformations|arm
Event|Event|SIMPLE_SEGMENT|11777,11780|false|false|false|||arm
Finding|Gene or Genome|SIMPLE_SEGMENT|11777,11780|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|11777,11780|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|SIMPLE_SEGMENT|11777,11780|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11777,11780|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11785,11788|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|11799,11808|false|false|false|C0009676|Confusion|confusion
Event|Event|SIMPLE_SEGMENT|11799,11808|false|false|false|||confusion
Finding|Finding|SIMPLE_SEGMENT|11799,11808|false|false|false|C0683369|Clouded consciousness|confusion
Event|Event|SIMPLE_SEGMENT|11812,11819|false|false|false|||trouble
Event|Event|SIMPLE_SEGMENT|11820,11828|false|false|false|||speaking
Event|Event|SIMPLE_SEGMENT|11832,11845|false|false|false|||understanding
Finding|Mental Process|SIMPLE_SEGMENT|11832,11845|false|false|false|C0162340|Comprehension|understanding
Event|Event|SIMPLE_SEGMENT|11864,11871|false|false|false|||walking
Event|Event|SIMPLE_SEGMENT|11873,11882|false|false|false|||dizziness
Finding|Sign or Symptom|SIMPLE_SEGMENT|11873,11882|false|false|false|C0012833;C0042571|Dizziness;Vertigo|dizziness
Event|Event|SIMPLE_SEGMENT|11887,11891|false|false|false|||loss
Finding|Finding|SIMPLE_SEGMENT|11887,11891|false|false|false|C5890125|Loss (adaptation)|loss
Finding|Finding|SIMPLE_SEGMENT|11887,11902|false|false|false|C0241981|Impairment of balance|loss of balance
Drug|Organic Chemical|SIMPLE_SEGMENT|11895,11902|false|false|false|C4319618|Balance (substance)|balance
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11895,11902|false|false|false|C4319618|Balance (substance)|balance
Event|Event|SIMPLE_SEGMENT|11895,11902|false|false|false|||balance
Finding|Finding|SIMPLE_SEGMENT|11895,11902|false|false|false|C0014653;C0560184|Ability to balance;Equilibrium|balance
Finding|Organism Function|SIMPLE_SEGMENT|11895,11902|false|false|false|C0014653;C0560184|Ability to balance;Equilibrium|balance
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|11895,11902|false|false|false|C2174421|examination of balance|balance
Event|Event|SIMPLE_SEGMENT|11907,11919|false|false|false|||coordination
Finding|Functional Concept|SIMPLE_SEGMENT|11907,11919|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|coordination
Finding|Idea or Concept|SIMPLE_SEGMENT|11907,11919|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|coordination
Finding|Physiologic Function|SIMPLE_SEGMENT|11907,11919|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|coordination
Finding|Finding|SIMPLE_SEGMENT|11930,11936|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|11930,11936|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Event|Event|SIMPLE_SEGMENT|11937,11946|false|false|false|||headaches
Finding|Sign or Symptom|SIMPLE_SEGMENT|11937,11946|false|false|false|C0018681|Headache|headaches
Event|Event|SIMPLE_SEGMENT|11961,11967|false|false|false|||reason
Finding|Idea or Concept|SIMPLE_SEGMENT|11961,11967|true|false|false|C0392360|Indication of (contextual qualifier)|reason
Procedure|Health Care Activity|SIMPLE_SEGMENT|11971,11979|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11980,11992|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|11980,11992|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|11980,11992|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

