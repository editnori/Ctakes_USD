 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|44,53|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|44,53|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|44,58|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|78,87|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|78,87|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|78,87|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|78,87|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|78,87|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|78,92|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|110,115|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|110,115|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|110,115|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|134,137|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|134,137|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|134,137|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|134,137|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|134,137|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|145,152|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|145,152|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|154,162|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|165,174|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|165,174|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|165,174|false|false|false|C0020517|Hypersensitivity|Allergies
Attribute|Clinical Attribute|SIMPLE_SEGMENT|186,195|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|186,195|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|186,195|false|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|198,220|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|206,210|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|SIMPLE_SEGMENT|206,210|false|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|SIMPLE_SEGMENT|206,220|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Event|Event|SIMPLE_SEGMENT|211,220|false|false|false|||Reactions
Event|Event|SIMPLE_SEGMENT|223,232|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|223,232|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|241,256|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|247,256|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|247,256|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|247,256|false|false|false|C5441521|Complaint (finding)|Complaint
Anatomy|Body Location or Region|SIMPLE_SEGMENT|258,263|false|false|false|C1548802|Body Site Modifier - Lower|Lower
Event|Activity|SIMPLE_SEGMENT|258,263|false|false|false|C2003888|Lower (action)|Lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|258,273|false|false|false|C0023216|Lower Extremity|Lower extremity
Finding|Pathologic Function|SIMPLE_SEGMENT|258,282|false|false|false|C0581394|Swelling of lower limb|Lower extremity swelling
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|264,273|false|false|false|C0015385|Limb structure|extremity
Finding|Sign or Symptom|SIMPLE_SEGMENT|264,282|false|false|false|C0158369|Swelling of limb|extremity swelling
Event|Event|SIMPLE_SEGMENT|274,282|false|false|false|||swelling
Finding|Finding|SIMPLE_SEGMENT|274,282|false|true|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|274,282|false|true|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Classification|SIMPLE_SEGMENT|285,290|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|291,299|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|291,299|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|303,321|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|312,321|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|312,321|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|312,321|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|312,321|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|312,321|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|SIMPLE_SEGMENT|330,337|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|330,337|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|330,337|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|330,337|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|330,340|false|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|330,356|false|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|330,356|false|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|341,348|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|341,348|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|341,356|false|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|349,356|false|false|false|C0221423|Illness (finding)|Illness
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|370,381|false|false|false|C0851145|on warfarin|on warfarin
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|373,381|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|SIMPLE_SEGMENT|373,381|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|373,381|false|false|false|C0043031|warfarin|warfarin
Event|Event|SIMPLE_SEGMENT|373,381|false|false|false|||warfarin
Drug|Organic Chemical|SIMPLE_SEGMENT|398,405|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|398,405|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Attribute|Clinical Attribute|SIMPLE_SEGMENT|406,411|false|false|false|C0232117|Pulse Rate|pulse
Event|Event|SIMPLE_SEGMENT|406,411|false|false|false|||pulse
Finding|Physiologic Function|SIMPLE_SEGMENT|406,411|false|false|false|C0391850|Physiologic pulse|pulse
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|406,411|false|false|false|C1947910|Pulse phenomenon|pulse
Procedure|Health Care Activity|SIMPLE_SEGMENT|406,411|false|false|false|C0034107|Pulse taking|pulse
Event|Event|SIMPLE_SEGMENT|429,436|false|false|false|||swollen
Finding|Finding|SIMPLE_SEGMENT|429,436|false|false|false|C0038999|Swelling|swollen
Finding|Sign or Symptom|SIMPLE_SEGMENT|441,448|false|false|false|C0030193|Pain|painful
Anatomy|Body Location or Region|SIMPLE_SEGMENT|449,455|false|false|false|C0003086|Ankle|ankles
Event|Event|SIMPLE_SEGMENT|467,477|false|false|false|||complaints
Finding|Finding|SIMPLE_SEGMENT|467,477|true|false|false|C5441521|Complaint (finding)|complaints
Event|Event|SIMPLE_SEGMENT|507,516|false|false|false|||concerned
Event|Event|SIMPLE_SEGMENT|538,546|false|false|false|||swelling
Finding|Finding|SIMPLE_SEGMENT|538,546|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|538,546|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Event|Event|SIMPLE_SEGMENT|556,565|false|false|false|||inability
Finding|Finding|SIMPLE_SEGMENT|556,573|false|false|false|C0560046|Unable to walk (finding)|inability to walk
Event|Event|SIMPLE_SEGMENT|569,573|false|false|false|||walk
Attribute|Clinical Attribute|SIMPLE_SEGMENT|582,586|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|582,586|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|582,586|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|582,586|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|SIMPLE_SEGMENT|595,601|false|false|false|C1561668|History of fall|a fall
Event|Event|SIMPLE_SEGMENT|597,601|false|false|false|||fall
Finding|Finding|SIMPLE_SEGMENT|597,601|false|false|false|C0085639|Falls|fall
Finding|Intellectual Product|SIMPLE_SEGMENT|622,626|false|false|false|C1561540|Transaction counts and value totals - week|week
Finding|Gene or Genome|SIMPLE_SEGMENT|627,630|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|SIMPLE_SEGMENT|632,639|false|false|false|||reports
Anatomy|Body Location or Region|SIMPLE_SEGMENT|643,647|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|643,647|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|643,647|true|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|643,647|true|false|false|C0876917|Procedure on head|head
Event|Event|SIMPLE_SEGMENT|648,654|false|false|false|||strike
Event|Occupational Activity|SIMPLE_SEGMENT|648,654|true|false|false|C0038452|Strikes, Employee|strike
Finding|Finding|SIMPLE_SEGMENT|689,693|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|689,693|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|689,693|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|710,715|false|false|false|C1550012|Local Remote Control State - Local|local
Event|Event|SIMPLE_SEGMENT|733,738|false|false|false|||found
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|749,758|false|false|false|C0549207|Bone structure of spine|vertebral
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|749,767|false|false|false|C0080179|Spinal Fractures|vertebral fracture
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|759,767|false|false|false|C0016658|Fracture|fracture
Event|Event|SIMPLE_SEGMENT|759,767|false|false|false|||fracture
Event|Event|SIMPLE_SEGMENT|790,795|false|false|false|||brace
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|790,795|false|false|false|C1828220|Application of brace (procedure)|brace
Event|Event|SIMPLE_SEGMENT|815,822|false|false|false|||wearing
Event|Event|SIMPLE_SEGMENT|853,857|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|853,857|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|853,857|false|false|false|C0582103|Medical Examination|exam
Event|Event|SIMPLE_SEGMENT|862,872|false|false|false|||remarkable
Finding|Finding|SIMPLE_SEGMENT|877,901|false|false|false|C2109101|swelling of both ankles|bilateral ankle swelling
Anatomy|Body Location or Region|SIMPLE_SEGMENT|887,892|false|false|false|C0003086;C0003087;C4284979|Ankle;Ankle joint structure;Lower extremity>Ankle|ankle
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|887,892|false|false|false|C0003086;C0003087;C4284979|Ankle;Ankle joint structure;Lower extremity>Ankle|ankle
Finding|Pathologic Function|SIMPLE_SEGMENT|887,901|false|false|false|C0235439|Ankle edema (finding)|ankle swelling
Event|Event|SIMPLE_SEGMENT|893,901|false|false|false|||swelling
Finding|Finding|SIMPLE_SEGMENT|893,901|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|893,901|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Finding|SIMPLE_SEGMENT|908,924|false|false|false|C1720001|3+ pitting edema|3+ pitting edema
Finding|Functional Concept|SIMPLE_SEGMENT|911,918|false|false|false|C0205323|Pitting|pitting
Finding|Finding|SIMPLE_SEGMENT|911,924|false|false|false|C0333243|Pitting edema|pitting edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|919,924|false|false|false|C1717255||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|919,924|false|false|false|C0013604|Edema|edema
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|926,930|false|false|false|C0009443;C0024117|Chronic Obstructive Airway Disease;Common Cold|cold
Drug|Organic Chemical|SIMPLE_SEGMENT|926,930|false|false|false|C0719425|Cold brand of chlorpheniramine-phenylpropanolamine|cold
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|926,930|false|false|false|C0719425|Cold brand of chlorpheniramine-phenylpropanolamine|cold
Event|Event|SIMPLE_SEGMENT|926,930|false|false|false|||cold
Finding|Organism Function|SIMPLE_SEGMENT|926,930|false|false|false|C0234192|Cold Sensation|cold
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|926,930|false|false|false|C0009264|Cold Temperature|cold
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|926,930|false|false|false|C0010412|Cold Therapy|cold
Finding|Finding|SIMPLE_SEGMENT|935,942|false|false|false|C0302133|Mottling|mottled
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|943,947|false|false|false|C0040357;C4299090|Lower extremity>Toes;Toes|toes
Drug|Food|SIMPLE_SEGMENT|979,985|false|false|false|C5890763||pulses
Event|Event|SIMPLE_SEGMENT|979,985|false|false|false|||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|979,985|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|979,985|false|false|false|C0034107|Pulse taking|pulses
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|994,1014|true|false|false|C0152027|Sensory Disorders|sensory disturbances
Event|Event|SIMPLE_SEGMENT|1002,1014|false|false|false|||disturbances
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1016,1019|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Hormone|SIMPLE_SEGMENT|1016,1019|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1016,1019|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Event|Event|SIMPLE_SEGMENT|1016,1019|false|false|false|||BNP
Finding|Gene or Genome|SIMPLE_SEGMENT|1016,1019|false|false|false|C1417808;C2982014|NPPB gene;NPPB wt Allele|BNP
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1016,1019|false|false|false|C1095989|Brain natriuretic peptide measurement|BNP
Event|Event|SIMPLE_SEGMENT|1024,1032|false|false|false|||elevated
Event|Event|SIMPLE_SEGMENT|1043,1046|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1043,1046|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|SIMPLE_SEGMENT|1047,1053|false|false|false|||showed
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1054,1063|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1054,1063|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|1054,1063|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|1054,1069|false|false|false|C0034063|Pulmonary Edema|pulmonary edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1064,1069|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|1064,1069|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|1064,1069|false|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|1071,1076|false|false|false|||LENIs
Event|Event|SIMPLE_SEGMENT|1082,1090|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|1082,1090|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|1082,1090|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1082,1090|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|SIMPLE_SEGMENT|1082,1094|false|false|false|C0205160|Negative|negative for
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1095,1098|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1095,1098|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1095,1098|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|SIMPLE_SEGMENT|1095,1098|false|false|false|||DVT
Event|Event|SIMPLE_SEGMENT|1115,1121|false|false|false|||showed
Event|Event|SIMPLE_SEGMENT|1125,1133|false|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|1125,1133|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|1125,1136|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1137,1148|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1137,1148|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1137,1157|true|false|false|C0031039|Pericardial effusion|pericardial effusion
Finding|Body Substance|SIMPLE_SEGMENT|1137,1157|true|false|false|C1253937|Pericardial effusion body substance|pericardial effusion
Event|Event|SIMPLE_SEGMENT|1149,1157|false|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|1149,1157|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|1149,1157|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|1149,1157|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1161,1164|false|false|false|C3498924|lamina IVC|IVC
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1161,1164|true|false|false|C4085887|Inspiratory Vital Capacity Test|IVC
Finding|Intellectual Product|SIMPLE_SEGMENT|1166,1172|false|false|false|C1705102|Volume (publication)|volume
Finding|Finding|SIMPLE_SEGMENT|1166,1182|false|false|false|C0546884|Hypovolemia|volume depletion
Event|Event|SIMPLE_SEGMENT|1173,1182|false|false|false|||depletion
Finding|Functional Concept|SIMPLE_SEGMENT|1173,1182|false|false|false|C0333668|Depletion|depletion
Drug|Organic Chemical|SIMPLE_SEGMENT|1207,1212|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1207,1212|false|false|false|C0699992|Lasix|Lasix
Event|Event|SIMPLE_SEGMENT|1207,1212|false|false|false|||Lasix
Event|Event|SIMPLE_SEGMENT|1214,1221|false|false|false|||Nursing
Finding|Organism Function|SIMPLE_SEGMENT|1214,1221|false|false|false|C0006147|Breast Feeding|Nursing
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1214,1221|false|false|false|C0028678|RNAx nursing therapy actions|Nursing
Event|Event|SIMPLE_SEGMENT|1232,1237|false|false|false|||noted
Event|Event|SIMPLE_SEGMENT|1246,1250|false|false|false|||able
Finding|Finding|SIMPLE_SEGMENT|1246,1250|false|false|false|C1299581|Able (qualifier value)|able
Event|Event|SIMPLE_SEGMENT|1255,1260|false|false|false|||stand
Finding|Finding|SIMPLE_SEGMENT|1255,1260|false|false|false|C0038137;C0596013|Does stand;standards characteristics|stand
Finding|Functional Concept|SIMPLE_SEGMENT|1255,1260|false|false|false|C0038137;C0596013|Does stand;standards characteristics|stand
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1265,1271|false|false|false|C0944911||weight
Event|Event|SIMPLE_SEGMENT|1265,1271|false|false|false|||weight
Finding|Finding|SIMPLE_SEGMENT|1265,1271|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|1265,1271|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|1265,1271|false|false|false|C1305866|Weighing patient|weight
Finding|Finding|SIMPLE_SEGMENT|1291,1295|false|false|false|C0085639|Falls|fall
Finding|Finding|SIMPLE_SEGMENT|1291,1300|false|false|false|C1268740|At increased risk for falls|fall risk
Event|Event|SIMPLE_SEGMENT|1296,1300|false|false|false|||risk
Finding|Idea or Concept|SIMPLE_SEGMENT|1296,1300|false|false|false|C0035647|Risk|risk
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1304,1309|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|spine
Anatomy|Cell Component|SIMPLE_SEGMENT|1304,1309|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|spine
Finding|Finding|SIMPLE_SEGMENT|1304,1309|false|false|false|C0150920|Spine Problem|spine
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1310,1314|false|false|false|C1561572;C1704608|Film Dosage Form;film - layer|film
Drug|Substance|SIMPLE_SEGMENT|1310,1314|false|false|false|C1561572;C1704608|Film Dosage Form;film - layer|film
Event|Event|SIMPLE_SEGMENT|1310,1314|false|false|false|||film
Finding|Intellectual Product|SIMPLE_SEGMENT|1310,1314|false|false|false|C4019020||film
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|1356,1365|true|false|false|C0016658|Fracture|fractures
Event|Event|SIMPLE_SEGMENT|1356,1365|false|false|false|||fractures
Finding|Finding|SIMPLE_SEGMENT|1356,1365|true|false|false|C4554413|Fractured|fractures
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|1370,1382|false|false|false|C0012691|Dislocations|dislocations
Event|Event|SIMPLE_SEGMENT|1370,1382|false|false|false|||dislocations
Event|Event|SIMPLE_SEGMENT|1390,1399|false|false|false|||triggered
Event|Event|SIMPLE_SEGMENT|1404,1415|false|false|false|||hypotension
Finding|Finding|SIMPLE_SEGMENT|1404,1415|false|false|false|C0020649|Hypotension|hypotension
Event|Event|SIMPLE_SEGMENT|1431,1442|false|false|false|||bradycardia
Finding|Finding|SIMPLE_SEGMENT|1431,1442|false|false|false|C0428977;C3812171|Bradycardia;Bradycardia by ECG Finding|bradycardia
Event|Event|SIMPLE_SEGMENT|1460,1469|false|false|false|||responded
Finding|Finding|SIMPLE_SEGMENT|1470,1474|false|false|false|C5575035|Well (answer to question)|well
Drug|Substance|SIMPLE_SEGMENT|1484,1489|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|1484,1489|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|1490,1497|false|false|false|||boluses
Event|Event|SIMPLE_SEGMENT|1516,1524|false|false|false|||transfer
Finding|Functional Concept|SIMPLE_SEGMENT|1516,1524|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|SIMPLE_SEGMENT|1516,1524|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|SIMPLE_SEGMENT|1516,1524|false|false|false|C4706767|Transfer (immobility management)|transfer
Event|Event|SIMPLE_SEGMENT|1534,1536|false|false|false|||HR
Finding|Finding|SIMPLE_SEGMENT|1578,1598|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|1583,1590|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|1583,1590|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|1583,1590|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|1583,1590|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1583,1590|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|1583,1598|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1591,1598|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1591,1598|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1591,1598|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1600,1605|false|false|false|C0378717|elongation factor DmS-II|DM II
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1607,1610|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|1607,1610|false|false|false|||HTN
Drug|Organic Chemical|SIMPLE_SEGMENT|1636,1644|false|false|false|C0699129|Coumadin|coumadin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1636,1644|false|false|false|C0699129|Coumadin|coumadin
Event|Event|SIMPLE_SEGMENT|1636,1644|false|false|false|||coumadin
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1646,1654|false|false|false|C0033572;C4266527|Prostate;Structure of prostate (body structure)|prostate
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1646,1654|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|prostate
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1646,1654|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|prostate
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1646,1657|false|false|false|C0376358|Malignant neoplasm of prostate|prostate CA
Event|Event|SIMPLE_SEGMENT|1655,1657|false|false|false|||CA
Event|Event|SIMPLE_SEGMENT|1659,1666|false|false|false|||treated
Finding|Functional Concept|SIMPLE_SEGMENT|1686,1692|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|1686,1700|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|1693,1700|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1693,1700|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1693,1700|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1693,1700|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|1706,1712|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|1706,1712|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|1706,1712|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|1706,1712|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|1706,1720|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|1713,1720|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1713,1720|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1713,1720|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1713,1720|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Event|Event|SIMPLE_SEGMENT|1742,1750|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|1742,1750|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|1742,1750|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1742,1750|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|1742,1755|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1742,1755|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|1751,1755|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|1751,1755|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1751,1755|false|false|false|C0582103|Medical Examination|Exam
Event|Event|SIMPLE_SEGMENT|1769,1771|false|false|false|||BP
Finding|Conceptual Entity|SIMPLE_SEGMENT|1776,1780|false|false|false|C1412365;C2945620;C3812647|ALPP gene;ALPP wt Allele;Palp - CHV concept|palp
Finding|Gene or Genome|SIMPLE_SEGMENT|1776,1780|false|false|false|C1412365;C2945620;C3812647|ALPP gene;ALPP wt Allele;Palp - CHV concept|palp
Event|Event|SIMPLE_SEGMENT|1808,1815|false|false|false|||GENERAL
Finding|Classification|SIMPLE_SEGMENT|1808,1815|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|1808,1815|false|false|false|C3812897|General medical service|GENERAL
Finding|Finding|SIMPLE_SEGMENT|1817,1821|false|false|false|C5575035|Well (answer to question)|Well
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1839,1842|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1839,1842|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1839,1842|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|1839,1842|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1839,1842|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|1839,1842|false|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|1839,1842|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Event|Event|SIMPLE_SEGMENT|1844,1855|false|false|false|||comfortable
Finding|Finding|SIMPLE_SEGMENT|1844,1855|false|false|false|C5546696|Feeling comfortable|comfortable
Event|Event|SIMPLE_SEGMENT|1857,1868|false|false|false|||appropriate
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1872,1877|false|false|false|C1512338|HEENT|HEENT
Event|Event|SIMPLE_SEGMENT|1886,1893|false|false|false|||sclerae
Event|Event|SIMPLE_SEGMENT|1894,1903|false|false|false|||anicteric
Finding|Finding|SIMPLE_SEGMENT|1894,1903|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1905,1908|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1905,1908|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1911,1916|false|false|false|C0018787;C4037974|Chest>Heart;Heart|HEART
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1911,1916|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|HEART
Event|Event|SIMPLE_SEGMENT|1911,1916|false|false|false|||HEART
Finding|Sign or Symptom|SIMPLE_SEGMENT|1911,1916|false|false|false|C0795691|HEART PROBLEM|HEART
Event|Event|SIMPLE_SEGMENT|1930,1939|false|false|false|||irregular
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|1948,1956|false|false|false|C0039155|Systole|systolic
Finding|Finding|SIMPLE_SEGMENT|1948,1972|false|false|false|C0694547|SYSTOLIC EJECTION MURMUR|systolic ejection murmur
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1957,1965|false|false|false|C0812388|Ejection time|ejection
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|1957,1965|false|false|false|C0336969|Ejection as a Sports activity|ejection
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|1957,1965|false|false|false|C0302131|Ejection as a Circumstance of Injury|ejection
Finding|Finding|SIMPLE_SEGMENT|1957,1972|false|false|false|C0277910|Ejection Murmurs|ejection murmur
Event|Event|SIMPLE_SEGMENT|1966,1972|false|false|false|||murmur
Finding|Finding|SIMPLE_SEGMENT|1966,1972|false|false|false|C0018808|Heart murmur|murmur
Event|Event|SIMPLE_SEGMENT|1974,1981|false|false|false|||loudest
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|1989,1992|false|false|false|C0262278;C4281534|Lunate Sulcus;lunate sulcus of the macaque|LUS
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2014,2019|false|false|false|C0024109|Lung|LUNGS
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2021,2024|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|SIMPLE_SEGMENT|2021,2024|false|false|false|||CTA
Finding|Gene or Genome|SIMPLE_SEGMENT|2021,2024|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2021,2024|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Finding|Idea or Concept|SIMPLE_SEGMENT|2044,2048|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Drug|Inorganic Chemical|SIMPLE_SEGMENT|2049,2052|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2049,2052|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|SIMPLE_SEGMENT|2049,2052|false|false|false|C0001861;C3536832|Air (substance);air|air
Finding|Finding|SIMPLE_SEGMENT|2049,2052|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|SIMPLE_SEGMENT|2049,2052|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|SIMPLE_SEGMENT|2049,2052|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2049,2061|false|false|false|C0001868|Air Movements|air movement
Event|Event|SIMPLE_SEGMENT|2053,2061|false|false|false|||movement
Finding|Organism Function|SIMPLE_SEGMENT|2053,2061|false|false|false|C0026649|Movement|movement
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2063,2067|false|false|true|C0231832|Respiratory rate|resp
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2063,2067|false|false|true|C0851355|Respiratory, thoracic and mediastinal disorders|resp
Event|Event|SIMPLE_SEGMENT|2068,2077|false|false|false|||unlabored
Finding|Functional Concept|SIMPLE_SEGMENT|2068,2077|false|false|false|C2983702|Unlabored|unlabored
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2082,2089|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2082,2089|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|SIMPLE_SEGMENT|2082,2089|false|false|false|||ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|2082,2089|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2107,2111|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|SIMPLE_SEGMENT|2107,2111|false|false|false|||soft
Event|Event|SIMPLE_SEGMENT|2122,2128|false|false|false|||masses
Event|Event|SIMPLE_SEGMENT|2132,2135|false|false|false|||HSM
Finding|Gene or Genome|SIMPLE_SEGMENT|2132,2135|true|false|false|C1537594|LRRC4B gene|HSM
Event|Event|SIMPLE_SEGMENT|2141,2148|false|false|false|||rebound
Event|Event|SIMPLE_SEGMENT|2149,2157|false|false|false|||guarding
Finding|Finding|SIMPLE_SEGMENT|2149,2157|false|false|false|C0427198|Protective muscle spasm|guarding
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2161,2172|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|2174,2182|false|false|false|C0009938|Contusions|Bruising
Event|Event|SIMPLE_SEGMENT|2174,2182|false|false|false|||Bruising
Finding|Finding|SIMPLE_SEGMENT|2174,2182|false|false|false|C2136686|reported bruising (history)|Bruising
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2190,2194|false|false|false|C0040357;C4299090|Lower extremity>Toes;Toes|toes
Finding|Functional Concept|SIMPLE_SEGMENT|2202,2206|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2202,2211|false|false|false|C0230461|Structure of left foot|left foot
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2207,2211|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|2207,2211|false|false|false|C0555980|Foot problem|foot
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2217,2222|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|2217,2222|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|2217,2222|false|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|2230,2240|false|false|false|||pronounced
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2248,2252|false|false|false|C0016504|Foot|feet
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2253,2259|false|false|false|C0003086|Ankle|ankles
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2271,2277|false|false|false|C0039866|Thigh structure|thighs
Event|Event|SIMPLE_SEGMENT|2288,2293|false|false|false|||Awake
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2295,2300|false|false|false|C5890168||alert
Drug|Organic Chemical|SIMPLE_SEGMENT|2295,2300|false|false|false|C0718338|Alert brand of caffeine|alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2295,2300|false|false|false|C0718338|Alert brand of caffeine|alert
Event|Event|SIMPLE_SEGMENT|2295,2300|false|false|false|||alert
Finding|Finding|SIMPLE_SEGMENT|2295,2300|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Functional Concept|SIMPLE_SEGMENT|2295,2300|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Intellectual Product|SIMPLE_SEGMENT|2295,2300|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Event|Event|SIMPLE_SEGMENT|2302,2312|false|false|false|||conversant
Event|Event|SIMPLE_SEGMENT|2322,2328|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|2322,2328|false|false|false|C1554187|Gender Status - Intact|intact
Procedure|Health Care Activity|SIMPLE_SEGMENT|2353,2362|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|SIMPLE_SEGMENT|2363,2367|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2363,2367|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2380,2385|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|2380,2385|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2380,2385|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|2386,2389|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|2395,2398|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2395,2398|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2395,2398|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2405,2408|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2405,2408|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|2405,2408|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2405,2408|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2415,2418|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2415,2418|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|2425,2428|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|2425,2428|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2425,2428|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2425,2428|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2425,2428|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|2432,2435|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2432,2435|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|2432,2435|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|2432,2435|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|2432,2435|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2432,2435|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|2441,2445|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2441,2445|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2460,2463|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2480,2485|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|2480,2485|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2480,2485|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2490,2493|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|SIMPLE_SEGMENT|2490,2493|false|false|false|||PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2490,2493|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2516,2521|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|2516,2521|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2516,2521|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|2516,2529|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2516,2529|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2516,2529|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2522,2529|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|2522,2529|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2522,2529|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|2522,2529|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2522,2529|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2522,2529|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|2576,2580|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2576,2580|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2576,2580|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2606,2611|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|2606,2611|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2606,2611|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2612,2615|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2612,2615|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|2612,2615|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|2612,2615|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|2612,2615|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|2612,2615|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|2612,2615|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2612,2615|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|2620,2623|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2620,2623|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2620,2623|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2620,2623|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|2620,2623|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|2620,2623|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|2620,2623|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2631,2634|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Drug|Enzyme|SIMPLE_SEGMENT|2631,2634|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Event|Event|SIMPLE_SEGMENT|2631,2634|false|false|false|||LDH
Finding|Finding|SIMPLE_SEGMENT|2631,2634|false|false|false|C0851148|Lifetime Drinking History|LDH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2631,2634|false|false|false|C0202113|Lactate dehydrogenase measurement|LDH
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2644,2647|false|false|false|C0010287|Creatine Kinase|CPK
Drug|Enzyme|SIMPLE_SEGMENT|2644,2647|false|false|false|C0010287|Creatine Kinase|CPK
Event|Event|SIMPLE_SEGMENT|2644,2647|false|false|false|||CPK
Finding|Gene or Genome|SIMPLE_SEGMENT|2644,2647|false|false|false|C1418571|PIK3C2A gene|CPK
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2644,2647|false|false|false|C0201973|Creatine kinase measurement|CPK
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2654,2661|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|SIMPLE_SEGMENT|2654,2661|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2689,2694|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|2689,2694|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2689,2694|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2695,2700|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|SIMPLE_SEGMENT|2695,2700|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|SIMPLE_SEGMENT|2695,2700|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2695,2700|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2716,2722|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Drug|Hormone|SIMPLE_SEGMENT|2716,2722|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Finding|Body Substance|SIMPLE_SEGMENT|2731,2740|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|2731,2740|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|2731,2740|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|2731,2740|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|SIMPLE_SEGMENT|2741,2745|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2741,2745|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2758,2763|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|2758,2763|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2758,2763|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|2764,2767|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|2772,2775|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2772,2775|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2772,2775|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2782,2785|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2782,2785|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|2782,2785|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2782,2785|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2792,2795|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2792,2795|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|2803,2806|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|2803,2806|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2803,2806|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2803,2806|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2803,2806|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|2810,2813|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2810,2813|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|2810,2813|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|2810,2813|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|2810,2813|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2810,2813|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|2819,2823|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2819,2823|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2838,2841|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2861,2866|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|2861,2866|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2861,2866|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2883,2888|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|2883,2888|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2883,2888|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Event|SIMPLE_SEGMENT|2912,2913|false|false|false|||-
Drug|Inorganic Chemical|SIMPLE_SEGMENT|2931,2935|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2931,2935|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2931,2935|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2960,2965|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|2960,2965|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2960,2965|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2966,2971|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|SIMPLE_SEGMENT|2966,2971|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|SIMPLE_SEGMENT|2966,2971|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2966,2971|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Event|Event|SIMPLE_SEGMENT|2988,2991|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2988,2991|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Intellectual Product|SIMPLE_SEGMENT|3000,3004|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3005,3029|false|false|false|C0018802|Congestive heart failure|congestive heart failure
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3016,3021|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3016,3021|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|3016,3021|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3016,3029|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Event|Event|SIMPLE_SEGMENT|3022,3029|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|3022,3029|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|3022,3029|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|3022,3029|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3044,3064|false|false|false|C0230147;C4299144|Chest>Mediastinum.superior;Superior mediastinum|superior mediastinum
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3053,3064|false|false|false|C0025066;C4037971|Chest>Mediastinum;Mediastinum|mediastinum
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3053,3064|false|false|false|C0025066;C4037971|Chest>Mediastinum;Mediastinum|mediastinum
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3053,3064|false|false|false|C0153956;C0496915|Benign tumor of mediastinum;Neoplasm of uncertain or unknown behavior of mediastinum|mediastinum
Event|Event|SIMPLE_SEGMENT|3053,3064|false|false|false|||mediastinum
Event|Event|SIMPLE_SEGMENT|3079,3088|false|false|false|||deviation
Finding|Finding|SIMPLE_SEGMENT|3079,3088|false|false|false|C1705236|Protocol Deviation|deviation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3097,3104|false|false|false|C0040578;C4299086|Neck+Chest>Trachea;Trachea|trachea
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3097,3104|false|false|false|C0040580;C0153953;C0154070|Benign neoplasm of trachea;Carcinoma in situ of trachea;Tracheal Diseases|trachea
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3097,3104|false|false|false|C0040580;C0153953;C0154070|Benign neoplasm of trachea;Carcinoma in situ of trachea;Tracheal Diseases|trachea
Event|Event|SIMPLE_SEGMENT|3097,3104|false|false|false|||trachea
Finding|Finding|SIMPLE_SEGMENT|3097,3104|false|false|false|C5848218|trachea findings|trachea
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3097,3104|false|false|false|C0872391|Procedure on trachea|trachea
Event|Event|SIMPLE_SEGMENT|3106,3113|false|false|false|||similar
Event|Event|SIMPLE_SEGMENT|3119,3127|false|false|false|||compared
Event|Event|SIMPLE_SEGMENT|3141,3146|false|false|false|||study
Finding|Intellectual Product|SIMPLE_SEGMENT|3141,3146|false|false|false|C1705923|Study Object|study
Procedure|Research Activity|SIMPLE_SEGMENT|3141,3146|false|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|study
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3148,3156|false|false|false|C2926606||Findings
Finding|Functional Concept|SIMPLE_SEGMENT|3148,3156|false|false|false|C2607943|findings aspects|Findings
Event|Event|SIMPLE_SEGMENT|3162,3169|false|false|false|||reflect
Event|Event|SIMPLE_SEGMENT|3174,3182|false|false|false|||presence
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3174,3182|false|false|false|C0392148|Providing presence (regime/therapy)|presence
Finding|Finding|SIMPLE_SEGMENT|3174,3185|false|false|false|C0150312|Present|presence of
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3188,3195|false|false|false|C0040132|Thyroid Gland|thyroid
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3188,3195|false|false|false|C0040128|Thyroid Diseases|thyroid
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3188,3195|false|false|false|C0040134;C3540038;C5781115|THYROID;THYROID DIAGNOSTIC RADIOPHARMACEUTICALS;thyroid (USP)|thyroid
Drug|Hormone|SIMPLE_SEGMENT|3188,3195|false|false|false|C0040134;C3540038;C5781115|THYROID;THYROID DIAGNOSTIC RADIOPHARMACEUTICALS;thyroid (USP)|thyroid
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|3188,3195|false|false|false|C0040134;C3540038;C5781115|THYROID;THYROID DIAGNOSTIC RADIOPHARMACEUTICALS;thyroid (USP)|thyroid
Drug|Organic Chemical|SIMPLE_SEGMENT|3188,3195|false|false|false|C0040134;C3540038;C5781115|THYROID;THYROID DIAGNOSTIC RADIOPHARMACEUTICALS;thyroid (USP)|thyroid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3188,3195|false|false|false|C0040134;C3540038;C5781115|THYROID;THYROID DIAGNOSTIC RADIOPHARMACEUTICALS;thyroid (USP)|thyroid
Procedure|Health Care Activity|SIMPLE_SEGMENT|3188,3195|false|false|false|C2228489|examination of thyroid|thyroid
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3188,3202|false|false|false|C0018021|Goiter|thyroid goiter
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3196,3202|false|false|false|C0018021|Goiter|goiter
Event|Event|SIMPLE_SEGMENT|3196,3202|false|false|false|||goiter
Event|Event|SIMPLE_SEGMENT|3208,3216|false|false|false|||clinical
Finding|Intellectual Product|SIMPLE_SEGMENT|3208,3216|false|false|false|C1315013|Clinical NEC (not elsewhere classified in LNC)|clinical
Event|Event|SIMPLE_SEGMENT|3218,3229|false|false|false|||correlation
Event|Event|SIMPLE_SEGMENT|3233,3244|false|false|false|||recommended
Event|Event|SIMPLE_SEGMENT|3253,3262|false|false|false|||indicated
Event|Event|SIMPLE_SEGMENT|3279,3288|false|false|false|||confirmed
Event|Event|SIMPLE_SEGMENT|3296,3298|false|false|false|||CT
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3306,3311|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|3306,3311|false|false|false|C0741025|Chest problem|chest
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3320,3325|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|spine
Anatomy|Cell Component|SIMPLE_SEGMENT|3320,3325|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|spine
Finding|Finding|SIMPLE_SEGMENT|3320,3325|false|false|false|C0150920|Spine Problem|spine
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3326,3330|false|false|false|C1561572;C1704608|Film Dosage Form;film - layer|film
Drug|Substance|SIMPLE_SEGMENT|3326,3330|false|false|false|C1561572;C1704608|Film Dosage Form;film - layer|film
Event|Event|SIMPLE_SEGMENT|3326,3330|false|false|false|||film
Finding|Intellectual Product|SIMPLE_SEGMENT|3326,3330|false|false|false|C4019020||film
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3357,3363|false|false|false|C0024090|Lumbar Region|lumbar
Finding|Gene or Genome|SIMPLE_SEGMENT|3364,3368|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Intellectual Product|SIMPLE_SEGMENT|3364,3368|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3369,3378|false|false|false|C0549207|Bone structure of spine|vertebral
Event|Event|SIMPLE_SEGMENT|3382,3388|false|false|false|||bodies
Event|Event|SIMPLE_SEGMENT|3393,3400|false|false|false|||present
Finding|Finding|SIMPLE_SEGMENT|3393,3400|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|SIMPLE_SEGMENT|3393,3400|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Functional Concept|SIMPLE_SEGMENT|3423,3435|false|false|false|C0011164;C1880269|Abnormal degeneration;biologic degeneration|degenerative
Finding|Pathologic Function|SIMPLE_SEGMENT|3423,3435|false|false|false|C0011164;C1880269|Abnormal degeneration;biologic degeneration|degenerative
Finding|Pathologic Function|SIMPLE_SEGMENT|3423,3443|false|false|false|C0011164|Abnormal degeneration|degenerative changes
Event|Event|SIMPLE_SEGMENT|3436,3443|false|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|3436,3443|false|false|false|C0392747|Changing|changes
Event|Event|SIMPLE_SEGMENT|3451,3455|false|false|false|||loss
Finding|Finding|SIMPLE_SEGMENT|3451,3455|false|false|false|C5890125|Loss (adaptation)|loss
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3459,3473|false|false|false|C0442106|Intervertebral|intervertebral
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3459,3478|false|false|false|C0021815|Intervertebral disc structure|intervertebral disc
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3474,3478|false|false|false|C1556138;C1621443|Disc - Body Part;death-inducing signaling complex location|disc
Anatomy|Cell Component|SIMPLE_SEGMENT|3474,3478|false|false|false|C1556138;C1621443|Disc - Body Part;death-inducing signaling complex location|disc
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3474,3478|false|false|false|C0993608|Disk Drug Form|disc
Finding|Finding|SIMPLE_SEGMENT|3474,3478|false|false|false|C1444662;C1696131|Disc (List bullets);Discontinued|disc
Finding|Intellectual Product|SIMPLE_SEGMENT|3474,3478|false|false|false|C1444662;C1696131|Disc (List bullets);Discontinued|disc
Event|Event|SIMPLE_SEGMENT|3479,3485|false|false|false|||height
Finding|Functional Concept|SIMPLE_SEGMENT|3516,3525|false|false|false|C0036429;C0334135|Sclerosis;Sclerotic (qualifier value)|sclerotic
Finding|Pathologic Function|SIMPLE_SEGMENT|3516,3525|false|false|false|C0036429;C0334135|Sclerosis;Sclerotic (qualifier value)|sclerotic
Event|Event|SIMPLE_SEGMENT|3526,3533|false|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|3526,3533|false|false|false|C0392747|Changing|changes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3539,3547|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3548,3558|false|false|false|C0015302;C1956089|External hyperostosis;Osteophyte|osteophyte
Finding|Pathologic Function|SIMPLE_SEGMENT|3548,3568|false|false|false|C5442360|Osteophyte formation|osteophyte formation
Event|Event|SIMPLE_SEGMENT|3559,3568|false|false|false|||formation
Finding|Functional Concept|SIMPLE_SEGMENT|3559,3568|false|false|false|C1522492|Formation|formation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|3559,3568|false|false|false|C0220781|Anabolism|formation
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|3583,3591|true|false|false|C0016658|Fracture|fracture
Event|Event|SIMPLE_SEGMENT|3583,3591|false|false|false|||fracture
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3595,3604|false|false|false|C0549207|Bone structure of spine|vertebral
Finding|Pathologic Function|SIMPLE_SEGMENT|3595,3616|true|false|false|C0262431|Compression fracture of vertebral column|vertebral compression
Event|Event|SIMPLE_SEGMENT|3605,3616|false|false|false|||compression
Finding|Functional Concept|SIMPLE_SEGMENT|3605,3616|true|false|false|C0332459;C4551657|Compressed structure|compression
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3605,3616|true|false|false|C0728907|Compression|compression
Procedure|Machine Activity|SIMPLE_SEGMENT|3605,3616|true|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3605,3616|true|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|3617,3626|true|false|false|C0000768;C0302142|Congenital Abnormality;Deformity|deformity
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|3617,3626|true|false|false|C0000768;C0302142|Congenital Abnormality;Deformity|deformity
Event|Event|SIMPLE_SEGMENT|3617,3626|false|false|false|||deformity
Finding|Finding|SIMPLE_SEGMENT|3617,3626|true|false|false|C2117111||deformity
Event|Event|SIMPLE_SEGMENT|3628,3638|false|false|false|||identified
Finding|Finding|SIMPLE_SEGMENT|3649,3655|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|3649,3655|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Intellectual Product|SIMPLE_SEGMENT|3656,3660|false|false|false|C1547225|Mild Severity of Illness Code|mild
Event|Event|SIMPLE_SEGMENT|3661,3666|false|false|false|||grade
Finding|Classification|SIMPLE_SEGMENT|3661,3666|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Finding|Finding|SIMPLE_SEGMENT|3661,3666|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Finding|Finding|SIMPLE_SEGMENT|3661,3668|false|false|false|C0475269;C0547053;C0687695;C4284291|First grade in elementary school;Grade 1 (qualifier value);Simpson Grade 1;Tumor grade G1|grade 1
Finding|Intellectual Product|SIMPLE_SEGMENT|3661,3668|false|false|false|C0475269;C0547053;C0687695;C4284291|First grade in elementary school;Grade 1 (qualifier value);Simpson Grade 1;Tumor grade G1|grade 1
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3679,3694|false|false|false|C1504511|Anterolisthesis|anterolisthesis
Event|Event|SIMPLE_SEGMENT|3679,3694|false|false|false|||anterolisthesis
Finding|Finding|SIMPLE_SEGMENT|3705,3711|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|3705,3711|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|SIMPLE_SEGMENT|3712,3724|false|false|false|||degenerative
Finding|Functional Concept|SIMPLE_SEGMENT|3712,3724|false|true|false|C0011164;C1880269|Abnormal degeneration;biologic degeneration|degenerative
Finding|Pathologic Function|SIMPLE_SEGMENT|3712,3724|false|true|false|C0011164;C1880269|Abnormal degeneration;biologic degeneration|degenerative
Event|Event|SIMPLE_SEGMENT|3728,3736|false|false|false|||etiology
Finding|Conceptual Entity|SIMPLE_SEGMENT|3728,3736|false|true|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|etiology
Finding|Functional Concept|SIMPLE_SEGMENT|3728,3736|false|true|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|etiology
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3738,3743|false|false|false|C0222679|Structure of articular surface of bone|Facet
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3745,3757|false|false|false|C0263630||hypertrophic
Event|Event|SIMPLE_SEGMENT|3745,3757|false|false|false|||hypertrophic
Finding|Functional Concept|SIMPLE_SEGMENT|3745,3757|false|false|false|C0020564;C0333959|Hypertrophic;Hypertrophy|hypertrophic
Finding|Pathologic Function|SIMPLE_SEGMENT|3745,3757|false|false|false|C0020564;C0333959|Hypertrophic;Hypertrophy|hypertrophic
Event|Event|SIMPLE_SEGMENT|3758,3765|false|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|3758,3765|false|false|false|C0392747|Changing|changes
Event|Event|SIMPLE_SEGMENT|3770,3775|false|false|false|||noted
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3787,3792|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|3787,3792|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3793,3799|false|false|false|C0024090|Lumbar Region|lumbar
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3793,3805|false|false|false|C0024091;C3887615|Bone structure of lumbar vertebra;Lumbar spine structure|lumbar spine
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3793,3805|false|false|false|C0024091;C3887615|Bone structure of lumbar vertebra;Lumbar spine structure|lumbar spine
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3800,3805|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|spine
Anatomy|Cell Component|SIMPLE_SEGMENT|3800,3805|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|spine
Finding|Finding|SIMPLE_SEGMENT|3800,3805|false|false|false|C0150920|Spine Problem|spine
Event|Event|SIMPLE_SEGMENT|3817,3826|false|false|false|||affecting
Event|Event|SIMPLE_SEGMENT|3841,3847|false|false|false|||levels
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3849,3857|false|false|false|C0005847|Blood Vessel|Vascular
Event|Event|SIMPLE_SEGMENT|3859,3873|false|false|false|||calcifications
Finding|Finding|SIMPLE_SEGMENT|3859,3873|true|false|false|C0006660;C2242558|Pathologic calcification, calcified structure;Physiologic calcification|calcifications
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3859,3873|true|false|false|C0006660;C2242558|Pathologic calcification, calcified structure;Physiologic calcification|calcifications
Event|Event|SIMPLE_SEGMENT|3878,3888|false|false|false|||visualized
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3894,3904|false|false|false|C0555898|sacroiliac|sacroiliac
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|3894,3911|false|false|false|C0036036|Sacroiliac joint structure|sacroiliac joints
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|3905,3911|false|false|false|C0022417;C0392905|Articular system;Joints|joints
Anatomy|Body System|SIMPLE_SEGMENT|3905,3911|false|false|false|C0022417;C0392905|Articular system;Joints|joints
Event|Event|SIMPLE_SEGMENT|3921,3930|false|false|false|||diastatic
Event|Event|SIMPLE_SEGMENT|3934,3944|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|3934,3944|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|3934,3944|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|3949,3957|true|false|false|C0016658|Fracture|fracture
Event|Event|SIMPLE_SEGMENT|3949,3957|false|false|false|||fracture
Event|Event|SIMPLE_SEGMENT|3958,3968|false|false|false|||identified
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3973,3980|false|false|false|C0881943||CT head
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3973,3980|false|false|false|C0202691|CAT scan of head|CT head
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3976,3980|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3976,3980|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3976,3980|false|false|false|C0362076|Problems with head|head
Event|Event|SIMPLE_SEGMENT|3976,3980|false|false|false|||head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3976,3980|false|false|false|C0876917|Procedure on head|head
Finding|Intellectual Product|SIMPLE_SEGMENT|3998,4003|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4004,4016|false|false|false|C0524466|Intracranial|intracranial
Finding|Functional Concept|SIMPLE_SEGMENT|4004,4016|false|false|false|C1522213|Intracranial Route of Administration|intracranial
Finding|Pathologic Function|SIMPLE_SEGMENT|4004,4027|true|false|false|C0151699|Intracranial Hemorrhage|intracranial hemorrhage
Event|Event|SIMPLE_SEGMENT|4017,4027|false|false|false|||hemorrhage
Finding|Pathologic Function|SIMPLE_SEGMENT|4017,4027|true|false|false|C0019080|Hemorrhage|hemorrhage
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4029,4034|true|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|4029,4034|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|4029,4034|true|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|4038,4043|false|false|false|||acute
Finding|Intellectual Product|SIMPLE_SEGMENT|4038,4043|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4045,4053|false|false|false|C0005847|Blood Vessel|vascular
Event|Event|SIMPLE_SEGMENT|4067,4077|false|false|false|||infarction
Finding|Pathologic Function|SIMPLE_SEGMENT|4067,4077|false|false|false|C0021308|Infarction|infarction
Event|Event|SIMPLE_SEGMENT|4079,4083|false|false|false|||Note
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4105,4121|false|false|false|C0014068|Encephalomalacia|encephalomalacia
Event|Event|SIMPLE_SEGMENT|4105,4121|false|false|false|||encephalomalacia
Event|Event|SIMPLE_SEGMENT|4122,4131|false|false|false|||involving
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4136,4149|false|false|false|C0030560|Parietal Lobe|parietal lobe
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4136,4149|false|false|false|C0153637|Malignant neoplasm of parietal lobe|parietal lobe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4145,4149|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|SIMPLE_SEGMENT|4145,4149|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Finding|Functional Concept|SIMPLE_SEGMENT|4157,4161|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Event|Event|SIMPLE_SEGMENT|4177,4186|false|false|false|||unchanged
Finding|Finding|SIMPLE_SEGMENT|4177,4186|false|false|false|C0442739||unchanged
Event|Governmental or Regulatory Activity|SIMPLE_SEGMENT|4198,4202|false|false|false|C1510751|Academic Research Enhancement Awards|area
Finding|Functional Concept|SIMPLE_SEGMENT|4225,4230|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Event|Event|SIMPLE_SEGMENT|4232,4240|false|false|false|||adjacent
Event|Event|SIMPLE_SEGMENT|4267,4276|false|false|false|||unchanged
Finding|Finding|SIMPLE_SEGMENT|4267,4276|false|false|false|C0442739||unchanged
Finding|Functional Concept|SIMPLE_SEGMENT|4285,4289|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4299,4310|false|false|false|C0025286|Meningioma|meningiomas
Event|Event|SIMPLE_SEGMENT|4299,4310|false|false|false|||meningiomas
Event|Event|SIMPLE_SEGMENT|4345,4354|false|false|false|||calcified
Finding|Idea or Concept|SIMPLE_SEGMENT|4361,4367|false|false|false|C1550462|Observation Interpretation - better|better
Event|Event|SIMPLE_SEGMENT|4368,4376|false|false|false|||depicted
Event|Event|SIMPLE_SEGMENT|4390,4393|false|false|false|||MRI
Finding|Gene or Genome|SIMPLE_SEGMENT|4390,4393|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4390,4393|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|SIMPLE_SEGMENT|4390,4393|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4410,4420|false|false|false|C0018827|Heart Ventricle|Ventricles
Finding|Finding|SIMPLE_SEGMENT|4457,4480|false|false|false|C5883508|Parenchymal volume loss|parenchymal volume loss
Finding|Intellectual Product|SIMPLE_SEGMENT|4469,4475|false|false|false|C1705102|Volume (publication)|volume
Event|Event|SIMPLE_SEGMENT|4476,4480|false|false|false|||loss
Finding|Finding|SIMPLE_SEGMENT|4476,4480|false|false|false|C5890125|Loss (adaptation)|loss
Finding|Functional Concept|SIMPLE_SEGMENT|4499,4514|false|false|false|C0333482|atherosclerotic|atherosclerotic
Event|Event|SIMPLE_SEGMENT|4515,4528|false|false|false|||calcification
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4515,4528|false|false|false|C0006660;C0006663;C1533591|Calcification;Calcinosis;Physiologic calcification|calcification
Finding|Pathologic Function|SIMPLE_SEGMENT|4515,4528|false|false|false|C0006660;C0006663;C1533591|Calcification;Calcinosis;Physiologic calcification|calcification
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4536,4543|false|false|false|C0007272|Carotid Arteries|carotid
Event|Event|SIMPLE_SEGMENT|4544,4551|false|false|false|||siphons
Finding|Finding|SIMPLE_SEGMENT|4568,4572|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|4587,4595|false|false|false|||segments
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|4610,4618|false|false|false|C0016658|Fracture|fracture
Event|Event|SIMPLE_SEGMENT|4610,4618|false|false|false|||fracture
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4624,4631|false|false|false|C0446908;C1521748;C4266570|Head>Mastoid;Mastoid process|mastoid
Procedure|Health Care Activity|SIMPLE_SEGMENT|4624,4631|false|false|false|C2228459|examination of mastoid region|mastoid
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4624,4641|false|false|false|C0229427|Pneumatic mastoid cell|mastoid air cells
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4632,4635|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4632,4635|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|SIMPLE_SEGMENT|4632,4635|false|false|false|C0001861;C3536832|Air (substance);air|air
Finding|Finding|SIMPLE_SEGMENT|4632,4635|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|SIMPLE_SEGMENT|4632,4635|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|SIMPLE_SEGMENT|4632,4635|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Anatomy|Cell|SIMPLE_SEGMENT|4636,4641|false|false|false|C0007634|Cells|cells
Event|Event|SIMPLE_SEGMENT|4646,4651|false|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|4646,4651|false|false|false|C1550016|Remote control command - Clear|clear
Event|Event|SIMPLE_SEGMENT|4654,4664|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|4654,4664|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|4654,4664|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|4669,4674|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4675,4687|false|false|false|C0524466|Intracranial|intracranial
Finding|Functional Concept|SIMPLE_SEGMENT|4675,4687|false|false|false|C1522213|Intracranial Route of Administration|intracranial
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|4688,4699|false|false|false|C0000768|Congenital Abnormality|abnormality
Event|Event|SIMPLE_SEGMENT|4688,4699|false|false|false|||abnormality
Finding|Finding|SIMPLE_SEGMENT|4688,4699|false|false|false|C1704258|Abnormality|abnormality
Event|Event|SIMPLE_SEGMENT|4705,4714|false|false|false|||unchanged
Finding|Finding|SIMPLE_SEGMENT|4705,4714|false|false|false|C0442739||unchanged
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4716,4724|false|false|false|C2926606||findings
Event|Event|SIMPLE_SEGMENT|4716,4724|false|false|false|||findings
Finding|Functional Concept|SIMPLE_SEGMENT|4716,4724|false|false|false|C2607943|findings aspects|findings
Event|Event|SIMPLE_SEGMENT|4738,4746|false|false|false|||infarcts
Finding|Pathologic Function|SIMPLE_SEGMENT|4738,4746|false|false|false|C0021308|Infarction|infarcts
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4751,4762|false|false|false|C0025286|Meningioma|meningiomas
Event|Event|SIMPLE_SEGMENT|4751,4762|false|false|false|||meningiomas
Event|Event|SIMPLE_SEGMENT|4777,4786|false|false|false|||Waveforms
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|4777,4786|false|false|false|C0450448|Waveforms|Waveforms
Finding|Functional Concept|SIMPLE_SEGMENT|4794,4800|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Finding|Intellectual Product|SIMPLE_SEGMENT|4794,4800|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4801,4808|false|false|false|C0015811|Femur|femoral
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4801,4814|false|false|false|C0015809|Femoral vein|femoral veins
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4809,4814|false|false|false|C0042449|Veins|veins
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4809,4814|false|false|false|C0398102|Procedure on vein|veins
Event|Event|SIMPLE_SEGMENT|4819,4828|false|false|false|||symmetric
Finding|Conceptual Entity|SIMPLE_SEGMENT|4819,4828|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|SIMPLE_SEGMENT|4819,4828|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Event|Event|SIMPLE_SEGMENT|4859,4868|false|false|false|||responses
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4872,4880|false|false|false|C0750122|valsalva|Valsalva
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4872,4890|false|false|false|C0042293|Valsalva Maneuver|Valsalva maneuvers
Event|Event|SIMPLE_SEGMENT|4881,4890|false|false|false|||maneuvers
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4900,4905|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|4900,4905|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4907,4918|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Finding|Functional Concept|SIMPLE_SEGMENT|4924,4930|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Finding|Intellectual Product|SIMPLE_SEGMENT|4924,4930|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4931,4938|false|false|false|C0015811|Femur|femoral
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4940,4948|false|false|false|C4489236|Proximal Resection Margin|proximal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4981,4988|false|false|false|C0015811|Femur|femoral
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4993,5002|false|false|false|C0442037|popliteal|popliteal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4993,5008|false|false|false|C0032652|Structure of popliteal vein|popliteal veins
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5003,5008|false|false|false|C0042449|Veins|veins
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5003,5008|false|false|false|C0398102|Procedure on vein|veins
Event|Event|SIMPLE_SEGMENT|5013,5019|false|false|false|||normal
Event|Event|SIMPLE_SEGMENT|5038,5053|false|false|false|||compressibility
Event|Event|SIMPLE_SEGMENT|5068,5072|false|false|false|||flow
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|5068,5072|false|false|false|C0806140|Flow|flow
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5076,5081|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|color
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|5076,5081|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|color
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5076,5089|false|false|false|C0474781|Color doppler ultrasound|color Doppler
Event|Event|SIMPLE_SEGMENT|5082,5089|false|false|false|||Doppler
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5082,5089|false|false|false|C0554756|Doppler studies|Doppler
Event|Event|SIMPLE_SEGMENT|5091,5099|false|false|false|||analysis
Finding|Functional Concept|SIMPLE_SEGMENT|5091,5099|false|false|false|C1524024|analysis aspect|analysis
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5091,5099|false|false|false|C0002778;C0936012|Analysis;Analysis of substances|analysis
Procedure|Research Activity|SIMPLE_SEGMENT|5091,5099|false|false|false|C0002778;C0936012|Analysis;Analysis of substances|analysis
Event|Event|SIMPLE_SEGMENT|5104,5112|false|false|false|||response
Finding|Finding|SIMPLE_SEGMENT|5104,5112|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Intellectual Product|SIMPLE_SEGMENT|5104,5112|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Mental Process|SIMPLE_SEGMENT|5104,5112|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|5116,5124|false|false|false|C0450448|Waveforms|waveform
Event|Event|SIMPLE_SEGMENT|5125,5137|false|false|false|||augmentation
Finding|Finding|SIMPLE_SEGMENT|5125,5137|false|false|false|C0332509|Increased size (finding)|augmentation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5125,5137|false|false|false|C1293122|Augmentation procedure|augmentation
Event|Event|SIMPLE_SEGMENT|5153,5157|false|false|false|||flow
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|5153,5157|false|false|false|C0806140|Flow|flow
Event|Event|SIMPLE_SEGMENT|5166,5176|false|false|false|||visualized
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5184,5193|false|false|false|C0751438|Posterior pituitary disease|posterior
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5194,5200|false|false|false|C0040184|Bone structure of tibia|tibial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5215,5220|false|false|false|C0042449|Veins|veins
Event|Event|SIMPLE_SEGMENT|5215,5220|false|false|false|||veins
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5215,5220|false|false|false|C0398102|Procedure on vein|veins
Event|Event|SIMPLE_SEGMENT|5229,5235|false|false|false|||calves
Event|Event|SIMPLE_SEGMENT|5237,5247|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|5237,5247|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|5237,5247|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5252,5256|false|false|false|C4318566|Deep Resection Margin|deep
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5252,5274|true|false|false|C0149871|Deep Vein Thrombosis|deep venous thrombosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5257,5263|false|false|false|C0042449|Veins|venous
Finding|Finding|SIMPLE_SEGMENT|5257,5274|true|false|false|C0042487;C0517555|Venous Thrombosis;Venous thrombosis after immobility|venous thrombosis
Finding|Pathologic Function|SIMPLE_SEGMENT|5257,5274|true|false|false|C0042487;C0517555|Venous Thrombosis;Venous thrombosis after immobility|venous thrombosis
Event|Event|SIMPLE_SEGMENT|5264,5274|false|false|false|||thrombosis
Finding|Pathologic Function|SIMPLE_SEGMENT|5264,5274|true|false|false|C0040053|Thrombosis|thrombosis
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5285,5290|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|5285,5290|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5285,5300|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5291,5300|false|false|false|C0015385|Limb structure|extremity
Event|Event|SIMPLE_SEGMENT|5308,5320|false|false|false|||MICROBIOLOGY
Finding|Functional Concept|SIMPLE_SEGMENT|5308,5320|false|false|false|C0025953;C1571921;C4049106|Microbiological;Microbiology - Laboratory Class;Microbiology Diagnostic Service Section ID|MICROBIOLOGY
Finding|Intellectual Product|SIMPLE_SEGMENT|5308,5320|false|false|false|C0025953;C1571921;C4049106|Microbiological;Microbiology - Laboratory Class;Microbiology Diagnostic Service Section ID|MICROBIOLOGY
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5308,5320|false|false|false|C0085672|Microbiology procedure|MICROBIOLOGY
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5328,5333|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Event|Event|SIMPLE_SEGMENT|5328,5333|false|false|false|||Blood
Finding|Body Substance|SIMPLE_SEGMENT|5328,5333|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5328,5341|false|false|false|C0200949|Blood culture|Blood culture
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5334,5341|false|false|false|C1706355|Culture Dose Form|culture
Event|Event|SIMPLE_SEGMENT|5334,5341|false|false|false|||culture
Finding|Functional Concept|SIMPLE_SEGMENT|5334,5341|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Finding|Idea or Concept|SIMPLE_SEGMENT|5334,5341|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5334,5341|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|culture
Event|Event|SIMPLE_SEGMENT|5347,5353|false|false|false|||growth
Finding|Finding|SIMPLE_SEGMENT|5347,5353|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5347,5353|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Finding|Organism Function|SIMPLE_SEGMENT|5347,5353|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Finding|Physiologic Function|SIMPLE_SEGMENT|5347,5353|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|5347,5353|true|false|false|C2911660|Growth action|growth
Finding|Intellectual Product|SIMPLE_SEGMENT|5365,5370|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|5371,5379|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5371,5386|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|5371,5386|false|false|false|C0489547|Hospital course|Hospital Course
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5406,5410|false|false|false|C0004238|Atrial Fibrillation|afib
Event|Event|SIMPLE_SEGMENT|5406,5410|false|false|false|||afib
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5406,5410|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|afib
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5416,5419|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5416,5419|false|false|false|C0018802|Congestive heart failure|CHF
Event|Event|SIMPLE_SEGMENT|5416,5419|false|false|false|||CHF
Event|Event|SIMPLE_SEGMENT|5420,5430|false|false|false|||presenting
Procedure|Health Care Activity|SIMPLE_SEGMENT|5436,5440|false|false|false|C1315068|Pulmonary ventilator management|pulm
Finding|Pathologic Function|SIMPLE_SEGMENT|5436,5446|false|false|false|C0034063|Pulmonary Edema|pulm edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5441,5446|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|5441,5446|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|5441,5446|false|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|5452,5461|false|false|false|||worsening
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5466,5471|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|5466,5471|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|5466,5471|false|false|false|C0013604|Edema|edema
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5477,5480|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5477,5480|false|false|false|C0018802|Congestive heart failure|CHF
Event|Event|SIMPLE_SEGMENT|5477,5480|false|false|false|||CHF
Finding|Intellectual Product|SIMPLE_SEGMENT|5492,5497|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Intellectual Product|SIMPLE_SEGMENT|5501,5508|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|5501,5508|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Event|Event|SIMPLE_SEGMENT|5509,5518|false|false|false|||worsening
Finding|Idea or Concept|SIMPLE_SEGMENT|5509,5518|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5522,5531|false|false|false|C0012000|Diastole|diastolic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5533,5557|false|false|false|C0018802|Congestive heart failure|congestive heart failure
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5544,5549|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5544,5549|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|5544,5549|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5544,5557|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Event|Event|SIMPLE_SEGMENT|5550,5557|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|5550,5557|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|5550,5557|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|5550,5557|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5571,5575|false|false|false|C0428772|Left ventricular ejection fraction|LVEF
Event|Event|SIMPLE_SEGMENT|5571,5575|false|false|false|||LVEF
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5571,5575|false|false|false|C3837267|LVEF (procedure)|LVEF
Event|Event|SIMPLE_SEGMENT|5594,5602|false|false|false|||decrease
Finding|Finding|SIMPLE_SEGMENT|5594,5602|false|false|false|C0392756|Reduced|decrease
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5606,5614|false|false|false|C0080078|Range of Motion, Articular|mobility
Event|Event|SIMPLE_SEGMENT|5606,5614|false|false|false|||mobility
Finding|Finding|SIMPLE_SEGMENT|5606,5614|false|false|false|C0425245|Mobility finding|mobility
Event|Event|SIMPLE_SEGMENT|5620,5624|false|false|false|||fall
Finding|Finding|SIMPLE_SEGMENT|5620,5624|false|false|false|C0085639|Falls|fall
Finding|Finding|SIMPLE_SEGMENT|5644,5650|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Idea or Concept|SIMPLE_SEGMENT|5644,5650|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Event|Event|SIMPLE_SEGMENT|5656,5665|false|false|false|||worsening
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5666,5671|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|5666,5671|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|5666,5671|false|false|false|C0013604|Edema|edema
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5682,5692|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|5682,5692|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|5682,5692|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Finding|Individual Behavior|SIMPLE_SEGMENT|5682,5707|false|false|false|C3489773|Medication Compliance|medication non-compliance
Event|Event|SIMPLE_SEGMENT|5716,5725|false|false|false|||worsening
Finding|Idea or Concept|SIMPLE_SEGMENT|5716,5725|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5733,5739|false|false|false|C0003483|Aorta|aortic
Finding|Pathologic Function|SIMPLE_SEGMENT|5733,5748|false|false|false|C0003507|Aortic Valve Stenosis|aortic stenosis
Event|Event|SIMPLE_SEGMENT|5740,5748|false|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|5740,5748|false|false|false|C1261287|Stenosis|stenosis
Event|Event|SIMPLE_SEGMENT|5766,5770|false|false|false|||echo
Procedure|Health Care Activity|SIMPLE_SEGMENT|5766,5770|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5766,5770|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Event|Event|SIMPLE_SEGMENT|5796,5807|false|false|false|||recommended
Event|Event|SIMPLE_SEGMENT|5816,5824|false|false|false|||repeated
Event|Event|SIMPLE_SEGMENT|5831,5841|false|false|false|||outpatient
Finding|Classification|SIMPLE_SEGMENT|5831,5841|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|5831,5841|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|SIMPLE_SEGMENT|5857,5864|false|false|false|||hypoxic
Finding|Pathologic Function|SIMPLE_SEGMENT|5857,5864|false|false|false|C0242184|Hypoxia|hypoxic
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5873,5877|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5873,5877|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5873,5877|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|5873,5877|false|false|false|C0740941|Lung Problem|lung
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5873,5882|false|false|false|C2228454|examination of lungs|lung exam
Event|Event|SIMPLE_SEGMENT|5878,5882|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|5878,5882|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|5878,5882|false|false|false|C0582103|Medical Examination|exam
Event|Event|SIMPLE_SEGMENT|5883,5892|false|false|false|||suggested
Event|Event|SIMPLE_SEGMENT|5903,5907|false|false|false|||pulm
Procedure|Health Care Activity|SIMPLE_SEGMENT|5903,5907|false|false|false|C1315068|Pulmonary ventilator management|pulm
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5909,5914|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|5909,5914|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|5909,5914|false|false|false|C0013604|Edema|edema
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5920,5924|false|false|false|C1140621|Leg|legs
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5920,5924|false|false|false|C5781420||legs
Event|Event|SIMPLE_SEGMENT|5930,5938|false|false|false|||elevated
Finding|Functional Concept|SIMPLE_SEGMENT|5943,5954|false|false|false|C0332459;C4551657|Compressed structure|compression
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|5943,5954|false|false|false|C0728907|Compression|compression
Procedure|Machine Activity|SIMPLE_SEGMENT|5943,5954|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5943,5954|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Event|Event|SIMPLE_SEGMENT|5955,5964|false|false|false|||stockings
Event|Event|SIMPLE_SEGMENT|5971,5975|false|false|false|||used
Drug|Organic Chemical|SIMPLE_SEGMENT|5981,5990|false|false|false|C0076840|torsemide|torsemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5981,5990|false|false|false|C0076840|torsemide|torsemide
Event|Event|SIMPLE_SEGMENT|5981,5990|false|false|false|||torsemide
Event|Event|SIMPLE_SEGMENT|5995,6000|false|false|false|||dosed
Event|Event|SIMPLE_SEGMENT|6028,6035|false|false|false|||unclear
Event|Event|SIMPLE_SEGMENT|6052,6060|false|false|false|||increase
Finding|Functional Concept|SIMPLE_SEGMENT|6052,6060|false|false|false|C0442805|Increase|increase
Event|Event|SIMPLE_SEGMENT|6082,6086|false|false|false|||dose
Finding|Body Substance|SIMPLE_SEGMENT|6097,6104|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6097,6104|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6097,6104|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|6119,6125|false|false|false|||unable
Finding|Finding|SIMPLE_SEGMENT|6119,6125|false|false|false|C1299582|Unable|unable
Event|Activity|SIMPLE_SEGMENT|6129,6136|false|false|false|C2986669|Clarify|clarify
Event|Event|SIMPLE_SEGMENT|6129,6136|false|false|false|||clarify
Event|Event|SIMPLE_SEGMENT|6148,6154|false|false|false|||slight
Finding|Finding|SIMPLE_SEGMENT|6148,6154|false|false|false|C5202796|Intensity and Distress 1|slight
Event|Event|SIMPLE_SEGMENT|6156,6167|false|false|false|||improvement
Finding|Conceptual Entity|SIMPLE_SEGMENT|6156,6167|false|false|false|C2986411|Improvement|improvement
Event|Event|SIMPLE_SEGMENT|6171,6179|false|false|false|||swelling
Finding|Finding|SIMPLE_SEGMENT|6171,6179|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|6171,6179|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Event|Event|SIMPLE_SEGMENT|6183,6192|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|6183,6192|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6183,6192|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6183,6192|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6183,6192|false|false|false|C0030685|Patient Discharge|discharge
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|6205,6210|false|false|false|C0000921|Accidental Falls|FALLS
Event|Event|SIMPLE_SEGMENT|6205,6210|false|false|false|||FALLS
Finding|Finding|SIMPLE_SEGMENT|6205,6210|false|false|false|C0085639|Falls|FALLS
Finding|Body Substance|SIMPLE_SEGMENT|6212,6219|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6212,6219|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6212,6219|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|6220,6227|false|false|false|||reports
Event|Event|SIMPLE_SEGMENT|6228,6235|false|false|false|||falling
Finding|Finding|SIMPLE_SEGMENT|6251,6258|false|false|false|C4534363|At home|at home
Event|Event|SIMPLE_SEGMENT|6254,6258|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|6254,6258|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|6254,6258|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|6254,6258|false|false|false|C1553498|home health encounter|home
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6269,6273|false|false|false|C0077275|triptorelin|trip
Drug|Hormone|SIMPLE_SEGMENT|6269,6273|false|false|false|C0077275|triptorelin|trip
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6269,6273|false|false|false|C0077275|triptorelin|trip
Event|Event|SIMPLE_SEGMENT|6269,6273|false|false|false|||trip
Finding|Gene or Genome|SIMPLE_SEGMENT|6269,6273|false|false|false|C1416921;C2239819;C2608049;C4085339|LRRFIP1 gene;PIK3IP1 gene;TRAIP gene;TRAIP wt Allele|trip
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|6269,6273|false|false|false|C0221188|Tripping|trip
Event|Event|SIMPLE_SEGMENT|6282,6291|false|false|false|||evaluated
Finding|Finding|SIMPLE_SEGMENT|6295,6303|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Finding|Functional Concept|SIMPLE_SEGMENT|6295,6303|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|6295,6303|false|false|false|C0031809|Physical Examination|physical
Finding|Intellectual Product|SIMPLE_SEGMENT|6295,6311|false|false|false|C1547999|Diagnostic Service Section ID - Physical Therapy|physical therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6295,6311|false|false|false|C0949766|Physical therapy|physical therapy
Event|Event|SIMPLE_SEGMENT|6304,6311|false|false|false|||therapy
Finding|Finding|SIMPLE_SEGMENT|6304,6311|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|SIMPLE_SEGMENT|6304,6311|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6304,6311|false|false|false|C0087111|Therapeutic procedure|therapy
Event|Event|SIMPLE_SEGMENT|6317,6321|false|false|false|||felt
Event|Event|SIMPLE_SEGMENT|6329,6337|false|false|false|||unsteady
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6345,6349|false|false|false|C0016504|Foot|feet
Event|Event|SIMPLE_SEGMENT|6354,6358|false|false|false|||safe
Finding|Intellectual Product|SIMPLE_SEGMENT|6354,6358|false|false|false|C4684764|SAFE-Biopharma Standard|safe
Event|Event|SIMPLE_SEGMENT|6363,6372|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|6363,6372|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6363,6372|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6363,6372|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6363,6372|false|false|false|C0030685|Patient Discharge|discharge
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6363,6377|false|false|false|C0184713|Discharge to home|discharge home
Event|Event|SIMPLE_SEGMENT|6373,6377|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|6373,6377|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|6373,6377|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|6373,6377|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|6423,6433|false|false|false|||instructed
Event|Event|SIMPLE_SEGMENT|6437,6445|false|false|false|||maintain
Event|Activity|SIMPLE_SEGMENT|6455,6459|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|6455,6459|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|6455,6459|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|6455,6459|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Idea or Concept|SIMPLE_SEGMENT|6475,6479|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|6475,6479|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|6475,6479|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|6483,6487|false|false|false|||help
Event|Event|SIMPLE_SEGMENT|6488,6495|false|false|false|||prevent
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|6504,6509|false|false|false|C0000921|Accidental Falls|falls
Event|Event|SIMPLE_SEGMENT|6504,6509|false|false|false|||falls
Finding|Finding|SIMPLE_SEGMENT|6504,6509|false|false|false|C0085639|Falls|falls
Event|Event|SIMPLE_SEGMENT|6536,6545|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|6536,6545|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|6547,6555|false|false|false|||Improved
Finding|Idea or Concept|SIMPLE_SEGMENT|6567,6571|false|false|false|C1552851|next - HtmlLinkType|next
Finding|Idea or Concept|SIMPLE_SEGMENT|6572,6575|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|6572,6575|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Finding|SIMPLE_SEGMENT|6578,6584|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|6578,6584|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|SIMPLE_SEGMENT|6585,6591|false|false|false|||closer
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6595,6603|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|SIMPLE_SEGMENT|6595,6603|false|false|false|||baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|6595,6603|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Drug|Organic Chemical|SIMPLE_SEGMENT|6616,6625|false|false|false|C0017642|glipizide|Glipizide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6616,6625|false|false|false|C0017642|glipizide|Glipizide
Event|Event|SIMPLE_SEGMENT|6616,6625|false|false|false|||Glipizide
Drug|Organic Chemical|SIMPLE_SEGMENT|6630,6635|false|false|false|C0875954|Actos|actos
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6630,6635|false|false|false|C0875954|Actos|actos
Event|Event|SIMPLE_SEGMENT|6630,6635|false|false|false|||actos
Event|Event|SIMPLE_SEGMENT|6636,6640|false|false|false|||held
Finding|Idea or Concept|SIMPLE_SEGMENT|6650,6658|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|SIMPLE_SEGMENT|6660,6667|false|false|false|||Covered
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6677,6684|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|6677,6684|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6677,6684|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|6677,6684|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|6677,6684|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6677,6684|false|false|false|C0202098|Insulin measurement|insulin
Event|Event|SIMPLE_SEGMENT|6685,6692|false|false|false|||sliding
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6693,6698|false|false|false|C0222045|Integumentary scale|scale
Event|Activity|SIMPLE_SEGMENT|6693,6698|false|false|false|C1947916|Scaling|scale
Event|Event|SIMPLE_SEGMENT|6693,6698|false|false|false|||scale
Finding|Conceptual Entity|SIMPLE_SEGMENT|6693,6698|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Finding|Intellectual Product|SIMPLE_SEGMENT|6693,6698|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6703,6707|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6703,6707|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|6703,6707|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|6703,6707|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6708,6719|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6708,6719|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|6708,6719|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|6708,6719|false|false|false|C4284232|Medications|medications
Event|Event|SIMPLE_SEGMENT|6720,6729|false|false|false|||restarted
Event|Event|SIMPLE_SEGMENT|6734,6743|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|6734,6743|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6734,6743|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6734,6743|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6734,6743|false|false|false|C0030685|Patient Discharge|discharge
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6750,6753|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|6750,6753|false|false|false|||HTN
Event|Event|SIMPLE_SEGMENT|6755,6764|false|false|false|||Continued
Drug|Organic Chemical|SIMPLE_SEGMENT|6765,6775|false|false|false|C0022251|isosorbide|isosorbide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6765,6775|false|false|false|C0022251|isosorbide|isosorbide
Event|Event|SIMPLE_SEGMENT|6765,6775|false|false|false|||isosorbide
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6780,6790|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6780,6790|false|false|false|C0065374|lisinopril|lisinopril
Event|Event|SIMPLE_SEGMENT|6780,6790|false|false|false|||lisinopril
Event|Event|SIMPLE_SEGMENT|6792,6796|false|false|false|||held
Finding|Idea or Concept|SIMPLE_SEGMENT|6805,6808|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|6805,6808|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|SIMPLE_SEGMENT|6821,6831|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6821,6831|false|false|false|C0025859|metoprolol|Metoprolol
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6821,6836|false|false|false|C4082236||Metoprolol dose
Event|Event|SIMPLE_SEGMENT|6832,6836|false|false|false|||dose
Event|Event|SIMPLE_SEGMENT|6841,6848|false|false|false|||lowered
Event|Event|SIMPLE_SEGMENT|6857,6860|false|false|false|||TID
Event|Event|SIMPLE_SEGMENT|6872,6883|false|false|false|||bradycardia
Finding|Finding|SIMPLE_SEGMENT|6872,6883|false|false|false|C0428977;C3812171|Bradycardia;Bradycardia by ECG Finding|bradycardia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6888,6892|false|false|false|C0004238|Atrial Fibrillation|Afib
Event|Event|SIMPLE_SEGMENT|6888,6892|false|false|false|||Afib
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6888,6892|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Afib
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6894,6897|false|false|false|C0368980|Coagulation tissue factor induced.INR|INR
Event|Event|SIMPLE_SEGMENT|6894,6897|false|false|false|||INR
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6894,6897|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6894,6897|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Event|Event|SIMPLE_SEGMENT|6909,6918|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|6909,6918|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|6924,6931|false|false|false|||unclear
Event|Event|SIMPLE_SEGMENT|6942,6947|false|false|false|||taken
Drug|Organic Chemical|SIMPLE_SEGMENT|6959,6967|false|false|false|C0699129|Coumadin|coumadin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6959,6967|false|false|false|C0699129|Coumadin|coumadin
Event|Event|SIMPLE_SEGMENT|6968,6972|false|false|false|||dose
Event|Event|SIMPLE_SEGMENT|6981,6990|false|false|false|||restarted
Event|Event|SIMPLE_SEGMENT|7017,7022|false|false|false|||noted
Event|Event|SIMPLE_SEGMENT|7040,7048|false|false|false|||switched
Event|Event|SIMPLE_SEGMENT|7052,7061|false|false|false|||alternate
Event|Event|SIMPLE_SEGMENT|7089,7099|false|false|false|||discharged
Finding|Idea or Concept|SIMPLE_SEGMENT|7105,7109|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|7105,7109|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|7105,7109|false|false|false|C1553498|home health encounter|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|7105,7118|false|false|false|C0020043|Home visit (procedure)|home services
Event|Event|SIMPLE_SEGMENT|7110,7118|false|false|false|||services
Event|Occupational Activity|SIMPLE_SEGMENT|7110,7118|false|false|false|C0557854|Services|services
Procedure|Health Care Activity|SIMPLE_SEGMENT|7110,7118|false|false|false|C1704289|Clinical Service|services
Event|Event|SIMPLE_SEGMENT|7122,7128|false|false|false|||follow
Event|Event|SIMPLE_SEGMENT|7129,7133|false|false|false|||INRs
Finding|Idea or Concept|SIMPLE_SEGMENT|7136,7148|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Event|Event|SIMPLE_SEGMENT|7149,7155|false|false|false|||ISSUES
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7157,7162|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Event|Event|SIMPLE_SEGMENT|7157,7162|false|false|false|||Blood
Finding|Body Substance|SIMPLE_SEGMENT|7157,7162|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7157,7170|false|false|false|C0200949|Blood culture|Blood culture
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7163,7170|false|false|false|C1706355|Culture Dose Form|culture
Event|Event|SIMPLE_SEGMENT|7163,7170|false|false|false|||culture
Finding|Functional Concept|SIMPLE_SEGMENT|7163,7170|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Finding|Idea or Concept|SIMPLE_SEGMENT|7163,7170|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7163,7170|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|culture
Event|Event|SIMPLE_SEGMENT|7179,7184|false|false|false|||needs
Event|Event|SIMPLE_SEGMENT|7191,7197|false|false|false|||follow
Event|Event|SIMPLE_SEGMENT|7206,7212|false|false|false|||growth
Finding|Finding|SIMPLE_SEGMENT|7206,7212|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|7206,7212|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Finding|Organism Function|SIMPLE_SEGMENT|7206,7212|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Finding|Physiologic Function|SIMPLE_SEGMENT|7206,7212|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|7206,7212|true|false|false|C2911660|Growth action|growth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7225,7236|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7225,7236|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|7225,7236|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|7225,7236|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|7225,7249|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|SIMPLE_SEGMENT|7240,7249|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|7240,7249|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Organic Chemical|SIMPLE_SEGMENT|7252,7263|false|false|false|C0002144|allopurinol|Allopurinol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7252,7263|false|false|false|C0002144|allopurinol|Allopurinol
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7279,7285|false|false|false|C0039225|Tablet Dosage Form|TABLET
Event|Event|SIMPLE_SEGMENT|7286,7290|false|false|false|||Take
Drug|Organic Chemical|SIMPLE_SEGMENT|7307,7321|false|false|false|C0042845;C3714801|Cyanocobalamin Drug Class;vitamin B12|Cyanocobalamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7307,7321|false|false|false|C0042845;C3714801|Cyanocobalamin Drug Class;vitamin B12|Cyanocobalamin
Drug|Vitamin|SIMPLE_SEGMENT|7307,7321|false|false|false|C0042845;C3714801|Cyanocobalamin Drug Class;vitamin B12|Cyanocobalamin
Event|Event|SIMPLE_SEGMENT|7327,7330|false|false|false|||MCG
Event|Event|SIMPLE_SEGMENT|7348,7352|false|false|false|||Take
Procedure|Health Care Activity|SIMPLE_SEGMENT|7348,7352|false|false|false|C1515187|Take|Take
Drug|Organic Chemical|SIMPLE_SEGMENT|7377,7390|false|false|false|C0011777|dexamethasone|Dexamethasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7377,7390|false|false|false|C0011777|dexamethasone|Dexamethasone
Event|Event|SIMPLE_SEGMENT|7377,7390|false|false|false|||Dexamethasone
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7406,7412|false|false|false|C0039225|Tablet Dosage Form|TABLET
Event|Event|SIMPLE_SEGMENT|7406,7412|false|false|false|||TABLET
Event|Event|SIMPLE_SEGMENT|7413,7417|false|false|false|||Take
Drug|Organic Chemical|SIMPLE_SEGMENT|7434,7443|false|false|false|C0017642|glipizide|Glipizide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7434,7443|false|false|false|C0017642|glipizide|Glipizide
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7457,7463|false|false|false|C0039225|Tablet Dosage Form|TABLET
Event|Event|SIMPLE_SEGMENT|7457,7463|false|false|false|||TABLET
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7475,7478|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7475,7478|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7475,7478|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|7475,7478|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|7475,7478|false|false|false|C1332410|BID gene|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7486,7495|false|false|false|C0120107|goserelin|Goserelin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7486,7495|false|false|false|C0120107|goserelin|Goserelin
Event|Event|SIMPLE_SEGMENT|7486,7495|false|false|false|||Goserelin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7486,7503|false|false|false|C0700476|goserelin acetate|Goserelin acetate
Drug|Hormone|SIMPLE_SEGMENT|7486,7503|false|false|false|C0700476|goserelin acetate|Goserelin acetate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7486,7503|false|false|false|C0700476|goserelin acetate|Goserelin acetate
Drug|Organic Chemical|SIMPLE_SEGMENT|7496,7503|false|false|false|C0000975|acetate|acetate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7496,7503|false|false|false|C0000975|acetate|acetate
Event|Event|SIMPLE_SEGMENT|7496,7503|false|false|false|||acetate
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7520,7527|false|false|false|C5444783||IMPLANT
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|7520,7527|false|false|false|C0332837|Traumatic implant|IMPLANT
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7520,7527|false|false|false|C1704229|Drug Implant|IMPLANT
Event|Event|SIMPLE_SEGMENT|7520,7527|false|false|false|||IMPLANT
Finding|Functional Concept|SIMPLE_SEGMENT|7520,7527|false|false|false|C1546675;C1711357|Administration via Implantation|IMPLANT
Finding|Intellectual Product|SIMPLE_SEGMENT|7520,7527|false|false|false|C1546675;C1711357|Administration via Implantation|IMPLANT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7520,7527|false|false|false|C0021107|Implantation procedure|IMPLANT
Event|Event|SIMPLE_SEGMENT|7539,7545|false|false|false|||QMONTH
Drug|Organic Chemical|SIMPLE_SEGMENT|7554,7564|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7554,7564|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|SIMPLE_SEGMENT|7554,7574|false|false|false|C0022252|isosorbide dinitrate|Isosorbide dinitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7554,7574|false|false|false|C0022252|isosorbide dinitrate|Isosorbide dinitrate
Event|Event|SIMPLE_SEGMENT|7565,7574|false|false|false|||dinitrate
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7588,7594|false|false|false|C0039225|Tablet Dosage Form|TABLET
Event|Event|SIMPLE_SEGMENT|7588,7594|false|false|false|||TABLET
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7606,7609|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7606,7609|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7606,7609|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|7606,7609|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|7606,7609|false|false|false|C1332410|BID gene|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7618,7628|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7618,7628|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7642,7648|false|false|false|C0039225|Tablet Dosage Form|TABLET
Event|Event|SIMPLE_SEGMENT|7649,7653|false|false|false|||Take
Drug|Organic Chemical|SIMPLE_SEGMENT|7670,7679|false|false|false|C0025242|memantine|Memantine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7670,7679|false|false|false|C0025242|memantine|Memantine
Drug|Organic Chemical|SIMPLE_SEGMENT|7690,7700|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7690,7700|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|7690,7709|false|false|false|C0700548|metoprolol tartrate|Metoprolol tartrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7690,7709|false|false|false|C0700548|metoprolol tartrate|Metoprolol tartrate
Drug|Organic Chemical|SIMPLE_SEGMENT|7701,7709|false|false|false|C0039328;C0144544|Tartrates;tartrate|tartrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7701,7709|false|false|false|C0039328;C0144544|Tartrates;tartrate|tartrate
Event|Event|SIMPLE_SEGMENT|7701,7709|false|false|false|||tartrate
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7723,7729|false|false|false|C0039225|Tablet Dosage Form|TABLET
Event|Event|SIMPLE_SEGMENT|7730,7734|false|false|false|||Take
Event|Event|SIMPLE_SEGMENT|7741,7744|false|false|false|||TID
Drug|Organic Chemical|SIMPLE_SEGMENT|7753,7763|false|false|false|C0068771|nilutamide|Nilutamide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7753,7763|false|false|false|C0068771|nilutamide|Nilutamide
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7779,7785|false|false|false|C0039225|Tablet Dosage Form|TABLET
Event|Event|SIMPLE_SEGMENT|7779,7785|false|false|false|||TABLET
Drug|Organic Chemical|SIMPLE_SEGMENT|7807,7820|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7807,7820|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Organic Chemical|SIMPLE_SEGMENT|7831,7840|false|false|false|C0030049|oxycodone|Oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7831,7840|false|false|false|C0030049|oxycodone|Oxycodone
Event|Event|SIMPLE_SEGMENT|7831,7840|false|false|false|||Oxycodone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7831,7840|false|false|false|C0524222|Oxycodone measurement|Oxycodone
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7851,7857|false|false|false|C0039225|Tablet Dosage Form|TABLET
Event|Event|SIMPLE_SEGMENT|7858,7862|false|false|false|||Take
Procedure|Health Care Activity|SIMPLE_SEGMENT|7858,7862|false|false|false|C1515187|Take|Take
Finding|Gene or Genome|SIMPLE_SEGMENT|7873,7876|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7877,7881|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|7877,7881|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|7877,7881|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|7877,7881|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Hormone|SIMPLE_SEGMENT|7889,7899|false|false|false|C0032952|prednisone|Prednisone
Drug|Organic Chemical|SIMPLE_SEGMENT|7889,7899|false|false|false|C0032952|prednisone|Prednisone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7889,7899|false|false|false|C0032952|prednisone|Prednisone
Event|Event|SIMPLE_SEGMENT|7900,7905|false|false|false|||Taper
Procedure|Health Care Activity|SIMPLE_SEGMENT|7900,7905|false|false|false|C0441640||Taper
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7913,7919|false|false|false|C0039225|Tablet Dosage Form|TABLET
Event|Event|SIMPLE_SEGMENT|7913,7919|false|false|false|||TABLET
Event|Event|SIMPLE_SEGMENT|7928,7930|false|false|false|||PO
Drug|Organic Chemical|SIMPLE_SEGMENT|7948,7959|false|false|false|C0074554|simvastatin|Simvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7948,7959|false|false|false|C0074554|simvastatin|Simvastatin
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7973,7979|false|false|false|C0039225|Tablet Dosage Form|TABLET
Event|Event|SIMPLE_SEGMENT|7980,7984|false|false|false|||Take
Event|Event|SIMPLE_SEGMENT|7991,7994|false|false|false|||QPM
Drug|Organic Chemical|SIMPLE_SEGMENT|8002,8011|false|false|false|C0076840|torsemide|Torsemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8002,8011|false|false|false|C0076840|torsemide|Torsemide
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8023,8029|false|false|false|C0039225|Tablet Dosage Form|TABLET
Event|Event|SIMPLE_SEGMENT|8030,8034|false|false|false|||Take
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|8051,8059|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|SIMPLE_SEGMENT|8051,8059|false|false|false|C0043031|warfarin|Warfarin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8051,8059|false|false|false|C0043031|warfarin|Warfarin
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|8051,8066|false|false|false|C0376218|warfarin sodium|Warfarin sodium
Drug|Organic Chemical|SIMPLE_SEGMENT|8051,8066|false|false|false|C0376218|warfarin sodium|Warfarin sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8051,8066|false|false|false|C0376218|warfarin sodium|Warfarin sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8060,8066|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|8060,8066|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8060,8066|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Event|Event|SIMPLE_SEGMENT|8060,8066|false|false|false|||sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|8060,8066|false|false|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8060,8066|false|false|false|C0337443|Sodium measurement|sodium
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8082,8088|false|false|false|C0039225|Tablet Dosage Form|TABLET
Event|Event|SIMPLE_SEGMENT|8082,8088|false|false|false|||TABLET
Event|Event|SIMPLE_SEGMENT|8089,8093|false|false|false|||Take
Event|Event|SIMPLE_SEGMENT|8097,8099|false|false|false|||PO
Event|Event|SIMPLE_SEGMENT|8103,8111|false|false|false|||directed
Event|Event|SIMPLE_SEGMENT|8117,8126|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|8117,8126|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8117,8126|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8117,8126|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8117,8126|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|8117,8138|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8127,8138|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8127,8138|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|8127,8138|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|8127,8138|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|8143,8156|false|false|false|C0011777|dexamethasone|dexamethasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8143,8156|false|false|false|C0011777|dexamethasone|dexamethasone
Event|Event|SIMPLE_SEGMENT|8143,8156|false|false|false|||dexamethasone
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8164,8170|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|8171,8174|false|false|false|||Sig
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8184,8190|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Intellectual Product|SIMPLE_SEGMENT|8194,8198|false|false|false|C1720092|Once - dosing instruction fragment|once
Finding|Idea or Concept|SIMPLE_SEGMENT|8202,8205|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|8202,8205|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|SIMPLE_SEGMENT|8212,8221|false|false|false|C0017642|glipizide|glipizide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8212,8221|false|false|false|C0017642|glipizide|glipizide
Event|Event|SIMPLE_SEGMENT|8212,8221|false|false|false|||glipizide
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8228,8234|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8248,8254|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|8248,8254|false|false|false|||Tablet
Event|Event|SIMPLE_SEGMENT|8255,8257|false|false|false|||PO
Finding|Intellectual Product|SIMPLE_SEGMENT|8258,8262|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8258,8268|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|SIMPLE_SEGMENT|8265,8268|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|8265,8268|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8275,8284|false|false|false|C0120107|goserelin|goserelin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8275,8284|false|false|false|C0120107|goserelin|goserelin
Event|Event|SIMPLE_SEGMENT|8275,8284|false|false|false|||goserelin
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8293,8300|false|false|false|C5444783||Implant
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|8293,8300|false|false|false|C0332837|Traumatic implant|Implant
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8293,8300|false|false|false|C1704229|Drug Implant|Implant
Event|Event|SIMPLE_SEGMENT|8293,8300|false|false|false|||Implant
Finding|Functional Concept|SIMPLE_SEGMENT|8293,8300|false|false|false|C1546675;C1711357|Administration via Implantation|Implant
Finding|Intellectual Product|SIMPLE_SEGMENT|8293,8300|false|false|false|C1546675;C1711357|Administration via Implantation|Implant
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8293,8300|false|false|false|C0021107|Implantation procedure|Implant
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8314,8321|false|false|false|C5444783||implant
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|8314,8321|false|false|false|C0332837|Traumatic implant|implant
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8314,8321|false|false|false|C1704229|Drug Implant|implant
Event|Event|SIMPLE_SEGMENT|8314,8321|false|false|false|||implant
Finding|Functional Concept|SIMPLE_SEGMENT|8314,8321|false|false|false|C1546675;C1711357|Administration via Implantation|implant
Finding|Intellectual Product|SIMPLE_SEGMENT|8314,8321|false|false|false|C1546675;C1711357|Administration via Implantation|implant
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8314,8321|false|false|false|C0021107|Implantation procedure|implant
Event|Event|SIMPLE_SEGMENT|8322,8334|false|false|false|||Subcutaneous
Finding|Functional Concept|SIMPLE_SEGMENT|8322,8334|false|false|false|C1522438|Subcutaneous Route of Administration|Subcutaneous
Event|Event|SIMPLE_SEGMENT|8339,8347|false|false|false|||directed
Drug|Organic Chemical|SIMPLE_SEGMENT|8354,8364|false|false|false|C0022251|isosorbide|isosorbide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8354,8364|false|false|false|C0022251|isosorbide|isosorbide
Event|Event|SIMPLE_SEGMENT|8354,8364|false|false|false|||isosorbide
Drug|Organic Chemical|SIMPLE_SEGMENT|8354,8374|false|false|false|C0022252|isosorbide dinitrate|isosorbide dinitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8354,8374|false|false|false|C0022252|isosorbide dinitrate|isosorbide dinitrate
Event|Event|SIMPLE_SEGMENT|8365,8374|false|false|false|||dinitrate
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8381,8387|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8401,8407|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|SIMPLE_SEGMENT|8420,8423|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|8420,8423|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8430,8440|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8430,8440|false|false|false|C0065374|lisinopril|lisinopril
Event|Event|SIMPLE_SEGMENT|8430,8440|false|false|false|||lisinopril
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8447,8453|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8467,8473|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|8467,8473|false|false|false|||Tablet
Event|Event|SIMPLE_SEGMENT|8474,8476|false|false|false|||PO
Finding|Intellectual Product|SIMPLE_SEGMENT|8477,8481|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8477,8487|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|SIMPLE_SEGMENT|8484,8487|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|8484,8487|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|SIMPLE_SEGMENT|8494,8504|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8494,8504|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|SIMPLE_SEGMENT|8494,8504|false|false|false|||metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|8494,8513|false|false|false|C0700548|metoprolol tartrate|metoprolol tartrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8494,8513|false|false|false|C0700548|metoprolol tartrate|metoprolol tartrate
Drug|Organic Chemical|SIMPLE_SEGMENT|8505,8513|false|false|false|C0039328;C0144544|Tartrates;tartrate|tartrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8505,8513|false|false|false|C0039328;C0144544|Tartrates;tartrate|tartrate
Event|Event|SIMPLE_SEGMENT|8505,8513|false|false|false|||tartrate
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8520,8526|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8540,8546|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|8540,8546|false|false|false|||Tablet
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8557,8562|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Event|Event|SIMPLE_SEGMENT|8557,8562|false|false|false|||times
Finding|Idea or Concept|SIMPLE_SEGMENT|8565,8568|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|8565,8568|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8579,8585|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|SIMPLE_SEGMENT|8590,8597|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|8605,8615|false|false|false|C0068771|nilutamide|nilutamide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8605,8615|false|false|false|C0068771|nilutamide|nilutamide
Event|Event|SIMPLE_SEGMENT|8605,8615|false|false|false|||nilutamide
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8623,8629|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8643,8649|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|8643,8649|false|false|false|||Tablet
Event|Event|SIMPLE_SEGMENT|8650,8652|false|false|false|||PO
Finding|Intellectual Product|SIMPLE_SEGMENT|8653,8657|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8653,8663|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|SIMPLE_SEGMENT|8660,8663|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|8660,8663|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|SIMPLE_SEGMENT|8670,8679|false|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8670,8679|false|false|false|C0030049|oxycodone|oxycodone
Event|Event|SIMPLE_SEGMENT|8670,8679|false|false|false|||oxycodone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8670,8679|false|false|false|C0524222|Oxycodone measurement|oxycodone
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8685,8691|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8705,8711|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|8739,8745|false|false|false|||needed
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8750,8754|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|8750,8754|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|8750,8754|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|8750,8754|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|8761,8772|false|false|false|C0074554|simvastatin|simvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8761,8772|false|false|false|C0074554|simvastatin|simvastatin
Event|Event|SIMPLE_SEGMENT|8761,8772|false|false|false|||simvastatin
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8779,8785|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8795,8801|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|8795,8801|false|false|false|||Tablet
Drug|Organic Chemical|SIMPLE_SEGMENT|8826,8835|false|false|false|C0076840|torsemide|torsemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8826,8835|false|false|false|C0076840|torsemide|torsemide
Event|Event|SIMPLE_SEGMENT|8826,8835|false|false|false|||torsemide
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8842,8848|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8862,8868|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|8862,8868|false|false|false|||Tablet
Event|Event|SIMPLE_SEGMENT|8869,8871|false|false|false|||PO
Finding|Intellectual Product|SIMPLE_SEGMENT|8872,8876|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8872,8882|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|SIMPLE_SEGMENT|8879,8882|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|8879,8882|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8893,8899|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|SIMPLE_SEGMENT|8904,8911|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|8920,8934|false|false|false|C0042845;C3714801|Cyanocobalamin Drug Class;vitamin B12|cyanocobalamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8920,8934|false|false|false|C0042845;C3714801|Cyanocobalamin Drug Class;vitamin B12|cyanocobalamin
Drug|Vitamin|SIMPLE_SEGMENT|8920,8934|false|false|false|C0042845;C3714801|Cyanocobalamin Drug Class;vitamin B12|cyanocobalamin
Event|Event|SIMPLE_SEGMENT|8920,8934|false|false|false|||cyanocobalamin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8920,8949|false|false|false|C0202252|VITAMIN B12 MEASUREMENT|cyanocobalamin (vitamin B-12)
Drug|Organic Chemical|SIMPLE_SEGMENT|8936,8943|false|false|false|C0042890|Vitamins|vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8936,8943|false|false|false|C0042890|Vitamins|vitamin
Drug|Vitamin|SIMPLE_SEGMENT|8936,8943|false|false|false|C0042890|Vitamins|vitamin
Drug|Organic Chemical|SIMPLE_SEGMENT|8936,8945|false|false|false|C0042849;C1704763;C5442122|B Vitamin Family;VITAMIN B;vitamin B complex|vitamin B
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8936,8945|false|false|false|C0042849;C1704763;C5442122|B Vitamin Family;VITAMIN B;vitamin B complex|vitamin B
Drug|Vitamin|SIMPLE_SEGMENT|8936,8945|false|false|false|C0042849;C1704763;C5442122|B Vitamin Family;VITAMIN B;vitamin B complex|vitamin B
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|8936,8948|false|false|false|C0042845;C0086024|cobalamins;vitamin B12|vitamin B-12
Drug|Organic Chemical|SIMPLE_SEGMENT|8936,8948|false|false|false|C0042845;C0086024|cobalamins;vitamin B12|vitamin B-12
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8936,8948|false|false|false|C0042845;C0086024|cobalamins;vitamin B12|vitamin B-12
Drug|Vitamin|SIMPLE_SEGMENT|8936,8948|false|false|false|C0042845;C0086024|cobalamins;vitamin B12|vitamin B-12
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8936,8948|false|false|false|C0202252|VITAMIN B12 MEASUREMENT|vitamin B-12
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8966,8972|false|false|false|C0302908;C1697794|Liquid Dosage Form;Liquid substance|Liquid
Drug|Substance|SIMPLE_SEGMENT|8966,8972|false|false|false|C0302908;C1697794|Liquid Dosage Form;Liquid substance|Liquid
Event|Event|SIMPLE_SEGMENT|8966,8972|false|false|false|||Liquid
Finding|Finding|SIMPLE_SEGMENT|8966,8972|false|false|false|C1304698|Liquid (finding)|Liquid
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8966,8972|false|false|false|C0301571|Liquid diet|Liquid
Finding|Intellectual Product|SIMPLE_SEGMENT|8995,8999|false|false|false|C1720092|Once - dosing instruction fragment|once
Finding|Intellectual Product|SIMPLE_SEGMENT|9002,9006|false|false|false|C1561540|Transaction counts and value totals - week|week
Drug|Organic Chemical|SIMPLE_SEGMENT|9014,9023|false|false|false|C0025242|memantine|memantine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9014,9023|false|false|false|C0025242|memantine|memantine
Event|Event|SIMPLE_SEGMENT|9014,9023|false|false|false|||memantine
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9030,9036|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9050,9056|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|SIMPLE_SEGMENT|9068,9071|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|9068,9071|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|SIMPLE_SEGMENT|9079,9090|false|false|false|C0002144|allopurinol|allopurinol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9079,9090|false|false|false|C0002144|allopurinol|allopurinol
Event|Event|SIMPLE_SEGMENT|9079,9090|false|false|false|||allopurinol
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9098,9104|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9118,9124|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|9125,9127|false|false|false|||PO
Finding|Intellectual Product|SIMPLE_SEGMENT|9128,9132|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9128,9138|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|SIMPLE_SEGMENT|9135,9138|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|9135,9138|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|9147,9155|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|SIMPLE_SEGMENT|9147,9155|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9147,9155|false|false|false|C0043031|warfarin|warfarin
Event|Event|SIMPLE_SEGMENT|9147,9155|false|false|false|||warfarin
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9163,9169|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|9170,9173|false|false|false|||Sig
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9183,9189|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9215,9222|false|false|false|C0039225|Tablet Dosage Form|tablets
Event|Event|SIMPLE_SEGMENT|9215,9222|false|false|false|||tablets
Drug|Organic Chemical|SIMPLE_SEGMENT|9252,9259|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9252,9259|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|SIMPLE_SEGMENT|9252,9259|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|SIMPLE_SEGMENT|9252,9261|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|SIMPLE_SEGMENT|9252,9261|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9252,9261|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|SIMPLE_SEGMENT|9252,9261|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9252,9261|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9273,9279|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|9273,9279|false|false|false|||Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9293,9299|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Intellectual Product|SIMPLE_SEGMENT|9303,9307|false|false|false|C1720092|Once - dosing instruction fragment|once
Finding|Idea or Concept|SIMPLE_SEGMENT|9311,9314|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|9311,9314|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9322,9329|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|9322,9329|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9322,9329|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|9322,9329|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|9322,9329|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9322,9329|false|false|false|C0202098|Insulin measurement|insulin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9322,9338|false|false|false|C0907402|insulin glargine|insulin glargine
Drug|Hormone|SIMPLE_SEGMENT|9322,9338|false|false|false|C0907402|insulin glargine|insulin glargine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9322,9338|false|false|false|C0907402|insulin glargine|insulin glargine
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9330,9338|false|false|false|C0907402|insulin glargine|glargine
Drug|Hormone|SIMPLE_SEGMENT|9330,9338|false|false|false|C0907402|insulin glargine|glargine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9330,9338|false|false|false|C0907402|insulin glargine|glargine
Event|Event|SIMPLE_SEGMENT|9330,9338|false|false|false|||glargine
Event|Event|SIMPLE_SEGMENT|9351,9360|false|false|false|||Cartridge
Finding|Intellectual Product|SIMPLE_SEGMENT|9351,9360|false|false|false|C1553461|Cartridge - package type|Cartridge
Event|Event|SIMPLE_SEGMENT|9382,9394|false|false|false|||Subcutaneous
Finding|Functional Concept|SIMPLE_SEGMENT|9382,9394|false|false|false|C1522438|Subcutaneous Route of Administration|Subcutaneous
Event|Event|SIMPLE_SEGMENT|9412,9421|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|9412,9421|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|9412,9421|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|9412,9421|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|9412,9421|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9412,9433|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|9412,9433|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9422,9433|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|9422,9433|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|9422,9433|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|SIMPLE_SEGMENT|9435,9439|false|false|false|||Home
Finding|Idea or Concept|SIMPLE_SEGMENT|9435,9439|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|9435,9439|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|9435,9439|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|SIMPLE_SEGMENT|9445,9452|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|9445,9452|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|SIMPLE_SEGMENT|9455,9463|false|false|false|||Facility
Finding|Intellectual Product|SIMPLE_SEGMENT|9455,9463|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|SIMPLE_SEGMENT|9471,9480|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|9471,9480|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|9471,9480|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|9471,9480|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|9471,9480|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|9471,9490|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9481,9490|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|9481,9490|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|9481,9490|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|9481,9490|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9481,9490|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Intellectual Product|SIMPLE_SEGMENT|9500,9505|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9500,9551|false|false|false|C2732749|Acute on chronic diastolic heart failure|Acute on chronic diastolic congestive heart failure
Finding|Intellectual Product|SIMPLE_SEGMENT|9509,9516|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|9509,9516|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9509,9551|false|false|false|C2711480|Chronic diastolic heart failure|chronic diastolic congestive heart failure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9517,9526|false|false|false|C0012000|Diastole|diastolic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9517,9551|false|false|false|C2183328|diastolic congestive heart failure|diastolic congestive heart failure
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9527,9551|false|false|false|C0018802|Congestive heart failure|congestive heart failure
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9538,9543|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|9538,9543|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|9538,9543|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9538,9551|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Event|Event|SIMPLE_SEGMENT|9544,9551|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|9544,9551|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|9544,9551|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|9544,9551|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Disorder|Neoplastic Process|SIMPLE_SEGMENT|9553,9562|false|false|false|C0027627|Neoplasm Metastasis|SECONDARY
Event|Event|SIMPLE_SEGMENT|9553,9562|false|false|false|||SECONDARY
Finding|Functional Concept|SIMPLE_SEGMENT|9553,9562|false|false|false|C1522484|metastatic qualifier|SECONDARY
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9563,9569|false|false|false|C0018792|Heart Atrium|Atrial
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9563,9582|false|false|false|C2926591||Atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9563,9582|false|false|false|C0004238|Atrial Fibrillation|Atrial fibrillation
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|9563,9582|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9570,9582|false|false|false|C0232197|Fibrillation|fibrillation
Event|Event|SIMPLE_SEGMENT|9570,9582|false|false|false|||fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9583,9591|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|Diabetes
Event|Event|SIMPLE_SEGMENT|9583,9591|false|false|false|||Diabetes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9592,9604|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|SIMPLE_SEGMENT|9592,9604|false|false|false|||Hypertension
Event|Event|SIMPLE_SEGMENT|9607,9616|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|9607,9616|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|9607,9616|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|9607,9616|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|9607,9616|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9617,9626|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9617,9626|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|9617,9626|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|9617,9626|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|9628,9634|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9628,9641|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|9628,9641|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9635,9641|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|9635,9641|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|9643,9648|false|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|9643,9648|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|9653,9661|false|false|false|||coherent
Finding|Finding|SIMPLE_SEGMENT|9653,9661|false|false|false|C4068804|Coherent|coherent
Event|Event|SIMPLE_SEGMENT|9663,9668|false|false|false|||Level
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9663,9685|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|9663,9685|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|SIMPLE_SEGMENT|9672,9685|false|false|false|||Consciousness
Finding|Finding|SIMPLE_SEGMENT|9672,9685|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|9672,9685|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9687,9692|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|9687,9692|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9687,9692|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|9687,9692|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|9687,9692|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|9687,9692|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|9687,9692|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|9697,9708|false|false|false|||interactive
Finding|Functional Concept|SIMPLE_SEGMENT|9697,9708|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|9710,9718|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|9710,9718|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|9710,9718|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9719,9725|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|9719,9725|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|9719,9725|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|SIMPLE_SEGMENT|9727,9737|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|9727,9737|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|9727,9737|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|9727,9737|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|SIMPLE_SEGMENT|9740,9748|false|false|false|||requires
Event|Event|SIMPLE_SEGMENT|9749,9759|false|false|false|||assistance
Finding|Social Behavior|SIMPLE_SEGMENT|9749,9759|false|false|false|C0018896|Helping Behavior|assistance
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9763,9766|false|false|false|C1454018|AICDA protein, human|aid
Drug|Enzyme|SIMPLE_SEGMENT|9763,9766|false|false|false|C1454018|AICDA protein, human|aid
Event|Event|SIMPLE_SEGMENT|9763,9766|false|false|false|||aid
Finding|Gene or Genome|SIMPLE_SEGMENT|9763,9766|false|false|false|C1421876;C3540469|AICDA gene;AICDA wt Allele|aid
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9763,9766|false|false|false|C0021588;C0280108|AID - Artificial insemination by donor;dacarbazine/doxorubicin/ifosfamide protocol|aid
Event|Event|SIMPLE_SEGMENT|9768,9774|false|false|false|||walker
Event|Event|SIMPLE_SEGMENT|9788,9797|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|9788,9797|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|9788,9797|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|9788,9797|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|9788,9797|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9788,9810|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|9788,9810|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|9788,9810|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9798,9810|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|9798,9810|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|9798,9810|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Event|Event|SIMPLE_SEGMENT|9832,9840|false|false|false|||admitted
Finding|Idea or Concept|SIMPLE_SEGMENT|9848,9856|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|SIMPLE_SEGMENT|9861,9869|false|false|false|||swelling
Finding|Finding|SIMPLE_SEGMENT|9861,9869|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|9861,9869|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9878,9882|false|false|false|C1140621|Leg|legs
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9878,9882|false|false|false|C5781420||legs
Finding|Finding|SIMPLE_SEGMENT|9885,9891|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|9885,9891|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9904,9909|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|9904,9909|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|9904,9909|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9904,9917|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Event|Event|SIMPLE_SEGMENT|9910,9917|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|9910,9917|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|9910,9917|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|9910,9917|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|SIMPLE_SEGMENT|9922,9931|false|false|false|||increased
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9937,9945|false|false|false|C0012798;C5399719|Diuretic [APC];Diuretics|diuretic
Event|Event|SIMPLE_SEGMENT|9937,9945|false|false|false|||diuretic
Event|Event|SIMPLE_SEGMENT|9966,9970|false|false|false|||work
Finding|Finding|SIMPLE_SEGMENT|9976,9984|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Finding|Functional Concept|SIMPLE_SEGMENT|9976,9984|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|9976,9984|false|false|false|C0031809|Physical Examination|physical
Finding|Intellectual Product|SIMPLE_SEGMENT|9976,9992|false|false|false|C1547999|Diagnostic Service Section ID - Physical Therapy|physical therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9976,9992|false|false|false|C0949766|Physical therapy|physical therapy
Event|Event|SIMPLE_SEGMENT|9985,9992|false|false|false|||therapy
Finding|Finding|SIMPLE_SEGMENT|9985,9992|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|SIMPLE_SEGMENT|9985,9992|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9985,9992|false|false|false|C0087111|Therapeutic procedure|therapy
Event|Event|SIMPLE_SEGMENT|10002,10007|false|false|false|||weigh
Event|Event|SIMPLE_SEGMENT|10039,10045|false|false|false|||doctor
Finding|Intellectual Product|SIMPLE_SEGMENT|10039,10045|false|false|false|C2348314|Doctor - Title|doctor
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10055,10061|false|false|false|C0944911||weight
Event|Event|SIMPLE_SEGMENT|10055,10061|false|false|false|||weight
Finding|Finding|SIMPLE_SEGMENT|10055,10061|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|10055,10061|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|10055,10061|false|false|false|C1305866|Weighing patient|weight
Event|Event|SIMPLE_SEGMENT|10062,10071|false|false|false|||increases
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10095,10105|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|10095,10105|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Event|Event|SIMPLE_SEGMENT|10106,10113|false|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|10106,10113|false|false|false|C0392747|Changing|changes
Finding|Idea or Concept|SIMPLE_SEGMENT|10117,10125|false|false|false|C0549178|Continuous|CONTINUE
Drug|Organic Chemical|SIMPLE_SEGMENT|10126,10135|false|false|false|C0076840|torsemide|torsemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10126,10135|false|false|false|C0076840|torsemide|torsemide
Event|Event|SIMPLE_SEGMENT|10126,10135|false|false|false|||torsemide
Event|Event|SIMPLE_SEGMENT|10150,10154|false|false|false|||help
Event|Event|SIMPLE_SEGMENT|10155,10161|false|false|false|||remove
Drug|Substance|SIMPLE_SEGMENT|10162,10167|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|10162,10167|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|10162,10167|false|false|false|C1546638|Fluid Specimen Code|fluid
Drug|Organic Chemical|SIMPLE_SEGMENT|10177,10187|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10177,10187|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|SIMPLE_SEGMENT|10177,10187|false|false|false|||metoprolol
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10210,10215|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|10210,10215|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|10210,10215|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|SIMPLE_SEGMENT|10210,10224|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Finding|Organism Function|SIMPLE_SEGMENT|10210,10224|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Procedure|Health Care Activity|SIMPLE_SEGMENT|10210,10224|false|false|false|C0005824|Blood pressure determination|blood pressure
Event|Event|SIMPLE_SEGMENT|10216,10224|false|false|false|||pressure
Finding|Finding|SIMPLE_SEGMENT|10216,10224|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|10216,10224|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|10216,10224|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|10216,10224|false|false|false|C0033095||pressure
Event|Event|SIMPLE_SEGMENT|10235,10238|false|false|false|||low
Finding|Finding|SIMPLE_SEGMENT|10235,10238|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|SIMPLE_SEGMENT|10235,10238|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Event|Event|SIMPLE_SEGMENT|10254,10266|false|false|false|||hospitalized
Event|Event|SIMPLE_SEGMENT|10274,10280|false|false|false|||doctor
Finding|Intellectual Product|SIMPLE_SEGMENT|10274,10280|false|false|false|C2348314|Doctor - Title|doctor
Event|Event|SIMPLE_SEGMENT|10285,10291|false|false|false|||decide
Event|Event|SIMPLE_SEGMENT|10296,10304|false|false|false|||increase
Finding|Idea or Concept|SIMPLE_SEGMENT|10322,10328|false|false|false|C1549636|Address type - Office|office
Procedure|Health Care Activity|SIMPLE_SEGMENT|10322,10334|false|false|false|C0028900|Office Visits|office visit
Event|Event|SIMPLE_SEGMENT|10329,10334|false|false|false|||visit
Finding|Social Behavior|SIMPLE_SEGMENT|10329,10334|false|false|false|C0545082|Visit|visit
Procedure|Health Care Activity|SIMPLE_SEGMENT|10338,10346|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10347,10359|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|10347,10359|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|10347,10359|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

