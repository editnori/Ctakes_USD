CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|Percocet|Drug|false|false||Percocet
null|Percocet|Drug|false|false||Percocetnull|Vicodin|Drug|false|false||Vicodin
null|Vicodin|Drug|false|false||Vicodinnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Abdominal Pain|Finding|false|false||Abdominal painnull|Abdomen|Anatomy|false|false||Abdominalnull|Abdominal (qualifier value)|Modifier|false|false||Abdominalnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Paracentesis|Procedure|false|false||Paracentesisnull|HIV Vaccine|Drug|false|false||HIV
null|HIV Vaccine|Drug|false|false||HIVnull|HIV Infections|Disorder|false|false||HIV
null|HIV|Disorder|false|false||HIVnull|Antiretroviral Therapy, Highly Active|Procedure|false|false||HAARTnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|SAT1 protein, human|Drug|false|false||sat
null|SAT1 protein, human|Drug|false|false||satnull|College Entrance Examination Board Scholastic Aptitude Test|Finding|false|false||sat
null|SAT1 wt Allele|Finding|false|false||sat
null|SAT1 gene|Finding|false|false||satnull|Santali language|Entity|false|false||satnull|Legal fine|Entity|false|false||finenull|Fine (qualifier value)|Modifier|false|false||finenull|On admission|Time|false|false||on admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|hepatitis C virus|Disorder|false|false||HCV
null|Hepatitis C|Disorder|false|false||HCVnull|Liver Cirrhosis|Disorder|false|false||cirrhosis
null|Cirrhosis|Disorder|false|false||cirrhosisnull|Ascites|Disorder|false|false||ascitesnull|Peritoneal Effusion|Finding|false|false||ascitesnull|Biweekly|Time|false|false||biweeklynull|Therapeutic brand of coal tar|Drug|false|false||therapeutic
null|Therapeutic brand of coal tar|Drug|false|false||therapeuticnull|Therapeutic - Location Service Code|Finding|false|false||therapeutic
null|Therapeutic|Finding|false|false||therapeuticnull|Therapeutic procedure|Procedure|false|false||therapeuticnull|Paracentesis|Procedure|false|false||paracentesesnull|Hepatic Encephalopathy|Disorder|false|false||hepatic encephalopathynull|Hepatic|Anatomy|false|false||hepaticnull|Encephalopathies|Disorder|false|false||encephalopathynull|Transplant|Finding|false|false||transplant
null|Transplanted organ and tissue status|Finding|false|false||transplantnull|Transplantation|Procedure|false|false||transplantnull|Transplanted tissue|Anatomy|false|false||transplantnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Comorbidity|Finding|false|false||comorbiditiesnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false||abdnull|ABD (body structure)|Anatomy|false|false||abd
null|Abdomen|Anatomy|false|false||abdnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Ascites|Disorder|false|false||ascitesnull|Peritoneal Effusion|Finding|false|false||ascitesnull|Paracentesis|Procedure|false|false||paracentesisnull|Last|Modifier|false|false||lastnull|Paracentesis|Procedure|false|false||paracentesisnull|Patient Outcome - Worsening|Finding|false|false||worseningnull|Worsening (qualifier value)|Modifier|false|false||worseningnull|Abdominal Pain|Finding|false|false||abdominal painnull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Constant - dosing instruction fragment|Finding|false|false||constantnull|Constant (qualifier)|Modifier|false|false||constantnull|Epigastric|Anatomy|false|false||epigastricnull|Food allergenic extracts|Drug|false|false||food
null|Food|Drug|false|false||food
null|Food allergenic extracts|Drug|false|false||foodnull|With intensity|Modifier|false|false||severity
null|Severities|Modifier|false|false||severitynull|Course|Time|false|false||coursenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|SON gene|Finding|false|false||sonnull|Son (person)|Subject|false|false||sonnull|Songhay Languages|Entity|false|false||sonnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Confusion|Disorder|false|false||confusionnull|Clouded consciousness|Finding|false|false||confusionnull|Alert brand of caffeine|Drug|false|false||alert
null|Alert brand of caffeine|Drug|false|false||alertnull|Mentally alert|Finding|false|false||alert
null|Consciousness clear|Finding|false|false||alert
null|Alert note|Finding|false|false||alert
null|Alert|Finding|false|false||alertnull|null|Attribute|false|false||alertnull|Oriented to place|Finding|false|false||orientednull|Orientation, Spatial|Modifier|false|false||orientednull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Recent|Time|false|false||recentlynull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Fever symptoms (finding)|Finding|true|false||fever
null|Fever|Finding|true|false||fevernull|Chills|Finding|true|false||chillsnull|Dyspnea|Finding|true|false||shortness of breathnull|null|Attribute|true|false||shortness of breathnull|Breath|Finding|false|false||breathnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Dysuria|Finding|false|false||dysurianull|Loose stool|Finding|false|false||loose stoolnull|Loose|Modifier|false|false||loosenull|2-(4-ethoxybenzyl)-1-diethylaminoethyl-5-isothiocyanatobenzimidazole|Drug|false|false||bit
null|2-(4-ethoxybenzyl)-1-diethylaminoethyl-5-isothiocyanatobenzimidazole|Drug|false|false||bit
null|PTPNS1 protein, human|Drug|false|false||bitnull|Breast-Impact of Treatment Scale|Finding|false|false||bit
null|PTPNS1 protein, human|Finding|false|false||bit
null|SIRPA gene|Finding|false|false||bit
null|SIRPA wt Allele|Finding|false|false||bitnull|bit - unit of measure|LabModifier|false|false||bitnull|Greater Than|LabModifier|false|false||more thannull|More|LabModifier|false|false||morenull|Usual|Modifier|false|false||usualnull|lactulose|Drug|false|false||lactulose
null|lactulose|Drug|false|false||lactulosenull|Use - dosing instruction imperative|Finding|false|false||use
null|utilization qualifier|Finding|false|false||use
null|Usage|Finding|false|false||usenull|Laboratory test finding|Lab|false|false||Labsnull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|lactate|Drug|false|false||lactate
null|lactate|Drug|false|false||lactate
null|Lactates|Drug|false|false||lactatenull|Lactic acid measurement|Procedure|false|false||lactatenull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||ASTnull|Atypical Spitz Nevus|Disorder|false|false||ASTnull|SLC17A5 wt Allele|Finding|false|false||AST
null|SLC17A5 gene|Finding|false|false||AST
null|GOT1 gene|Finding|false|false||ASTnull|Asterion|Anatomy|false|false||ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Leukocytosis|Disorder|true|false||leukocytosisnull|Blood leukocyte number above reference range|Finding|true|false||leukocytosisnull|Ascitic Fluid|Finding|false|false||Ascitic fluidnull|Ascitic|Modifier|false|false||Asciticnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Leukocytes|Anatomy|false|false||WBCnull|morphine sulfate|Drug|false|false||Morphine Sulfate
null|morphine sulfate|Drug|false|false||Morphine Sulfatenull|morphine|Drug|false|false||Morphine
null|morphine|Drug|false|false||Morphinenull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||Sulfate
null|Sulfates, Inorganic|Drug|false|false||Sulfate
null|sulfate ion|Drug|false|false||Sulfate
null|sulfate ion|Drug|false|false||Sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||Sulfatenull|Once - dosing instruction fragment|Finding|false|false||ONCEnull|Once (schedule frequency)|Time|false|false||ONCEnull|MR1 gene|Finding|false|false||MR1
null|PNKD gene|Finding|false|false||MR1null|Cocktail|Drug|false|false||cocktailnull|hepatitis C virus|Disorder|false|false||HCV
null|Hepatitis C|Disorder|false|false||HCVnull|Liver Cirrhosis|Disorder|false|false||Cirrhosis
null|Cirrhosis|Disorder|false|false||Cirrhosisnull|Genotype determination|Procedure|false|false||genotypenull|Genotype|Subject|false|false||genotypenull|HIV Vaccine|Drug|false|false||HIV
null|HIV Vaccine|Drug|false|false||HIVnull|HIV Infections|Disorder|false|false||HIV
null|HIV|Disorder|false|false||HIVnull|Antiretroviral Therapy, Highly Active|Procedure|false|false||HAARTnull|CD4 Count determination procedure|Procedure|false|false||CD4 count
null|CD4 Expressing Cell Count|Procedure|false|false||CD4 countnull|T-Cell Surface Glycoprotein CD4, human|Drug|false|false||CD4
null|T-Cell Surface Glycoprotein CD4, human|Drug|false|false||CD4
null|CD4 Antigens|Drug|false|false||CD4
null|CD4 Antigens|Drug|false|false||CD4null|CD4 Antigens|Finding|false|false||CD4
null|CD4 gene|Finding|false|false||CD4null|Count Dosing Unit|LabModifier|false|false||count
null|Count|LabModifier|false|false||countnull|HIV viral load|Procedure|false|false||HIV viral loadnull|HIV Vaccine|Drug|false|false||HIV
null|HIV Vaccine|Drug|false|false||HIVnull|HIV Infections|Disorder|false|false||HIV
null|HIV|Disorder|false|false||HIVnull|Viral Load result|Finding|false|false||viral loadnull|Viral load (procedure)|Procedure|false|false||viral loadnull|Viral|Finding|false|false||viralnull|Load - Remote control command|Finding|false|false||loadnull|Load Device|Device|false|false||loadnull|Loading Technique|Event|false|false||loadnull|Undetectable|Attribute|false|false||undetectablenull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|bentiromide|Drug|false|false||PFT
null|bentiromide|Drug|false|false||PFTnull|fluorouracil/melphalan/tamoxifen|Procedure|false|false||PFT
null|Pulmonary function tests|Procedure|false|false||PFTnull|area PFt|Anatomy|false|false||PFTnull|Forced Vital Capacity|Lab|false|false||FVCnull|Pulmonary Function Test/Forced Expiratory Volume 1|Procedure|false|false||FEV1null|null|Attribute|false|false||FEV1null|Volume expired during 1.0 s of forced expiration|LabModifier|false|false||FEV1null|MAJOR AFFECTIVE DISORDER 4|Disorder|false|false||Bipolar Affective Disorder
null|MAJOR AFFECTIVE DISORDER 9|Disorder|false|false||Bipolar Affective Disorder
null|Bipolar Disorder|Disorder|false|false||Bipolar Affective Disorder
null|MAJOR AFFECTIVE DISORDER 2|Disorder|false|false||Bipolar Affective Disorder
null|MAJOR AFFECTIVE DISORDER 1|Disorder|false|false||Bipolar Affective Disorder
null|MAJOR AFFECTIVE DISORDER 8|Disorder|false|false||Bipolar Affective Disorder
null|MAJOR AFFECTIVE DISORDER 6|Disorder|false|false||Bipolar Affective Disorder
null|MAJOR AFFECTIVE DISORDER 7|Disorder|false|false||Bipolar Affective Disordernull|Bipolar|Modifier|false|false||Bipolarnull|Mood Disorders|Disorder|false|false||Affective Disordernull|Disease|Disorder|false|false||Disordernull|6-pyruvoyl-tetrahydropterin synthase deficiency|Disorder|false|false||PTSD
null|Post-Traumatic Stress Disorder|Disorder|false|false||PTSDnull|cocaine|Drug|false|false||cocaine
null|cocaine|Drug|false|false||cocaine
null|cocaine|Drug|false|false||cocaine
null|cocaine|Drug|false|false||cocainenull|Poisoning by cocaine|Disorder|false|false||cocainenull|Cocaine measurement|Procedure|false|false||cocainenull|heroin abuse|Disorder|false|false||heroin abusenull|heroin|Drug|false|false||heroin
null|heroin|Drug|false|false||heroin
null|heroin|Drug|false|false||heroinnull|Poisoning by heroin|Disorder|false|false||heroinnull|Drug abuse|Disorder|false|false||abusenull|Victim of abuse (finding)|Finding|false|false||abusenull|Abuse|Event|false|false||abusenull|Malignant neoplasm of skin|Disorder|false|false||of skin cancernull|Malignant neoplasm of skin|Disorder|false|false||skin cancernull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false||skinnull|Skin Specimen Source Code|Finding|false|false||skin
null|Skin Specimen|Finding|false|false||skinnull|Skin, Human|Anatomy|false|false||skin
null|Skin|Anatomy|false|false||skinnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Patient-Reported|Finding|false|false||patient reportnull|Report source - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Relationship modifier - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Report (document)|Finding|false|false||reportnull|Reporting|Procedure|false|false||reportnull|null|Attribute|false|false||reportnull|Total|Modifier|false|false||totalnull|Sibling|Subject|false|false||siblingsnull|Brother - courtesy title|Finding|false|false||brother
null|Relationship - Brother|Finding|false|false||brothernull|Brothers|Subject|false|false||brothernull|In Touch|Device|false|false||in touchnull|Touch Perception|Finding|false|false||touch
null|Touch sensation|Finding|false|false||touchnull|Therapeutic Touch|Procedure|false|false||touchnull|Tactile|Modifier|false|false||touchnull|Awareness|Finding|true|false||awarenull|Known|Modifier|false|false||knownnull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Disease|Disorder|false|false||diseasenull|ErbB Receptors|Drug|false|false||her family
null|ErbB Receptors|Drug|false|false||her familynull|ErbB Receptors|Finding|false|false||her familynull|Entity Name Part Type - family|Finding|false|false||family
null|Last Name|Finding|false|false||family
null|Living Arrangement - Family|Finding|false|false||family
null|Family (taxonomic)|Finding|false|false||family
null|Family Collection|Finding|false|false||familynull|Family|Subject|false|false||familynull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|physical examination (physical finding)|Finding|false|false||PHYSICAL EXAMnull|Physical Examination|Procedure|false|false||PHYSICAL EXAMnull|physical examination (physical finding)|Finding|false|false||PHYSICAL
null|Physical|Finding|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||PHYSICALnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GENERALnull|General medical service|Procedure|false|false||GENERALnull|Generalized|Modifier|false|false||GENERALnull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|RIGHT SIDE (USED TO IDENTIFY PROCEDURES PERFORMED ON THE RIGHT SIDE OF THE BODY)|Modifier|false|false||right side
null|Right|Modifier|false|false||right sidenull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Side|Modifier|false|false||sidenull|HEENT|Anatomy|false|false||HEENTnull|Pupil equal round and reacting to light|Finding|false|false||PERRLnull|Anicteric|Finding|false|false||anictericnull|Scleral Diseases|Disorder|false|false||scleranull|examination of sclera|Procedure|false|false||scleranull|Sclera|Anatomy|false|false||scleranull|Pink color|Modifier|false|false||pinknull|Malignant neoplasm of conjunctiva|Disorder|false|false||conjunctiva
null|Benign neoplasm of conjunctiva|Disorder|false|false||conjunctiva
null|Conjunctival Diseases|Disorder|false|false||conjunctivanull|Specimen Type - Conjunctiva|Finding|false|false||conjunctiva
null|null|Finding|false|false||conjunctivanull|examination of conjunctiva|Procedure|false|false||conjunctiva
null|Procedure on conjunctiva|Procedure|false|false||conjunctivanull|Structure of palpebral conjunctiva|Anatomy|false|false||conjunctiva
null|conjunctiva|Anatomy|false|false||conjunctivanull|Myelofibrosis|Disorder|false|false||MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false||MMMnull|Language Ability Proficiency - Good|Finding|false|false||good
null|Language Proficiency - Good|Finding|false|false||goodnull|Specimen Quality - Good|Modifier|false|false||good
null|Good|Modifier|false|false||goodnull|Dentition|Anatomy|false|false||dentition
null|Tooth structure|Anatomy|false|false||dentitionnull|Passive joint movement of neck (finding)|Finding|false|false||NECK
null|Neck problem|Finding|false|false||NECKnull|dendritic spine neck|Anatomy|false|false||NECK
null|Neck|Anatomy|false|false||NECKnull|Supple neck|Finding|false|false||supple necknull|Supple|Finding|false|false||supplenull|Passive joint movement of neck (finding)|Finding|false|false||neck
null|Neck problem|Finding|false|false||necknull|dendritic spine neck|Anatomy|false|false||neck
null|Neck|Anatomy|false|false||necknull|Leukocyte adhesion deficiency type 1|Disorder|true|false||LAD
null|Leukocyte adhesion deficiency|Disorder|true|false||LADnull|ITGB2 wt Allele|Finding|true|false||LAD
null|DLD gene|Finding|true|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false||LADnull|Ladino Language|Entity|true|false||LADnull|Jugular venous engorgement|Finding|true|false||JVDnull|Cardiac attachment|Finding|false|false||CARDIACnull|Heart|Anatomy|false|false||CARDIACnull|Cardiac - anatomy qualifier|Modifier|false|false||CARDIACnull|Heart murmur|Finding|true|false||murmursnull|Pericardial friction rub|Finding|true|false||rubsnull|Lung diseases|Disorder|false|false||LUNGnull|Lung Problem|Finding|false|false||LUNGnull|Chest>Lung|Anatomy|false|false||LUNG
null|Lung|Anatomy|false|false||LUNGnull|cetrimonium bromide|Drug|false|false||CTABnull|Wheezing|Finding|true|false||wheezesnull|Basilar Rales|Finding|true|false||rales
null|Rales|Finding|true|false||ralesnull|Rhonchi|Finding|true|false||rhonchinull|Use of accessory muscles|Finding|true|false||use of accessory musclesnull|Use of|Finding|true|false||use ofnull|Use - dosing instruction imperative|Finding|true|false||use
null|utilization qualifier|Finding|true|false||use
null|Usage|Finding|true|false||usenull|Accessory skeletal muscle|Disorder|false|false||accessory musclesnull|Accessory|Device|false|false||accessorynull|Set of muscles|Anatomy|false|false||muscles
null|Muscle (organ)|Anatomy|false|false||muscles
null|Muscle Tissue|Anatomy|false|false||musclesnull|Malignant neoplasm of abdomen|Disorder|false|false||ABDOMENnull|Abdomen problem|Finding|false|false||ABDOMENnull|Abdomen|Anatomy|false|false||ABDOMEN
null|Abdominal Cavity|Anatomy|false|false||ABDOMENnull|Dilated|Finding|false|false||distendednull|Distended|Modifier|false|false||distendednull|Fluid thrill in abdomen|Finding|false|false||fluid wavenull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|WASF1 gene|Finding|false|false||wavenull|null|Phenomenon|false|false||wavenull|Tension|Disorder|true|false||tensenull|Feeling tense|Finding|true|false||tensenull|All extremities|Anatomy|false|false||EXTREMITIES
null|Limb structure|Anatomy|false|false||EXTREMITIESnull|Cyanosis|Finding|true|false||cyanosisnull|Clubbing|Disorder|true|false||clubbingnull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|PURPOSE (pharmacologic preparation)|Drug|false|false||purpose
null|PURPOSE (pharmacologic preparation)|Drug|false|false||purposenull|Purpose|Finding|false|false||purposenull|null|Drug|false|false||PULSESnull|Physiologic pulse|Finding|false|false||PULSESnull|Pulse taking|Procedure|false|false||PULSESnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Neurology speciality|Title|false|false||NEUROnull|Neurologic (qualifier value)|Modifier|false|false||NEUROnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|abscisic aldehyde oxidase activity|Finding|false|false||AAO3null|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||SKIN
null|Skin and subcutaneous tissue disorders|Disorder|false|false||SKINnull|Skin Specimen Source Code|Finding|false|false||SKIN
null|Skin Specimen|Finding|false|false||SKINnull|Skin, Human|Anatomy|false|false||SKIN
null|Skin|Anatomy|false|false||SKINnull|Feels warm|Finding|false|false||warmnull|warming process|Phenomenon|false|false||warmnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Excoriation|Disorder|true|false||excoriationsnull|Lesion|Finding|true|false||lesionsnull|Skin rash|Finding|false|false||rashes
null|Exanthema|Finding|false|false||rashesnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|physical examination (physical finding)|Finding|false|false||PHYSICAL EXAMnull|Physical Examination|Procedure|false|false||PHYSICAL EXAMnull|physical examination (physical finding)|Finding|false|false||PHYSICAL
null|Physical|Finding|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||PHYSICALnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GENERALnull|General medical service|Procedure|false|false||GENERALnull|Generalized|Modifier|false|false||GENERALnull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|RIGHT SIDE (USED TO IDENTIFY PROCEDURES PERFORMED ON THE RIGHT SIDE OF THE BODY)|Modifier|false|false||right side
null|Right|Modifier|false|false||right sidenull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Side|Modifier|false|false||sidenull|HEENT|Anatomy|false|false||HEENTnull|Pupil equal round and reacting to light|Finding|false|false||PERRLnull|Anicteric|Finding|false|false||anictericnull|Scleral Diseases|Disorder|false|false||scleranull|examination of sclera|Procedure|false|false||scleranull|Sclera|Anatomy|false|false||scleranull|Pink color|Modifier|false|false||pinknull|Malignant neoplasm of conjunctiva|Disorder|false|false||conjunctiva
null|Benign neoplasm of conjunctiva|Disorder|false|false||conjunctiva
null|Conjunctival Diseases|Disorder|false|false||conjunctivanull|Specimen Type - Conjunctiva|Finding|false|false||conjunctiva
null|null|Finding|false|false||conjunctivanull|examination of conjunctiva|Procedure|false|false||conjunctiva
null|Procedure on conjunctiva|Procedure|false|false||conjunctivanull|Structure of palpebral conjunctiva|Anatomy|false|false||conjunctiva
null|conjunctiva|Anatomy|false|false||conjunctivanull|Myelofibrosis|Disorder|false|false||MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false||MMMnull|Language Ability Proficiency - Good|Finding|false|false||good
null|Language Proficiency - Good|Finding|false|false||goodnull|Specimen Quality - Good|Modifier|false|false||good
null|Good|Modifier|false|false||goodnull|Dentition|Anatomy|false|false||dentition
null|Tooth structure|Anatomy|false|false||dentitionnull|Passive joint movement of neck (finding)|Finding|false|false||NECK
null|Neck problem|Finding|false|false||NECKnull|dendritic spine neck|Anatomy|false|false||NECK
null|Neck|Anatomy|false|false||NECKnull|Supple neck|Finding|false|false||supple necknull|Supple|Finding|false|false||supplenull|Passive joint movement of neck (finding)|Finding|false|false||neck
null|Neck problem|Finding|false|false||necknull|dendritic spine neck|Anatomy|false|false||neck
null|Neck|Anatomy|false|false||necknull|Leukocyte adhesion deficiency type 1|Disorder|true|false||LAD
null|Leukocyte adhesion deficiency|Disorder|true|false||LADnull|ITGB2 wt Allele|Finding|true|false||LAD
null|DLD gene|Finding|true|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false||LADnull|Ladino Language|Entity|true|false||LADnull|Jugular venous engorgement|Finding|true|false||JVDnull|Cardiac attachment|Finding|false|false||CARDIACnull|Heart|Anatomy|false|false||CARDIACnull|Cardiac - anatomy qualifier|Modifier|false|false||CARDIACnull|Heart murmur|Finding|true|false||murmursnull|Pericardial friction rub|Finding|true|false||rubsnull|Lung diseases|Disorder|false|false||LUNGnull|Lung Problem|Finding|false|false||LUNGnull|Chest>Lung|Anatomy|false|false||LUNG
null|Lung|Anatomy|false|false||LUNGnull|cetrimonium bromide|Drug|false|false||CTABnull|Wheezing|Finding|true|false||wheezesnull|Basilar Rales|Finding|true|false||rales
null|Rales|Finding|true|false||ralesnull|Rhonchi|Finding|true|false||rhonchinull|Use of accessory muscles|Finding|true|false||use of accessory musclesnull|Use of|Finding|true|false||use ofnull|Use - dosing instruction imperative|Finding|true|false||use
null|utilization qualifier|Finding|true|false||use
null|Usage|Finding|true|false||usenull|Accessory skeletal muscle|Disorder|false|false||accessory musclesnull|Accessory|Device|false|false||accessorynull|Set of muscles|Anatomy|false|false||muscles
null|Muscle (organ)|Anatomy|false|false||muscles
null|Muscle Tissue|Anatomy|false|false||musclesnull|Malignant neoplasm of abdomen|Disorder|false|false||ABDOMENnull|Abdomen problem|Finding|false|false||ABDOMENnull|Abdomen|Anatomy|false|false||ABDOMEN
null|Abdominal Cavity|Anatomy|false|false||ABDOMENnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|Decreasing|Finding|false|false||decreased
null|Reduced|Finding|false|false||decreasednull|Decreased|LabModifier|false|false||decreasednull|Pathological Dilatation|Finding|true|false||distension
null|Distention|Finding|true|false||distensionnull|Tension|Disorder|true|false||tensenull|Feeling tense|Finding|true|false||tensenull|All extremities|Anatomy|false|false||EXTREMITIES
null|Limb structure|Anatomy|false|false||EXTREMITIESnull|Cyanosis|Finding|true|false||cyanosisnull|Clubbing|Disorder|true|false||clubbingnull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|PURPOSE (pharmacologic preparation)|Drug|false|false||purpose
null|PURPOSE (pharmacologic preparation)|Drug|false|false||purposenull|Purpose|Finding|false|false||purposenull|null|Drug|false|false||PULSESnull|Physiologic pulse|Finding|false|false||PULSESnull|Pulse taking|Procedure|false|false||PULSESnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Neurology speciality|Title|false|false||NEUROnull|Neurologic (qualifier value)|Modifier|false|false||NEUROnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|abscisic aldehyde oxidase activity|Finding|false|false||AAO3null|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||SKIN
null|Skin and subcutaneous tissue disorders|Disorder|false|false||SKINnull|Skin Specimen Source Code|Finding|false|false||SKIN
null|Skin Specimen|Finding|false|false||SKINnull|Skin, Human|Anatomy|false|false||SKIN
null|Skin|Anatomy|false|false||SKINnull|Feels warm|Finding|false|false||warmnull|warming process|Phenomenon|false|false||warmnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Excoriation|Disorder|true|false||excoriationsnull|Lesion|Finding|true|false||lesionsnull|Skin rash|Finding|false|false||rashes
null|Exanthema|Finding|false|false||rashesnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||ASTnull|Atypical Spitz Nevus|Disorder|false|false||ASTnull|SLC17A5 wt Allele|Finding|false|false||AST
null|SLC17A5 gene|Finding|false|false||AST
null|GOT1 gene|Finding|false|false||ASTnull|Asterion|Anatomy|false|false||ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Alkaline Phosphatase|Drug|false|false||AlkPhos
null|Alkaline Phosphatase|Drug|false|false||AlkPhosnull|Blood albumin|Procedure|false|false||BLOOD Albuminnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Albumin|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumin|Drug|false|false||Albuminnull|Albumin metabolic function|Finding|false|false||Albumin
null|ALB gene|Finding|false|false||Albuminnull|Albumin measurement|Procedure|false|false||Albuminnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|lactate in blood (lab test)|Procedure|false|false||BLOOD Lactatenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|lactate|Drug|false|false||Lactate
null|lactate|Drug|false|false||Lactate
null|Lactates|Drug|false|false||Lactatenull|Lactic acid measurement|Procedure|false|false||Lactatenull|Laboratory test finding|Lab|false|false||LABSnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Ascites|Disorder|false|false||ASCITESnull|Peritoneal Effusion|Finding|false|false||ASCITESnull|Leukocytes|Anatomy|false|false||WBCnull|5'-Inosinic acid, 2'-deoxy-2'-fluoro-, homopolymer|Drug|false|false||Polys
null|Poly A|Drug|false|false||Polysnull|Lymph|Finding|false|false||Lymphsnull|Monos|Drug|false|false||Monos
null|Mono-S|Drug|false|false||Monos
null|Monos|Drug|false|false||Monosnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Ascites|Disorder|false|false||ASCITESnull|Peritoneal Effusion|Finding|false|false||ASCITESnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Microbiology Diagnostic Service Section ID|Finding|false|false||MICROBIOLOGY
null|Microbiological|Finding|false|false||MICROBIOLOGY
null|Microbiology - Laboratory Class|Finding|false|false||MICROBIOLOGYnull|Microbiology procedure|Procedure|false|false||MICROBIOLOGYnull|Science of Microbiology|Title|false|false||MICROBIOLOGYnull|Peritoneal fluid (substance)|Finding|false|false||PERITONEAL FLUIDnull|Peritoneal fluid analysis|Procedure|false|false||PERITONEAL FLUIDnull|peritoneal|Anatomy|false|false||PERITONEAL
null|Peritoneum|Anatomy|false|false||PERITONEALnull|fluid - substance|Drug|false|false||FLUID
null|Liquid substance|Drug|false|false||FLUIDnull|Fluid Specimen Code|Finding|false|false||FLUIDnull|Fluid behavior|Modifier|false|false||FLUIDnull|Gram's stain|Drug|false|false||GRAM STAIN
null|Gram's stain|Drug|false|false||GRAM STAINnull|Bacterial stain, routine|Procedure|false|false||GRAM STAINnull|gram|LabModifier|false|false||GRAMnull|Stains|Drug|false|false||STAINnull|Staining method|Procedure|false|false||STAINnull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|granulocyte|Anatomy|false|false||POLYMORPHONUCLEAR LEUKOCYTES
null|neutrophil|Anatomy|false|false||POLYMORPHONUCLEAR LEUKOCYTESnull|Specimen Type - Leukocytes|Finding|true|false||LEUKOCYTES
null|null|Finding|true|false||LEUKOCYTESnull|Leukocytes|Anatomy|false|false||LEUKOCYTESnull|Microorganisms seen|Finding|false|false||MICROORGANISMS SEENnull|Microorganism|Entity|true|false||MICROORGANISMSnull|fluid - substance|Drug|false|false||FLUID
null|Liquid substance|Drug|false|false||FLUIDnull|Fluid Specimen Code|Finding|false|false||FLUIDnull|Fluid behavior|Modifier|false|false||FLUIDnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Growth & development aspects|Finding|true|false||GROWTH
null|Tissue Growth|Finding|true|false||GROWTH
null|Growth|Finding|true|false||GROWTH
null|growth aspects|Finding|true|false||GROWTHnull|Growth action|Phenomenon|true|false||GROWTHnull|Anaerobic microbial culture|Procedure|false|false||ANAEROBIC CULTUREnull|Anaerobic|Modifier|false|false||ANAEROBICnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Preliminary|Time|false|false||Preliminarynull|Growth & development aspects|Finding|true|false||GROWTH
null|Tissue Growth|Finding|true|false||GROWTH
null|Growth|Finding|true|false||GROWTH
null|growth aspects|Finding|true|false||GROWTHnull|Growth action|Phenomenon|true|false||GROWTHnull|Vancomycin-Resistant Enterococci|Entity|false|false||VREnull|Toxicology screen, general (procedure)|Procedure|false|false||screen
null|Disease Screening|Procedure|false|false||screen
null|Screening for cancer|Procedure|false|false||screen
null|Screening procedure|Procedure|false|false||screennull|Screen Device|Device|false|false||screennull|Vancomycin-Resistant Enterococci|Entity|true|false||VREnull|Imaging problem|Finding|false|false||IMAGINGnull|Diagnostic Imaging|Procedure|false|false||IMAGING
null|Imaging Techniques|Procedure|false|false||IMAGINGnull|Imaging Technology|Title|false|false||IMAGINGnull|Scientific Study|Procedure|false|false||STUDIESnull|Plain chest X-ray|Procedure|false|false||CXRnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Cardiovascular disease+Pulmonary disease|Disorder|false|false||cardiopulmonarynull|Cardiopulmonary|Anatomy|false|false||cardiopulmonarynull|Process Pharmacologic Substance|Drug|true|false||processnull|Process (qualifier value)|Finding|true|false||processnull|bony process|Anatomy|false|false||processnull|Process|Phenomenon|true|false||processnull|Cirrhotic|Modifier|false|false||Cirrhoticnull|Mild splenomegaly|Finding|false|false||mild splenomegalynull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Splenomegaly|Finding|false|false||splenomegalynull|Ascites|Disorder|false|false||ascitesnull|Peritoneal Effusion|Finding|false|false||ascitesnull|Solid Dose Form|Drug|false|false||solid
null|solid substance|Drug|false|false||solidnull|Solid|Modifier|false|false||solidnull|Left lobe of liver|Anatomy|false|false||left lobe of the livernull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|AKT1S1 wt Allele|Finding|false|false||lobe
null|AKT1S1 gene|Finding|false|false||lobenull|lobe|Anatomy|false|false||lobenull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|patient appearance regarding mental status exam|Procedure|false|false||appearancenull|null|Attribute|false|false||appearancenull|Personal appearance|Subject|false|false||appearancenull|Appearance|Modifier|false|false||appearancenull|Kind of quantity - Appearance|LabModifier|false|false||appearancenull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||ASTnull|Atypical Spitz Nevus|Disorder|false|false||ASTnull|SLC17A5 wt Allele|Finding|false|false||AST
null|SLC17A5 gene|Finding|false|false||AST
null|GOT1 gene|Finding|false|false||ASTnull|Asterion|Anatomy|false|false||ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Alkaline Phosphatase|Drug|false|false||AlkPhos
null|Alkaline Phosphatase|Drug|false|false||AlkPhosnull|Blood albumin|Procedure|false|false||BLOOD Albuminnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Albumin|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumin|Drug|false|false||Albuminnull|Albumin metabolic function|Finding|false|false||Albumin
null|ALB gene|Finding|false|false||Albuminnull|Albumin measurement|Procedure|false|false||Albuminnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|HIV Vaccine|Drug|false|false||HIV
null|HIV Vaccine|Drug|false|false||HIVnull|HIV Infections|Disorder|false|false||HIV
null|HIV|Disorder|false|false||HIVnull|Antiretroviral Therapy, Highly Active|Procedure|false|false||HAARTnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|hepatitis C virus|Disorder|false|false||HCV
null|Hepatitis C|Disorder|false|false||HCVnull|Liver Cirrhosis|Disorder|false|false||cirrhosis
null|Cirrhosis|Disorder|false|false||cirrhosisnull|Decompensated|Modifier|false|false||decompensatednull|Ascites|Disorder|false|false||ascitesnull|Peritoneal Effusion|Finding|false|false||ascitesnull|Biweekly|Time|false|false||biweeklynull|Therapeutic brand of coal tar|Drug|false|false||therapeutic
null|Therapeutic brand of coal tar|Drug|false|false||therapeuticnull|Therapeutic - Location Service Code|Finding|false|false||therapeutic
null|Therapeutic|Finding|false|false||therapeuticnull|Therapeutic procedure|Procedure|false|false||therapeuticnull|Paracentesis|Procedure|false|false||paracentesesnull|Hepatic Encephalopathy|Disorder|false|false||hepatic encephalopathynull|Hepatic|Anatomy|false|false||hepaticnull|Encephalopathies|Disorder|false|false||encephalopathynull|Transplant|Finding|false|false||transplant
null|Transplanted organ and tissue status|Finding|false|false||transplantnull|Transplantation|Procedure|false|false||transplantnull|Transplanted tissue|Anatomy|false|false||transplantnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Comorbidity|Finding|false|false||comorbiditiesnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false||abdnull|ABD (body structure)|Anatomy|false|false||abd
null|Abdomen|Anatomy|false|false||abdnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Goals of Care|Procedure|false|false||Goals of carenull|What subject filter - Goals|Finding|false|false||Goals
null|objective (goal)|Finding|false|false||Goals
null|treatment goals|Finding|false|false||Goalsnull|null|Attribute|false|false||Goalsnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|desire|Finding|false|false||desirenull|peace|Finding|false|false||peacenull|Feel Tired question|Finding|false|false||tired
null|Fatigue|Finding|false|false||tired
null|Feeling tired|Finding|false|false||tirednull|Fighting|Finding|false|false||fightingnull|End-stage|Modifier|false|false||end stagenull|Endoglin, human|Drug|false|false||end
null|Endoglin, human|Drug|false|false||endnull|end - ActRelationshipCheckpoint|Finding|false|false||end
null|ENG gene|Finding|false|false||end
null|ENG wt Allele|Finding|false|false||endnull|Stop (qualifier value)|Time|false|false||endnull|End|Modifier|false|false||endnull|Tumor stage|Attribute|false|false||stagenull|Stage|Time|false|false||stage
null|Phase|Time|false|false||stagenull|Liver diseases|Disorder|false|false||liver disease
null|Hepatobiliary Disorder|Disorder|false|false||liver diseasenull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Disease|Disorder|false|false||diseasenull|Language Ability Proficiency - Good|Finding|false|false||good
null|Language Proficiency - Good|Finding|false|false||goodnull|Specimen Quality - Good|Modifier|false|false||good
null|Good|Modifier|false|false||goodnull|Quality|Modifier|false|false||qualitynull|Life|Finding|false|false||lifenull|Laser-Induced Fluorescence Endoscopy|Procedure|false|false||lifenull|Representation (action)|Event|false|false||representativenull|Hospice Care|Procedure|false|false||hospicenull|Hospice (environment)|Device|false|false||hospicenull|Hospice (environment)|Entity|false|false||hospicenull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Hospice Care|Procedure|false|false||hospicenull|Hospice (environment)|Device|false|false||hospicenull|Hospice (environment)|Entity|false|false||hospicenull|conversation|Finding|false|false||conversationnull|Disabled Person Code - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|Relationship modifier - Patient|Finding|false|false||patient
null|null|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|CODE STATUS|Procedure|false|false||code statusnull|MDF Attribute Type - Code|Finding|false|false||code
null|A Codes|Finding|false|false||code
null|Code|Finding|false|false||codenull|Coding|Event|false|false||codenull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|Probably|Finding|false|false||probably
null|Probable diagnosis|Finding|false|false||probablynull|daunorubicin|Drug|false|false||DNR
null|daunorubicin|Drug|false|false||DNRnull|Do-Not-Resuscitate Orders|Finding|false|false||DNR
null|Do not resuscitate status|Finding|false|false||DNRnull|null|Attribute|false|false||DNRnull|SON gene|Finding|false|false||sonnull|Son (person)|Subject|false|false||sonnull|Songhay Languages|Entity|false|false||sonnull|Hereditary Coproporphyria|Disorder|false|false||HCPnull|PTPN6 wt Allele|Finding|false|false||HCP
null|CPOX gene|Finding|false|false||HCP
null|AMBP wt Allele|Finding|false|false||HCP
null|PTPN6 gene|Finding|false|false||HCP
null|AMBP gene|Finding|false|false||HCPnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Full|Modifier|false|false||fullnull|MDF Attribute Type - Code|Finding|false|false||code
null|A Codes|Finding|false|false||code
null|Code|Finding|false|false||codenull|Coding|Event|false|false||codenull|null|Finding|false|false||catheternull|catheter device|Device|false|false||catheter
null|XXX>Catheter|Device|false|false||catheternull|Paracentesis|Procedure|false|false||paracentesesnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Hospice Care|Procedure|false|false||hospicenull|Hospice (environment)|Device|false|false||hospicenull|Hospice (environment)|Entity|false|false||hospicenull|hepatitis C virus|Disorder|false|false||HCV
null|Hepatitis C|Disorder|false|false||HCVnull|Liver Cirrhosis|Disorder|false|false||cirrhosis
null|Cirrhosis|Disorder|false|false||cirrhosisnull|Ascites|Disorder|false|false||ascitesnull|Peritoneal Effusion|Finding|false|false||ascitesnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Presentation|Finding|false|false||presentednull|Patient Outcome - Worsening|Finding|false|false||worseningnull|Worsening (qualifier value)|Modifier|false|false||worseningnull|Ascites|Disorder|false|false||ascitesnull|Peritoneal Effusion|Finding|false|false||ascitesnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Initially|Time|false|false||initiallynull|tramadol|Drug|false|false||tramadol
null|tramadol|Drug|false|false||tramadolnull|Tramadol measurement (procedure)|Procedure|false|false||tramadolnull|morphine|Drug|false|false||morphine
null|morphine|Drug|false|false||morphinenull|Paracentesis|Procedure|false|false||paracentesisnull|removal technique|Procedure|false|false||removal
null|Excision|Procedure|false|false||removal
null|Extraction|Procedure|false|false||removalnull|Removing (action)|Event|false|false||removalnull|Albumin|Drug|false|false||albumin
null|Albumins|Drug|false|false||albumin
null|Albumins|Drug|false|false||albumin
null|Albumin|Drug|false|false||albuminnull|Albumin metabolic function|Finding|false|false||albumin
null|ALB gene|Finding|false|false||albuminnull|Albumin measurement|Procedure|false|false||albuminnull|Scientific Study|Procedure|false|false||Studiesnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Improvement|Finding|false|false||improvementnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Hyperkalemia|Finding|false|false||Hyperkalemia
null|Serum potassium level above reference range|Finding|false|false||Hyperkalemianull|Hospitalization|Procedure|false|false||hospitalizationnull|Hyperkalemia|Finding|false|false||hyperkalemia
null|Serum potassium level above reference range|Finding|false|false||hyperkalemianull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|Changing|Finding|true|false||changesnull|Changed status|LabModifier|false|false||changesnull|Aftercare|Procedure|false|false||After treatmentnull|Post-Therapy|Time|false|false||After treatmentnull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|calcium gluconate|Drug|false|false||calcium gluconate
null|calcium gluconate|Drug|false|false||calcium gluconatenull|CALCIUM SUPPLEMENTS|Drug|false|false||calcium
null|calcium|Drug|false|false||calcium
null|calcium|Drug|false|false||calcium
null|calcium|Drug|false|false||calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||calcium
null|Calcium, Dietary|Drug|false|false||calcium
null|Calcium [EPC]|Drug|false|false||calcium
null|Calcium Drug Class|Drug|false|false||calciumnull|Calcium metabolic function|Finding|false|false||calciumnull|Calcium measurement|Procedure|false|false||calciumnull|gluconate|Drug|false|false||gluconate
null|Gluconates|Drug|false|false||gluconate
null|Gluconates|Drug|false|false||gluconate
null|gluconate|Drug|false|false||gluconate
null|gluconate|Drug|false|false||gluconatenull|insulin, regular, human|Drug|false|false||insulin
null|Insulin [EPC]|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulinnull|INS gene|Finding|false|false||insulinnull|Insulin measurement|Procedure|false|false||insulinnull|persistently|Finding|false|false||persistentlynull|Hepatic Encephalopathy|Disorder|false|false||Hepatic encephalopathynull|Hepatic|Anatomy|false|false||Hepaticnull|Encephalopathies|Disorder|false|false||encephalopathynull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Mental state|Finding|false|false||mental statusnull|null|Attribute|false|false||mental status
null|null|Attribute|false|false||mental statusnull|Psyche structure|Finding|false|false||mentalnull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|On admission|Time|false|false||on admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|rifaximin|Drug|false|false||rifaximin
null|rifaximin|Drug|false|false||rifaximinnull|lactulose|Drug|false|false||lactulose
null|lactulose|Drug|false|false||lactulosenull|In-House|Finding|false|false||in-housenull|House (environment)|Device|false|false||housenull|Home environment|Modifier|false|false||housenull|At discharge|Time|false|false||at dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Chronic - Admission Level of Care Code|Finding|false|false||CHRONICnull|Provision of recurring care for chronic illness|Procedure|false|false||CHRONICnull|chronic|Time|false|false||CHRONICnull|Hyponatremia|Disorder|false|false||Hyponatremianull|Has patient|Finding|false|false||patient hasnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Asymptomatic diagnosis of|Finding|false|false||asymptomatic
null|Asymptomatic (finding)|Finding|false|false||asymptomaticnull|Hyponatremia|Disorder|false|false||hyponatremianull|most likely|Finding|false|false||most likelynull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Hyponatremia|Disorder|false|false||hyponatremianull|Relate - vinyl resin|Drug|false|false||relatednull|Role Link Type - related|Finding|false|false||related
null|Related (finding)|Finding|false|false||relatednull|Definitely Related to Intervention|Modifier|false|false||related
null|Relationships|Modifier|false|false||relatednull|Liver diseases|Disorder|false|false||liver disease
null|Hepatobiliary Disorder|Disorder|false|false||liver diseasenull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Disease|Disorder|false|false||diseasenull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|aldosterone|Drug|false|false||aldosterone
null|aldosterone|Drug|false|false||aldosterone
null|aldosterone|Drug|false|false||aldosteronenull|Aldosterone measurement|Procedure|false|false||aldosteronenull|Fracture of second cervical vertebra|Disorder|false|false||axisnull|Axis vertebra|Anatomy|false|false||axisnull|Genus Axis|Entity|false|false||axisnull|Axis|Modifier|false|false||axisnull|DYSFUNCTION - SKIN DISORDERS|Disorder|false|false||dysfunctionnull|Dysfunction|Finding|false|false||dysfunction
null|physiopathological|Finding|false|false||dysfunction
null|Functional disorder|Finding|false|false||dysfunctionnull|Relate - vinyl resin|Drug|false|false||relatednull|Role Link Type - related|Finding|false|false||related
null|Related (finding)|Finding|false|false||relatednull|Definitely Related to Intervention|Modifier|false|false||related
null|Relationships|Modifier|false|false||relatednull|Liver diseases|Disorder|false|false||liver disease
null|Hepatobiliary Disorder|Disorder|false|false||liver diseasenull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Disease|Disorder|false|false||diseasenull|Asymptomatic diagnosis of|Finding|false|false||asymptomatic
null|Asymptomatic (finding)|Finding|false|false||asymptomaticnull|Hospitalization|Procedure|false|false||hospitalizationnull|furosemide|Drug|false|false||furosemide
null|furosemide|Drug|false|false||furosemidenull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Twice weekly|Time|false|false||twice weeklynull|Weekly|Time|false|false||weeklynull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|HIV Vaccine|Drug|false|false||HIV
null|HIV Vaccine|Drug|false|false||HIVnull|HIV Infections|Disorder|false|false||HIV
null|HIV|Disorder|false|false||HIVnull|Emtricitabine- and tenofovir-containing product|Drug|false|false||Emtricitabine-Tenofovir
null|Emtricitabine- and tenofovir-containing product|Drug|false|false||Emtricitabine-Tenofovirnull|emtricitabine|Drug|false|false||Emtricitabine
null|emtricitabine|Drug|false|false||Emtricitabinenull|tenofovir|Drug|false|false||Tenofovir
null|tenofovir|Drug|false|false||Tenofovirnull|Truvada|Drug|false|false||Truvada
null|Truvada|Drug|false|false||Truvadanull|raltegravir|Drug|false|false||Raltegravir
null|raltegravir|Drug|false|false||Raltegravirnull|In-House|Finding|false|false||in-housenull|House (environment)|Device|false|false||housenull|Home environment|Modifier|false|false||housenull|At discharge|Time|false|false||at dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|fluticasone|Drug|false|false||fluticasone
null|fluticasone|Drug|false|false||fluticasonenull|tiotropium|Drug|false|false||tiotropium
null|tiotropium|Drug|false|false||tiotropiumnull|albuterol|Drug|false|false||albuterol
null|albuterol|Drug|false|false||albuterolnull|In-House|Finding|false|false||in-housenull|House (environment)|Device|false|false||housenull|Home environment|Modifier|false|false||housenull|At discharge|Time|false|false||at dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Marketing basis - Transitional|Finding|false|false||TRANSITIONALnull|Transitional cell morphology|Modifier|false|false||TRANSITIONALnull|Peritoneal Fluid Culture|Procedure|false|false||peritoneal fluid culturenull|Peritoneal fluid (substance)|Finding|false|false||peritoneal fluidnull|Peritoneal fluid analysis|Procedure|false|false||peritoneal fluidnull|peritoneal|Anatomy|false|false||peritoneal
null|Peritoneum|Anatomy|false|false||peritonealnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Culture Dose Form|Drug|false|false||culturenull|Culture (Anthropological)|Finding|false|false||culture
null|Cultural aspects|Finding|false|false||culturenull|Microbial culture (procedure)|Procedure|false|false||culture
null|Laboratory culture|Procedure|false|false||culturenull|Query Status Code - new|Finding|false|false||New
null|Act Status - new|Finding|false|false||Newnull|Newar Language|Entity|false|false||Newnull|New|Modifier|false|false||Newnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|furosemide|Drug|false|false||Furosemide
null|furosemide|Drug|false|false||Furosemidenull|Daily|Time|false|false||dailynull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Hyperkalemia|Finding|false|false||hyperkalemia
null|Serum potassium level above reference range|Finding|false|false||hyperkalemianull|Hyponatremia|Disorder|false|false||hyponatremianull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Biweekly|Time|false|false||biweeklynull|Script|Finding|false|false||scriptnull|Once a week|Time|false|false||once weeklynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Weekly|Time|false|false||weeklynull|lab results|Finding|false|false||Lab resultsnull|AML Lab Table|Finding|false|false||Lab
null|LAT2 gene|Finding|false|false||Lab
null|EWS Lab Table|Finding|false|false||Labnull|Laboratory|Device|false|false||Labnull|Labrador retriever|Entity|false|false||Lab
null|Laboratory|Entity|false|false||Labnull|Send (transmission)|Finding|false|false||sentnull|conversation|Finding|false|false||conversationnull|Catheter placement|Procedure|false|false||catheter placementnull|null|Finding|false|false||catheternull|catheter device|Device|false|false||catheter
null|XXX>Catheter|Device|false|false||catheternull|null|Procedure|false|false||placement
null|Implantation procedure|Procedure|false|false||placement
null|Clinical act of insertion|Procedure|false|false||placementnull|Placement|Modifier|false|false||placementnull|CODE STATUS|Procedure|false|false||code statusnull|MDF Attribute Type - Code|Finding|false|false||code
null|A Codes|Finding|false|false||code
null|Code|Finding|false|false||codenull|Coding|Event|false|false||codenull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|Twice weekly|Time|false|false||twice weeklynull|Weekly|Time|false|false||weeklynull|Paracentesis|Procedure|false|false||paracentesesnull|MDF Attribute Type - Code|Finding|false|false||Code
null|A Codes|Finding|false|false||Code
null|Code|Finding|false|false||Codenull|Coding|Event|false|false||Codenull|Full|Modifier|false|false||fullnull|emergency contact|Finding|false|false||Emergency Contactnull|Consent Non-Disclosure Reason - Emergency|Finding|false|false||Emergency
null|Admission Type - Emergency|Finding|false|false||Emergency
null|Referral category - Emergency|Finding|false|false||Emergency
null|Emergencies [Disease/Finding]|Finding|false|false||Emergency
null|Consent Bypass Reason - Emergency|Finding|false|false||Emergency
null|Level of Care - Emergency|Finding|false|false||Emergency
null|Certification patient type - Emergency|Finding|false|false||Emergency
null|Encounter Admission Source - emergency|Finding|false|false||Emergency
null|Patient Class - Emergency|Finding|false|false||Emergency
null|Visit Priority Code - Emergency|Finding|false|false||Emergencynull|emergency encounter|Procedure|false|false||Emergencynull|Emergency Situation|Phenomenon|false|false||Emergencynull|Specialty Type - Emergency|Title|false|false||Emergencynull|Bale out|Time|false|false||Emergencynull|Contact - HL7 Attribution|Finding|false|false||Contact
null|Contact with|Finding|false|false||Contact
null|Communication Contact|Finding|false|false||Contactnull|contact person|Subject|false|false||Contactnull|Physical contact|Phenomenon|false|false||Contactnull|Personal Contact|Event|false|false||Contactnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Accurate (qualifier value)|Modifier|false|false||accuratenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|calcium carbonate|Drug|false|false||Calcium Carbonate
null|calcium carbonate|Drug|false|false||Calcium Carbonatenull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|carbonate ion|Drug|false|false||Carbonate
null|Carbonates|Drug|false|false||Carbonate
null|Carbonates|Drug|false|false||Carbonatenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Emtricitabine- and tenofovir-containing product|Drug|false|false||Emtricitabine-Tenofovir
null|Emtricitabine- and tenofovir-containing product|Drug|false|false||Emtricitabine-Tenofovirnull|emtricitabine|Drug|false|false||Emtricitabine
null|emtricitabine|Drug|false|false||Emtricitabinenull|tenofovir|Drug|false|false||Tenofovir
null|tenofovir|Drug|false|false||Tenofovirnull|Truvada|Drug|false|false||Truvada
null|Truvada|Drug|false|false||Truvadanull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|Daily|Time|false|false||DAILYnull|fluticasone propionate|Drug|false|false||Fluticasone Propionate
null|fluticasone propionate|Drug|false|false||Fluticasone Propionatenull|fluticasone|Drug|false|false||Fluticasone
null|fluticasone|Drug|false|false||Fluticasonenull|propionate|Drug|false|false||Propionate
null|Propionates|Drug|false|false||Propionatenull|Puff Dosing Unit|LabModifier|false|false||PUFF
null|Picofarad|LabModifier|false|false||PUFFnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|lactulose|Drug|false|false||Lactulose
null|lactulose|Drug|false|false||Lactulosenull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|raltegravir|Drug|false|false||Raltegravir
null|raltegravir|Drug|false|false||Raltegravirnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|rifaximin|Drug|false|false||Rifaximin
null|rifaximin|Drug|false|false||Rifaximinnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|tramadol|Drug|false|false||TraMADOL
null|tramadol|Drug|false|false||TraMADOLnull|Tramadol measurement (procedure)|Procedure|false|false||TraMADOLnull|Ultram|Drug|false|false||Ultram
null|Ultram|Drug|false|false||Ultramnull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|albuterol sulfate|Drug|false|false||albuterol sulfate
null|albuterol sulfate|Drug|false|false||albuterol sulfatenull|albuterol|Drug|false|false||albuterol
null|albuterol|Drug|false|false||albuterolnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfate
null|Sulfates, Inorganic|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfatenull|mcg/actuation|LabModifier|false|false||mcg/actuationnull|microgram|LabModifier|false|false||mcgnull|Actuation (unit of presentation)|LabModifier|false|false||actuationnull|Inhalation Route of Administration|Finding|false|false||inhalation
null|Inspiration (function)|Finding|false|false||inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||inhalationnull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Wheezing|Finding|false|false||Wheezingnull|tiotropium bromide|Drug|false|false||Tiotropium Bromide
null|tiotropium bromide|Drug|false|false||Tiotropium Bromidenull|tiotropium|Drug|false|false||Tiotropium
null|tiotropium|Drug|false|false||Tiotropiumnull|Bromides|Drug|false|false||Bromidenull|Bromides measurement|Procedure|false|false||Bromidenull|capsule (pharmacologic)|Drug|false|false||CAPnull|CATARACT, ANTERIOR POLAR|Disorder|false|false||CAPnull|BRD4 wt Allele|Finding|false|false||CAP
null|HACD1 gene|Finding|false|false||CAP
null|SERPINB6 gene|Finding|false|false||CAP
null|BRD4 gene|Finding|false|false||CAP
null|CAP1 gene|Finding|false|false||CAP
null|SORBS1 gene|Finding|false|false||CAP
null|LNPEP gene|Finding|false|false||CAPnull|CAP Regimen|Procedure|false|false||CAP
null|cisplatin/cyclophosphamide/doxorubicin protocol|Procedure|false|false||CAP
null|cyclophosphamide/doxorubicin/prednisone protocol|Procedure|false|false||CAPnull|Cap (physical object)|Device|false|false||CAP
null|Syringe Caps|Device|false|false||CAP
null|Cap device|Device|false|false||CAPnull|College of American Pathologists|Subject|false|false||CAPnull|Controlled Attenuation Parameter|Modifier|false|false||CAPnull|Capsule Dosing Unit|LabModifier|false|false||CAPnull|Daily|Time|false|false||DAILYnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|albuterol sulfate|Drug|false|false||albuterol sulfate
null|albuterol sulfate|Drug|false|false||albuterol sulfatenull|albuterol|Drug|false|false||albuterol
null|albuterol|Drug|false|false||albuterolnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfate
null|Sulfates, Inorganic|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfatenull|mcg/actuation|LabModifier|false|false||mcg/actuationnull|microgram|LabModifier|false|false||mcgnull|Actuation (unit of presentation)|LabModifier|false|false||actuationnull|Inhalation Route of Administration|Finding|false|false||inhalation
null|Inspiration (function)|Finding|false|false||inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||inhalationnull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Wheezing|Finding|false|false||Wheezingnull|calcium carbonate|Drug|false|false||Calcium Carbonate
null|calcium carbonate|Drug|false|false||Calcium Carbonatenull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|carbonate ion|Drug|false|false||Carbonate
null|Carbonates|Drug|false|false||Carbonate
null|Carbonates|Drug|false|false||Carbonatenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Emtricitabine- and tenofovir-containing product|Drug|false|false||Emtricitabine-Tenofovir
null|Emtricitabine- and tenofovir-containing product|Drug|false|false||Emtricitabine-Tenofovirnull|emtricitabine|Drug|false|false||Emtricitabine
null|emtricitabine|Drug|false|false||Emtricitabinenull|tenofovir|Drug|false|false||Tenofovir
null|tenofovir|Drug|false|false||Tenofovirnull|Truvada|Drug|false|false||Truvada
null|Truvada|Drug|false|false||Truvadanull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|Daily|Time|false|false||DAILYnull|fluticasone propionate|Drug|false|false||Fluticasone Propionate
null|fluticasone propionate|Drug|false|false||Fluticasone Propionatenull|fluticasone|Drug|false|false||Fluticasone
null|fluticasone|Drug|false|false||Fluticasonenull|propionate|Drug|false|false||Propionate
null|Propionates|Drug|false|false||Propionatenull|Puff Dosing Unit|LabModifier|false|false||PUFF
null|Picofarad|LabModifier|false|false||PUFFnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|lactulose|Drug|false|false||Lactulose
null|lactulose|Drug|false|false||Lactulosenull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|raltegravir|Drug|false|false||Raltegravir
null|raltegravir|Drug|false|false||Raltegravirnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|rifaximin|Drug|false|false||Rifaximin
null|rifaximin|Drug|false|false||Rifaximinnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|tiotropium bromide|Drug|false|false||Tiotropium Bromide
null|tiotropium bromide|Drug|false|false||Tiotropium Bromidenull|tiotropium|Drug|false|false||Tiotropium
null|tiotropium|Drug|false|false||Tiotropiumnull|Bromides|Drug|false|false||Bromidenull|Bromides measurement|Procedure|false|false||Bromidenull|capsule (pharmacologic)|Drug|false|false||CAPnull|CATARACT, ANTERIOR POLAR|Disorder|false|false||CAPnull|BRD4 wt Allele|Finding|false|false||CAP
null|HACD1 gene|Finding|false|false||CAP
null|SERPINB6 gene|Finding|false|false||CAP
null|BRD4 gene|Finding|false|false||CAP
null|CAP1 gene|Finding|false|false||CAP
null|SORBS1 gene|Finding|false|false||CAP
null|LNPEP gene|Finding|false|false||CAPnull|CAP Regimen|Procedure|false|false||CAP
null|cisplatin/cyclophosphamide/doxorubicin protocol|Procedure|false|false||CAP
null|cyclophosphamide/doxorubicin/prednisone protocol|Procedure|false|false||CAPnull|Cap (physical object)|Device|false|false||CAP
null|Syringe Caps|Device|false|false||CAP
null|Cap device|Device|false|false||CAPnull|College of American Pathologists|Subject|false|false||CAPnull|Controlled Attenuation Parameter|Modifier|false|false||CAPnull|Capsule Dosing Unit|LabModifier|false|false||CAPnull|Daily|Time|false|false||DAILYnull|tramadol|Drug|false|false||TraMADOL
null|tramadol|Drug|false|false||TraMADOLnull|Tramadol measurement (procedure)|Procedure|false|false||TraMADOLnull|Ultram|Drug|false|false||Ultram
null|Ultram|Drug|false|false||Ultramnull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|furosemide|Drug|false|false||Furosemide
null|furosemide|Drug|false|false||Furosemidenull|Daily|Time|false|false||DAILYnull|furosemide|Drug|false|false||furosemide
null|furosemide|Drug|false|false||furosemidenull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Daily|Time|false|false||dailynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|Referral category - Outpatient|Finding|false|false||Outpatient
null|Patient Class - Outpatient|Finding|false|false||Outpatientnull|Outpatients|Subject|false|false||Outpatientnull|AML Lab Table|Finding|false|false||Lab
null|LAT2 gene|Finding|false|false||Lab
null|EWS Lab Table|Finding|false|false||Labnull|Laboratory|Device|false|false||Labnull|Labrador retriever|Entity|false|false||Lab
null|Laboratory|Entity|false|false||Labnull|Work|Event|false|false||Worknull|Biweekly|Time|false|false||biweeklynull|Bone Morphogenetic Proteins|Drug|false|false||BMP
null|Bone Morphogenetic Proteins|Drug|false|false||BMPnull|carmustine/methotrexate/procarbazine protocol|Procedure|false|false||BMPnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|hepatitis C virus|Disorder|false|false||HCV
null|Hepatitis C|Disorder|false|false||HCVnull|Liver Cirrhosis|Disorder|false|false||cirrhosis
null|Cirrhosis|Disorder|false|false||cirrhosisnull|Hyperkalemia|Finding|false|false||Hyperkalemia
null|Serum potassium level above reference range|Finding|false|false||Hyperkalemianull|Neoplasm Metastasis|Disorder|false|false||SECONDARYnull|metastatic qualifier|Finding|false|false||SECONDARYnull|Secondary to|Modifier|false|false||SECONDARYnull|second (number)|LabModifier|false|false||SECONDARYnull|Diagnosis|Procedure|false|false||DIAGNOSESnull|HIV Vaccine|Drug|false|false||HIV
null|HIV Vaccine|Drug|false|false||HIVnull|HIV Infections|Disorder|false|false||HIV
null|HIV|Disorder|false|false||HIVnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Hyponatremia|Disorder|false|false||Hyponatremianull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|FBXW7-AS1 gene|Finding|false|false||Dearnull|Production Class Code - Pleasure|Finding|false|false||pleasure
null|pleasurable emotion|Finding|false|false||pleasurenull|Pleasure - Animals raised for recreation|Entity|false|false||pleasurenull|Abdominal Pain|Finding|false|false||abdominal painnull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Malignant neoplasm of abdomen|Disorder|false|false||abdomennull|Abdomen problem|Finding|false|false||abdomennull|Abdomen|Anatomy|false|false||abdomen
null|Abdominal Cavity|Anatomy|false|false||abdomennull|Liver Cirrhosis|Disorder|false|false||cirrhosis
null|Cirrhosis|Disorder|false|false||cirrhosisnull|Paracentesis|Procedure|false|false||paracentesisnull|Much|Finding|false|false||muchnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Potassium increased|Finding|false|false||high potassiumnull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Potassium Drug Class|Drug|false|false||potassium
null|Dietary Potassium|Drug|false|false||potassium
null|potassium|Drug|false|false||potassium
null|potassium|Drug|false|false||potassium
null|potassium|Drug|false|false||potassium
null|Potassium supplement|Drug|false|false||potassium
null|Potassium supplement|Drug|false|false||potassiumnull|Potassium metabolic function|Finding|false|false||potassiumnull|Potassium measurement|Procedure|false|false||potassiumnull|Hospitalization|Procedure|false|false||hospitalizationnull|CAME|Drug|false|false||camenull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|desire|Finding|false|false||desirenull|Representation (action)|Event|false|false||representativenull|Hospice Care|Procedure|false|false||hospicenull|Hospice (environment)|Device|false|false||hospicenull|Hospice (environment)|Entity|false|false||hospicenull|Paracentesis|Procedure|false|false||paracentesesnull|Catheter placement|Procedure|false|false||catheter placementnull|null|Finding|false|false||catheternull|catheter device|Device|false|false||catheter
null|XXX>Catheter|Device|false|false||catheternull|null|Procedure|false|false||placement
null|Implantation procedure|Procedure|false|false||placement
null|Clinical act of insertion|Procedure|false|false||placementnull|Placement|Modifier|false|false||placementnull|Hospice Care|Procedure|false|false||hospicenull|Hospice (environment)|Device|false|false||hospicenull|Hospice (environment)|Entity|false|false||hospicenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Hospice Care|Procedure|false|false||hospicenull|Hospice (environment)|Device|false|false||hospicenull|Hospice (environment)|Entity|false|false||hospicenull|Vitelliform Macular Dystrophy|Disorder|false|false||bestnull|BEST1 wt Allele|Finding|false|false||best
null|BEST1 gene|Finding|false|false||bestnull|best (quality)|Modifier|false|false||bestnull|Care team|Finding|false|false||care teamnull|null|Attribute|false|false||care teamnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Team|Subject|false|false||teamnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions