 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|44,53|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|44,53|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|44,58|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|78,87|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|78,87|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|78,87|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|78,87|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|78,87|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|78,92|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|110,115|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|110,115|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|110,115|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|134,137|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|134,137|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|134,137|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|134,137|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|134,137|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|145,152|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|145,152|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|SIMPLE_SEGMENT|154,166|true|false|false|||NEUROSURGERY
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|154,166|true|false|false|C0524850|Neurosurgical Procedures|NEUROSURGERY
Finding|Body Substance|Allergies|181,188|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Allergies|181,188|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Allergies|181,188|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Allergies|189,197|true|false|false|||recorded
Attribute|Clinical Attribute|Allergies|217,226|true|false|false|C1717415||Allergies
Event|Event|Allergies|217,226|true|false|false|||Allergies
Finding|Pathologic Function|Allergies|217,226|true|false|false|C0020517|Hypersensitivity|Allergies
Drug|Pharmacologic Substance|Allergies|230,235|true|false|false|C0013227|Pharmaceutical Preparations|Drugs
Event|Event|Allergies|230,235|true|false|false|||Drugs
Procedure|Therapeutic or Preventive Procedure|Allergies|230,235|true|false|false|C3687832|Drugs - dental services|Drugs
Event|Event|Allergies|238,247|true|false|false|||Attending
Finding|Functional Concept|Allergies|238,247|true|false|false|C1999232|Attending (action)|Attending
Finding|Finding|Chief Complaint|273,277|false|false|false|C0016928|Gait|Gait
Finding|Finding|Chief Complaint|273,289|false|false|false|C0231686|Gait, Unsteady|Gait instability
Event|Event|Chief Complaint|278,289|false|false|false|||instability
Finding|Finding|Chief Complaint|278,289|false|false|false|C1444783|Instability|instability
Finding|Finding|Chief Complaint|291,305|false|false|false|C0743800|multiple falls|multiple falls
Disorder|Injury or Poisoning|Chief Complaint|300,305|false|false|false|C0000921|Accidental Falls|falls
Event|Event|Chief Complaint|300,305|false|false|false|||falls
Finding|Finding|Chief Complaint|300,305|false|false|false|C0085639|Falls|falls
Finding|Classification|Chief Complaint|308,313|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|314,322|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|314,322|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|326,344|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|335,344|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|335,344|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|335,344|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|335,344|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|335,344|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|History of Present Illness|394,402|false|false|false|||pleasant
Finding|Mental Process|History of Present Illness|394,402|false|false|false|C2987187|Pleasant|pleasant
Finding|Functional Concept|History of Present Illness|403,408|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|403,415|false|false|false|C0230370|Structure of right hand|right handed
Finding|Idea or Concept|History of Present Illness|420,424|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|History of Present Illness|420,424|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|History of Present Illness|429,433|false|false|false|||male
Finding|Finding|History of Present Illness|429,433|false|false|false|C1706180|Male Gender|male
Disorder|Disease or Syndrome|History of Present Illness|439,443|false|false|false|C0004238|Atrial Fibrillation|Afib
Lab|Laboratory or Test Result|History of Present Illness|439,443|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Afib
Drug|Organic Chemical|History of Present Illness|449,457|false|false|false|C0699129|Coumadin|coumadin
Drug|Pharmacologic Substance|History of Present Illness|449,457|false|false|false|C0699129|Coumadin|coumadin
Event|Event|History of Present Illness|449,457|false|false|false|||coumadin
Event|Event|History of Present Illness|472,483|false|false|false|||independent
Finding|Finding|History of Present Illness|472,483|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|independent
Finding|Idea or Concept|History of Present Illness|472,483|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|independent
Event|Event|History of Present Illness|485,491|false|false|false|||living
Finding|Idea or Concept|History of Present Illness|520,524|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Event|Event|History of Present Illness|525,530|false|false|false|||state
Finding|Functional Concept|History of Present Illness|525,530|false|false|false|C1442792|State|state
Finding|Finding|History of Present Illness|525,540|false|false|false|C0683314|personal health|state of health
Event|Event|History of Present Illness|534,540|false|false|false|||health
Finding|Idea or Concept|History of Present Illness|534,540|false|false|false|C0018684|Health|health
Finding|Idea or Concept|History of Present Illness|556,560|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|History of Present Illness|556,560|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Finding|History of Present Illness|570,574|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|History of Present Illness|570,574|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|History of Present Illness|570,574|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|History of Present Illness|585,592|false|false|false|||reports
Event|Event|History of Present Illness|601,606|false|false|false|||began
Event|Event|History of Present Illness|614,621|false|false|false|||periods
Finding|Organism Function|History of Present Illness|614,621|false|false|false|C0025344|Menstruation|periods
Event|Event|History of Present Illness|625,637|false|false|false|||disorganized
Event|Event|History of Present Illness|639,645|false|false|false|||speech
Finding|Organism Function|History of Present Illness|639,645|false|false|false|C0037817|Speech|speech
Procedure|Diagnostic Procedure|History of Present Illness|639,645|false|false|false|C0846595|Speech assessment|speech
Finding|Finding|History of Present Illness|650,654|false|false|false|C0016928|Gait|gait
Finding|Finding|History of Present Illness|650,666|false|false|false|C0231686|Gait, Unsteady|gait instability
Event|Event|History of Present Illness|655,666|false|false|false|||instability
Finding|Finding|History of Present Illness|655,666|false|false|false|C1444783|Instability|instability
Finding|Finding|History of Present Illness|684,690|true|false|false|C1561668|History of fall|a fall
Event|Event|History of Present Illness|686,690|true|false|false|||fall
Finding|Finding|History of Present Illness|686,690|true|true|false|C0085639|Falls|fall
Finding|Gene or Genome|History of Present Illness|707,710|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|History of Present Illness|719,724|false|false|false|||broke
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|733,737|false|false|false|C0035561|Bone structure of rib|ribs
Drug|Food|History of Present Illness|745,751|false|false|false|C0009237|Coffee|coffee
Event|Event|History of Present Illness|752,757|false|false|false|||table
Finding|Intellectual Product|History of Present Illness|752,757|false|false|false|C1706074|Data Table|table
Anatomy|Body Location or Region|History of Present Illness|780,784|true|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|780,784|true|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|History of Present Illness|780,784|true|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|780,784|true|false|false|C0876917|Procedure on head|head
Disorder|Injury or Poisoning|History of Present Illness|780,791|true|false|false|C0018674|Craniocerebral Trauma|head trauma
Disorder|Injury or Poisoning|History of Present Illness|785,791|true|false|false|C1368081;C3263723;C3714660|Physical trauma;Trauma;Traumatic injury|trauma
Event|Event|History of Present Illness|785,791|true|false|false|||trauma
Procedure|Health Care Activity|History of Present Illness|785,791|true|false|false|C0548346|Trauma assessment and care|trauma
Event|Event|History of Present Illness|804,811|true|false|false|||scanned
Event|Event|History of Present Illness|818,821|true|false|false|||OSH
Event|Event|History of Present Illness|836,842|false|false|false|||speech
Finding|Organism Function|History of Present Illness|836,842|false|false|false|C0037817|Speech|speech
Procedure|Diagnostic Procedure|History of Present Illness|836,842|false|false|false|C0846595|Speech assessment|speech
Event|Event|History of Present Illness|847,859|false|false|false|||unsteadiness
Finding|Finding|History of Present Illness|847,859|false|false|false|C0427108|General unsteadiness|unsteadiness
Event|Event|History of Present Illness|865,870|false|false|false|||waxed
Event|Event|History of Present Illness|875,880|false|false|false|||waned
Event|Event|History of Present Illness|918,925|false|false|false|||reports
Finding|Finding|History of Present Illness|940,944|false|false|false|C4281574|Much|much
Event|Event|History of Present Illness|945,953|false|false|false|||improved
Event|Event|History of Present Illness|963,968|false|false|false|||takes
Drug|Pharmacologic Substance|History of Present Illness|973,982|false|false|false|C0012798|Diuretics|diuretics
Event|Event|History of Present Illness|973,982|false|false|false|||diuretics
Event|Event|History of Present Illness|994,1000|false|false|false|||period
Finding|Organism Function|History of Present Illness|994,1000|false|false|false|C0025344|Menstruation|period
Procedure|Research Activity|History of Present Illness|994,1000|false|false|false|C2347804|Clinical Trial Period|period
Event|Event|History of Present Illness|1008,1012|false|false|false|||lost
Event|Event|History of Present Illness|1018,1021|false|false|false|||lbs
Procedure|Laboratory Procedure|History of Present Illness|1018,1021|false|false|false|C3161851|liquid-based cytology (procedure)|lbs
Event|Event|History of Present Illness|1042,1049|false|false|false|||sorting
Event|Event|History of Present Illness|1050,1056|false|false|false|||papers
Finding|Intellectual Product|History of Present Illness|1076,1081|false|false|false|C1706074|Data Table|table
Event|Event|History of Present Illness|1091,1095|false|false|false|||fell
Event|Event|History of Present Illness|1101,1109|false|false|false|||standing
Event|Event|History of Present Illness|1125,1134|false|false|false|||dizziness
Finding|Sign or Symptom|History of Present Illness|1125,1134|false|false|false|C0012833;C0042571|Dizziness;Vertigo|dizziness
Event|Event|History of Present Illness|1139,1146|true|false|false|||reports
Event|Event|History of Present Illness|1151,1154|true|false|false|||LOC
Anatomy|Body Location or Region|History of Present Illness|1159,1163|true|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1159,1163|true|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|History of Present Illness|1159,1163|true|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1159,1163|true|false|false|C0876917|Procedure on head|head
Disorder|Injury or Poisoning|History of Present Illness|1159,1170|true|false|false|C0018674|Craniocerebral Trauma|head trauma
Disorder|Injury or Poisoning|History of Present Illness|1164,1170|true|false|false|C1368081;C3263723;C3714660|Physical trauma;Trauma;Traumatic injury|trauma
Event|Event|History of Present Illness|1164,1170|true|false|false|||trauma
Procedure|Health Care Activity|History of Present Illness|1164,1170|true|false|false|C0548346|Trauma assessment and care|trauma
Event|Event|History of Present Illness|1179,1183|true|false|false|||able
Finding|Finding|History of Present Illness|1179,1183|true|false|false|C1299581|Able (qualifier value)|able
Event|Event|History of Present Illness|1187,1192|true|false|false|||stand
Event|Event|History of Present Illness|1198,1200|false|false|false|||up
Event|Event|History of Present Illness|1205,1213|false|false|false|||continue
Finding|Idea or Concept|History of Present Illness|1205,1213|false|false|false|C0549178|Continuous|continue
Event|Event|History of Present Illness|1219,1223|false|false|false|||work
Event|Occupational Activity|History of Present Illness|1219,1223|false|false|false|C0043227|Work|work
Event|Event|History of Present Illness|1234,1240|false|false|false|||placed
Event|Event|History of Present Illness|1266,1269|false|false|false|||got
Event|Event|History of Present Illness|1283,1287|false|false|false|||fell
Event|Event|History of Present Illness|1315,1321|true|false|false|||denies
Event|Event|History of Present Illness|1326,1329|true|false|false|||LOC
Anatomy|Body Location or Region|History of Present Illness|1333,1337|true|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1333,1337|true|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|History of Present Illness|1333,1337|true|false|false|C0362076|Problems with head|head
Event|Event|History of Present Illness|1333,1337|true|false|false|||head
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1333,1337|true|false|false|C0876917|Procedure on head|head
Disorder|Injury or Poisoning|History of Present Illness|1339,1345|true|false|false|C1368081;C3263723;C3714660|Physical trauma;Trauma;Traumatic injury|trauma
Event|Event|History of Present Illness|1339,1345|true|false|false|||trauma
Procedure|Health Care Activity|History of Present Illness|1339,1345|true|false|false|C0548346|Trauma assessment and care|trauma
Event|Event|History of Present Illness|1347,1354|true|false|false|||blaming
Event|Event|History of Present Illness|1359,1370|false|false|false|||instability
Finding|Finding|History of Present Illness|1359,1370|false|false|false|C1444783|Instability|instability
Event|Event|History of Present Illness|1379,1387|false|false|false|||weakness
Finding|Sign or Symptom|History of Present Illness|1379,1387|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1400,1406|true|false|false|C0040408|Tongue|tongue
Disorder|Neoplastic Process|History of Present Illness|1400,1406|true|false|false|C0153933|Benign neoplasm of tongue|tongue
Event|Event|History of Present Illness|1400,1406|true|false|false|||tongue
Procedure|Health Care Activity|History of Present Illness|1400,1406|true|false|false|C0872394|Procedure on tongue|tongue
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|1400,1413|true|false|false|C0241424|Tongue biting|tongue biting
Disorder|Injury or Poisoning|History of Present Illness|1407,1413|true|false|false|C0005658|bite injury|biting
Event|Event|History of Present Illness|1407,1413|true|false|false|||biting
Finding|Physiologic Function|History of Present Illness|1407,1413|true|false|false|C2584293|Biting|biting
Event|Event|History of Present Illness|1417,1421|true|false|false|||loss
Finding|Finding|History of Present Illness|1417,1421|true|false|false|C5890125|Loss (adaptation)|loss
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1425,1430|true|false|false|C0021853|Intestines|bowel
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1431,1438|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|History of Present Illness|1431,1438|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1431,1438|false|false|false|C0872388|Procedures on bladder|bladder
Finding|Finding|History of Present Illness|1431,1449|false|false|false|C0876938;C4319531|Bladder Continence Question;Urinary bladder control|bladder continence
Finding|Intellectual Product|History of Present Illness|1431,1449|false|false|false|C0876938;C4319531|Bladder Continence Question;Urinary bladder control|bladder continence
Event|Event|History of Present Illness|1439,1449|false|false|false|||continence
Disorder|Disease or Syndrome|History of Present Illness|1463,1466|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Event|Event|History of Present Illness|1463,1466|false|false|false|||bed
Finding|Intellectual Product|History of Present Illness|1463,1466|false|false|false|C2346952|Bachelor of Education|bed
Event|Event|History of Present Illness|1498,1510|false|false|false|||presentation
Finding|Idea or Concept|History of Present Illness|1498,1510|false|false|false|C0449450|Presentation|presentation
Event|Event|History of Present Illness|1525,1534|false|false|false|||concerned
Disorder|Injury or Poisoning|History of Present Illness|1545,1550|false|false|false|C0000921|Accidental Falls|falls
Event|Event|History of Present Illness|1545,1550|false|false|false|||falls
Finding|Finding|History of Present Illness|1545,1550|false|false|false|C0085639|Falls|falls
Event|Event|History of Present Illness|1555,1562|false|false|false|||brought
Attribute|Clinical Attribute|History of Present Illness|1594,1603|false|false|false|C0945731||diagnosis
Event|Event|History of Present Illness|1594,1603|false|false|false|||diagnosis
Finding|Classification|History of Present Illness|1594,1603|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|History of Present Illness|1594,1603|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|History of Present Illness|1594,1603|false|false|false|C0011900|Diagnosis|diagnosis
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1607,1612|false|false|false|C0378717|elongation factor DmS-II|DM II
Finding|Idea or Concept|History of Present Illness|1630,1635|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|History of Present Illness|1630,1635|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Gene or Genome|History of Present Illness|1636,1639|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|History of Present Illness|1649,1656|false|false|false|||started
Anatomy|Body Space or Junction|History of Present Illness|1657,1661|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|History of Present Illness|1657,1661|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|History of Present Illness|1657,1661|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|History of Present Illness|1657,1661|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Pharmacologic Substance|History of Present Illness|1657,1675|false|false|false|C0359086|Oral hypoglycemic|oral hypoglycemics
Drug|Pharmacologic Substance|History of Present Illness|1662,1675|false|false|false|C0020616|Hypoglycemic Agents|hypoglycemics
Event|Event|History of Present Illness|1662,1675|false|false|false|||hypoglycemics
Event|Event|History of Present Illness|1689,1696|false|false|false|||reports
Finding|Finding|History of Present Illness|1704,1707|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|History of Present Illness|1704,1707|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Event|Event|History of Present Illness|1716,1720|false|false|false|||home
Finding|Idea or Concept|History of Present Illness|1716,1720|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|History of Present Illness|1716,1720|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|History of Present Illness|1716,1720|false|false|false|C1553498|home health encounter|home
Event|Event|History of Present Illness|1729,1733|false|false|false|||seen
Finding|Intellectual Product|History of Present Illness|1764,1768|false|false|false|C1561540|Transaction counts and value totals - week|week
Attribute|Clinical Attribute|History of Present Illness|1794,1801|false|false|false|C0881943||CT head
Procedure|Diagnostic Procedure|History of Present Illness|1794,1801|false|false|false|C0202691|CAT scan of head|CT head
Anatomy|Body Location or Region|History of Present Illness|1797,1801|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1797,1801|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|History of Present Illness|1797,1801|false|false|false|C0362076|Problems with head|head
Event|Event|History of Present Illness|1797,1801|false|false|false|||head
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1797,1801|false|false|false|C0876917|Procedure on head|head
Event|Event|History of Present Illness|1808,1817|false|false|false|||completed
Finding|Intellectual Product|History of Present Illness|1832,1836|false|false|false|C1561540|Transaction counts and value totals - week|week
Anatomy|Body Location or Region|History of Present Illness|1853,1857|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1853,1857|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|History of Present Illness|1853,1857|false|false|false|C0362076|Problems with head|head
Event|Event|History of Present Illness|1853,1857|false|false|false|||head
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1853,1857|false|false|false|C0876917|Procedure on head|head
Event|Event|History of Present Illness|1862,1869|false|false|false|||scanned
Event|Event|History of Present Illness|1876,1884|true|false|false|||revealed
Event|Event|History of Present Illness|1888,1893|true|false|false|||bleed
Finding|Pathologic Function|History of Present Illness|1888,1893|true|false|false|C0019080|Hemorrhage|bleed
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1907,1919|false|false|false|C0016733|frontal lobe|frontal lobe
Disorder|Neoplastic Process|History of Present Illness|1907,1919|false|false|false|C0153635|malignant neoplasm of frontal lobe|frontal lobe
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1915,1919|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|History of Present Illness|1915,1919|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Event|Event|History of Present Illness|1932,1936|false|false|false|||mass
Finding|Finding|History of Present Illness|1932,1936|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|History of Present Illness|1932,1936|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|History of Present Illness|1932,1936|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Anatomy|Cell Component|History of Present Illness|1968,1975|true|false|false|C1660780|midline cell component|midline
Finding|Finding|History of Present Illness|1968,1981|true|false|false|C4086580|Midline Shift|midline shift
Event|Event|History of Present Illness|1976,1981|true|false|false|||shift
Finding|Functional Concept|History of Present Illness|1976,1981|true|false|false|C0333051|shift displacement|shift
Phenomenon|Phenomenon or Process|History of Present Illness|1976,1981|true|false|false|C2347509|Physical Shift|shift
Event|Event|History of Present Illness|1983,1995|false|false|false|||Neurosurgery
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1983,1995|false|false|false|C0524850|Neurosurgical Procedures|Neurosurgery
Event|Event|History of Present Illness|2000,2009|false|false|false|||contacted
Event|Event|History of Present Illness|2014,2024|false|false|false|||evaluation
Finding|Idea or Concept|History of Present Illness|2014,2024|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|History of Present Illness|2014,2024|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Event|Event|History of Present Illness|2033,2037|false|false|false|||mass
Finding|Finding|History of Present Illness|2033,2037|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|History of Present Illness|2033,2037|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|History of Present Illness|2033,2037|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Finding|History of Present Illness|2046,2054|false|false|false|C0332149|Possible|possible
Attribute|Clinical Attribute|History of Present Illness|2055,2059|false|false|false|C5890809||role
Event|Event|History of Present Illness|2055,2059|false|false|false|||role
Finding|Conceptual Entity|History of Present Illness|2055,2059|false|false|false|C0035820;C1704326;C1705809;C1705811;C1705812;C3871154|NCI Thesaurus Role;Role;Security Role Object;Social Role;Terminology Role Entity;role - RoleClass|role
Finding|Intellectual Product|History of Present Illness|2055,2059|false|false|false|C0035820;C1704326;C1705809;C1705811;C1705812;C3871154|NCI Thesaurus Role;Role;Security Role Object;Social Role;Terminology Role Entity;role - RoleClass|role
Finding|Social Behavior|History of Present Illness|2055,2059|false|false|false|C0035820;C1704326;C1705809;C1705811;C1705812;C3871154|NCI Thesaurus Role;Role;Security Role Object;Social Role;Terminology Role Entity;role - RoleClass|role
Finding|Body Substance|History of Present Illness|2067,2074|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|2067,2074|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|2067,2074|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|2084,2092|false|false|false|||symptoms
Finding|Functional Concept|History of Present Illness|2084,2092|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|History of Present Illness|2084,2092|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Drug|Amino Acid, Peptide, or Protein|Past Medical History|2120,2125|false|false|false|C0378717|elongation factor DmS-II|DM II
Disorder|Disease or Syndrome|Past Medical History|2127,2130|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|Past Medical History|2127,2130|false|false|false|||HTN
Drug|Organic Chemical|Past Medical History|2156,2164|false|false|false|C0699129|Coumadin|coumadin
Drug|Pharmacologic Substance|Past Medical History|2156,2164|false|false|false|C0699129|Coumadin|coumadin
Event|Event|Past Medical History|2156,2164|false|false|false|||coumadin
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2166,2174|false|false|false|C0033572;C4266527|Prostate;Structure of prostate (body structure)|prostate
Disorder|Disease or Syndrome|Past Medical History|2166,2174|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|prostate
Disorder|Neoplastic Process|Past Medical History|2166,2174|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|prostate
Disorder|Neoplastic Process|Past Medical History|2166,2177|false|false|false|C0376358|Malignant neoplasm of prostate|prostate CA
Event|Event|Past Medical History|2175,2177|false|false|false|||CA
Event|Event|Past Medical History|2179,2186|false|false|false|||treated
Finding|Finding|General Exam|2277,2289|false|false|false|C4533677|at admission|At Admission
Event|Event|General Exam|2280,2289|false|false|false|||Admission
Procedure|Health Care Activity|General Exam|2280,2289|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Event|Event|General Exam|2293,2296|false|false|false|||Gen
Finding|Classification|General Exam|2293,2296|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Finding|Gene or Genome|General Exam|2293,2296|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Event|Event|General Exam|2305,2316|false|false|false|||comfortable
Finding|Finding|General Exam|2305,2316|false|false|false|C5546696|Feeling comfortable|comfortable
Disorder|Disease or Syndrome|General Exam|2318,2321|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|2318,2321|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|2318,2321|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|2318,2321|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|2318,2321|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|General Exam|2318,2321|false|false|false|||NAD
Finding|Finding|General Exam|2318,2321|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|General Exam|2323,2328|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|General Exam|2330,2336|false|false|false|C0034121|Pupil|Pupils
Event|Event|General Exam|2346,2350|false|false|false|||EOMs
Finding|Functional Concept|General Exam|2346,2350|false|false|false|C0241886|Extraocular|EOMs
Event|Event|General Exam|2351,2357|false|false|false|||intact
Finding|Finding|General Exam|2351,2357|false|false|false|C1554187|Gender Status - Intact|intact
Anatomy|Body Part, Organ, or Organ Component|General Exam|2362,2367|false|false|false|C0024109|Lung|Lungs
Drug|Amino Acid, Peptide, or Protein|General Exam|2369,2372|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|General Exam|2369,2372|false|false|false|||CTA
Finding|Gene or Genome|General Exam|2369,2372|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|General Exam|2369,2372|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Anatomy|Body Part, Organ, or Organ Component|General Exam|2386,2393|false|false|false|C0018787|Heart|Cardiac
Finding|Intellectual Product|General Exam|2386,2393|false|false|false|C1314974|Cardiac attachment|Cardiac
Finding|Finding|General Exam|2416,2435|false|false|false|C0232258|Pansystolic murmur|holosystolic murmur
Event|Event|General Exam|2429,2435|false|false|false|||murmur
Finding|Finding|General Exam|2429,2435|false|false|false|C0018808|Heart murmur|murmur
Anatomy|Body Location or Region|General Exam|2437,2440|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|Abd
Disorder|Cell or Molecular Dysfunction|General Exam|2437,2440|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|Abd
Disorder|Disease or Syndrome|General Exam|2442,2446|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|General Exam|2442,2446|false|false|false|||Soft
Event|Event|General Exam|2448,2450|false|false|false|||NT
Event|Event|General Exam|2464,2468|false|false|false|||Warm
Finding|Finding|General Exam|2464,2468|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|2464,2468|false|false|false|C0687712|warming process|Warm
Finding|Finding|General Exam|2473,2477|false|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|2478,2486|false|false|false|||perfused
Finding|Mental Process|General Exam|2495,2501|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|General Exam|2495,2508|false|false|false|C0488568;C0488569||Mental status
Finding|Finding|General Exam|2495,2508|false|false|false|C0278060|Mental state|Mental status
Attribute|Clinical Attribute|General Exam|2502,2508|false|false|false|C5889824||status
Event|Event|General Exam|2502,2508|false|false|false|||status
Finding|Idea or Concept|General Exam|2502,2508|false|false|false|C1546481|What subject filter - Status|status
Event|Event|General Exam|2510,2515|false|false|false|||Awake
Finding|Finding|General Exam|2510,2515|false|false|false|C0234422|Awake (finding)|Awake
Event|Event|General Exam|2520,2531|false|false|false|||cooperative
Event|Event|General Exam|2537,2541|false|false|false|||exam
Finding|Functional Concept|General Exam|2537,2541|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|General Exam|2537,2541|false|false|false|C0582103|Medical Examination|exam
Event|Event|General Exam|2550,2556|false|false|false|||affect
Finding|Mental Process|General Exam|2550,2556|false|false|false|C0001721|Affect (mental function)|affect
Procedure|Health Care Activity|General Exam|2550,2556|false|false|false|C2237113|assessment of affect|affect
Event|Event|General Exam|2558,2569|false|false|false|||Orientation
Finding|Mental Process|General Exam|2558,2569|false|false|false|C0029266|Mental Orientation|Orientation
Event|Event|General Exam|2571,2579|false|false|false|||Oriented
Finding|Finding|General Exam|2571,2579|false|false|false|C1961028|Oriented to place|Oriented
Finding|Finding|General Exam|2571,2589|false|false|false|C1961030|Oriented to person|Oriented to person
Attribute|Clinical Attribute|General Exam|2583,2589|false|false|false|C5890614||person
Event|Event|General Exam|2583,2589|false|false|false|||person
Finding|Intellectual Product|General Exam|2583,2589|false|false|false|C1522390|Person Info|person
Event|Activity|General Exam|2591,2596|false|false|false|C1882509|put - instruction imperative|place
Event|Event|General Exam|2591,2596|false|false|false|||place
Finding|Functional Concept|General Exam|2591,2596|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|General Exam|2591,2596|false|false|false|C1533810||place
Event|Event|General Exam|2608,2614|false|false|false|||Recall
Event|Governmental or Regulatory Activity|General Exam|2608,2614|false|false|false|C1705180|Recall (activity)|Recall
Finding|Mental Process|General Exam|2608,2614|false|false|false|C0034770|Mental Recall|Recall
Event|Event|General Exam|2620,2627|false|false|false|||objects
Procedure|Therapeutic or Preventive Procedure|General Exam|2631,2640|false|false|false|C0886384|5 minutes Office visit|5 minutes
Event|Event|General Exam|2633,2640|false|false|false|||minutes
Attribute|Clinical Attribute|General Exam|2642,2650|false|false|false|C2706915||Language
Event|Event|General Exam|2642,2650|false|false|false|||Language
Finding|Intellectual Product|General Exam|2642,2650|false|false|false|C0033348|Programming Languages|Language
Event|Event|General Exam|2652,2658|false|false|false|||Speech
Finding|Organism Function|General Exam|2652,2658|false|false|false|C0037817|Speech|Speech
Procedure|Diagnostic Procedure|General Exam|2652,2658|false|false|false|C0846595|Speech assessment|Speech
Event|Event|General Exam|2662,2668|false|false|false|||fluent
Finding|Idea or Concept|General Exam|2670,2674|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Event|Event|General Exam|2675,2688|false|false|false|||comprehension
Finding|Mental Process|General Exam|2675,2688|false|false|false|C0162340|Comprehension|comprehension
Event|Event|General Exam|2690,2700|false|false|false|||Difficulty
Finding|Finding|General Exam|2690,2700|false|false|false|C1299586|Has difficulty doing (qualifier value)|Difficulty
Finding|Finding|General Exam|2690,2705|false|false|false|C0332218|Difficult (qualifier value)|Difficulty with
Event|Event|General Exam|2706,2716|false|false|false|||repitition
Event|Event|General Exam|2718,2724|false|false|false|||Naming
Finding|Mental Process|General Exam|2718,2724|false|false|false|C0233735|Naming (function)|Naming
Event|Event|General Exam|2725,2731|false|false|false|||intact
Finding|Finding|General Exam|2725,2731|false|false|false|C1554187|Gender Status - Intact|intact
Disorder|Mental or Behavioral Dysfunction|General Exam|2736,2746|true|false|false|C0013362|Dysarthria|dysarthria
Event|Event|General Exam|2736,2746|true|false|false|||dysarthria
Event|Event|General Exam|2761,2767|true|false|false|||errors
Anatomy|Body Part, Organ, or Organ Component|General Exam|2770,2777|false|false|false|C0037303|Bone structure of cranium|Cranial
Anatomy|Body Part, Organ, or Organ Component|General Exam|2770,2784|false|false|false|C0010268|Cranial Nerves|Cranial Nerves
Disorder|Neoplastic Process|General Exam|2770,2784|false|false|false|C0004992;C0496937|Benign neoplasm of cranial nerves;Neoplasm of uncertain or unknown behavior of cranial nerves|Cranial Nerves
Anatomy|Body Part, Organ, or Organ Component|General Exam|2778,2784|false|false|false|C0027740|Nerve|Nerves
Event|Event|General Exam|2793,2799|true|false|false|||tested
Anatomy|Body Part, Organ, or Organ Component|General Exam|2804,2810|false|false|false|C0034121|Pupil|Pupils
Event|Event|General Exam|2819,2824|false|false|false|||round
Event|Event|General Exam|2829,2837|false|false|false|||reactive
Procedure|Therapeutic or Preventive Procedure|General Exam|2829,2837|false|false|false|C4722408|Reactive Therapy|reactive
Finding|Finding|General Exam|2829,2846|false|false|false|C4068744|Reactive to light|reactive to light
Drug|Amino Acid, Peptide, or Protein|General Exam|2841,2846|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|General Exam|2841,2846|false|false|false|C1570446|TNFSF14 protein, human|light
Event|Event|General Exam|2841,2846|false|false|false|||light
Finding|Finding|General Exam|2841,2846|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|General Exam|2841,2846|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|General Exam|2841,2846|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|General Exam|2841,2846|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|General Exam|2841,2846|false|false|false|C0031765|Phototherapy|light
Finding|Functional Concept|General Exam|2867,2873|false|false|false|C0234621|Visual|Visual
Event|Event|General Exam|2874,2880|false|false|false|||fields
Event|Event|General Exam|2885,2889|false|false|false|||full
Event|Event|General Exam|2893,2906|false|false|false|||confrontation
Finding|Finding|General Exam|2893,2906|false|false|false|C0518608|Social confrontation skill|confrontation
Procedure|Diagnostic Procedure|General Exam|2893,2906|false|false|false|C0700282;C1444674|Confrontation;Confrontation visual field test|confrontation
Procedure|Therapeutic or Preventive Procedure|General Exam|2893,2906|false|false|false|C0700282;C1444674|Confrontation;Confrontation visual field test|confrontation
Finding|Functional Concept|General Exam|2921,2932|true|false|false|C0241886|Extraocular|Extraocular
Procedure|Diagnostic Procedure|General Exam|2921,2942|true|false|false|C2228439|examination of extraocular movements|Extraocular movements
Event|Event|General Exam|2933,2942|true|false|false|||movements
Finding|Organism Function|General Exam|2933,2942|true|false|false|C0026649|Movement|movements
Event|Event|General Exam|2943,2949|true|false|false|||intact
Finding|Finding|General Exam|2943,2949|true|false|false|C1554187|Gender Status - Intact|intact
Disorder|Disease or Syndrome|General Exam|2970,2979|true|false|false|C0028738|Nystagmus|nystagmus
Event|Event|General Exam|2970,2979|true|false|false|||nystagmus
Anatomy|Body Part, Organ, or Organ Component|General Exam|2984,2987|false|false|false|C2338708;C3496273;C3496274|Lamina VII of gray matter of spinal cord;layer VII (Cajal);lobule VII|VII
Finding|Intellectual Product|General Exam|2984,2987|false|false|false|C0445385|Roman numeral VII|VII
Anatomy|Body Location or Region|General Exam|2989,2995|false|false|false|C0015450|Face|Facial
Event|Event|General Exam|2996,3004|false|false|false|||strength
Finding|Idea or Concept|General Exam|2996,3004|false|false|false|C0808080|Strength (attribute)|strength
Event|Event|General Exam|3009,3018|false|false|false|||sensation
Finding|Finding|General Exam|3009,3018|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|General Exam|3009,3018|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|General Exam|3009,3018|false|false|false|C2229507|sensory exam|sensation
Event|Event|General Exam|3019,3025|false|false|false|||intact
Finding|Finding|General Exam|3019,3025|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|General Exam|3030,3039|false|false|false|||symmetric
Finding|Conceptual Entity|General Exam|3030,3039|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|General Exam|3030,3039|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Anatomy|Body Part, Organ, or Organ Component|General Exam|3041,3045|false|false|false|C0228488;C2327388|Cerebellar pyramis;Lamina VIII of gray matter of spinal cord|VIII
Finding|Gene or Genome|General Exam|3041,3045|false|false|false|C0445599;C1413661|COX8A gene;Roman numeral VIII|VIII
Finding|Intellectual Product|General Exam|3041,3045|false|false|false|C0445599;C1413661|COX8A gene;Roman numeral VIII|VIII
Event|Event|General Exam|3047,3054|false|false|false|||Hearing
Finding|Finding|General Exam|3047,3054|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|Hearing
Finding|Physiologic Function|General Exam|3047,3054|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|Hearing
Event|Event|General Exam|3055,3061|false|false|false|||intact
Finding|Finding|General Exam|3055,3061|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|General Exam|3065,3070|false|false|false|||voice
Finding|Idea or Concept|General Exam|3065,3070|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Intellectual Product|General Exam|3065,3070|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Organism Function|General Exam|3065,3070|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Anatomy|Body Part, Organ, or Organ Component|General Exam|3079,3086|false|false|false|C0700374|Palate|Palatal
Event|Event|General Exam|3087,3096|false|false|false|||elevation
Procedure|Therapeutic or Preventive Procedure|General Exam|3087,3096|false|false|false|C0439775|Elevation procedure|elevation
Event|Event|General Exam|3097,3108|false|false|false|||symmetrical
Finding|Finding|General Exam|3097,3108|false|false|false|C0332516|Symmetrical|symmetrical
Anatomy|Body Part, Organ, or Organ Component|General Exam|3114,3133|false|false|false|C0224153|Structure of sternocleidomastoid muscle|Sternocleidomastoid
Anatomy|Body Part, Organ, or Organ Component|General Exam|3138,3147|false|false|false|C0224361|Structure of trapezius muscle|trapezius
Event|Event|General Exam|3148,3154|false|false|false|||normal
Anatomy|Body Part, Organ, or Organ Component|General Exam|3173,3179|true|false|false|C0040408|Tongue|Tongue
Disorder|Neoplastic Process|General Exam|3173,3179|true|false|false|C0153933|Benign neoplasm of tongue|Tongue
Procedure|Health Care Activity|General Exam|3173,3179|true|false|false|C0872394|Procedure on tongue|Tongue
Finding|Finding|General Exam|3173,3187|true|false|false|C3693372|tongue midline|Tongue midline
Anatomy|Cell Component|General Exam|3180,3187|true|false|false|C1660780|midline cell component|midline
Event|Event|General Exam|3196,3210|true|false|false|||fasciculations
Finding|Sign or Symptom|General Exam|3196,3210|true|false|false|C0015644|Muscular fasciculation|fasciculations
Event|Event|General Exam|3213,3218|false|false|false|||Motor
Finding|Functional Concept|General Exam|3213,3218|false|false|false|C1513492|motor movement|Motor
Drug|Biomedical or Dental Material|General Exam|3227,3231|false|false|false|C0012173;C1337615|Bulk (conceptual);Dietary Fiber|bulk
Drug|Food|General Exam|3227,3231|false|false|false|C0012173;C1337615|Bulk (conceptual);Dietary Fiber|bulk
Event|Event|General Exam|3227,3231|false|false|false|||bulk
Event|Event|General Exam|3236,3240|false|false|false|||tone
Finding|Finding|General Exam|3257,3265|true|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Finding|Idea or Concept|General Exam|3257,3265|true|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Disorder|Disease or Syndrome|General Exam|3257,3275|true|false|false|C0013384|Dyskinetic syndrome|abnormal movements
Finding|Finding|General Exam|3257,3275|true|false|false|C0558189|Abnormal movement|abnormal movements
Event|Event|General Exam|3266,3275|true|false|false|||movements
Finding|Organism Function|General Exam|3266,3275|true|false|false|C0026649|Movement|movements
Event|Event|General Exam|3277,3284|true|false|false|||tremors
Finding|Sign or Symptom|General Exam|3277,3284|true|false|false|C0040822|Tremor|tremors
Finding|Idea or Concept|General Exam|3286,3294|false|false|false|C0808080|Strength (attribute)|Strength
Finding|Social Behavior|General Exam|3300,3305|false|false|false|C0032863|Power (Psychology)|power
Finding|Intellectual Product|General Exam|3322,3326|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Finding|Pathologic Function|General Exam|3335,3349|false|false|false|C1504476|Pronator drift|pronator drift
Event|Event|General Exam|3344,3349|false|false|false|||drift
Finding|Finding|General Exam|3351,3355|false|false|false|C0016928|Gait|Gait
Finding|Finding|General Exam|3351,3364|false|false|false|C0231686|Gait, Unsteady|Gait unsteady
Event|Event|General Exam|3356,3364|false|false|false|||unsteady
Procedure|Diagnostic Procedure|General Exam|3366,3379|false|false|false|C1656968|rhomberg test|rhomberg test
Anatomy|Body Location or Region|General Exam|3375,3379|false|false|false|C4318744|Test - temporal region|test
Event|Event|General Exam|3375,3379|false|false|false|||test
Finding|Functional Concept|General Exam|3375,3379|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|General Exam|3375,3379|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|General Exam|3375,3379|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|General Exam|3375,3379|false|false|false|C0022885|Laboratory Procedures|test
Event|Event|General Exam|3385,3397|false|false|false|||unsteadiness
Finding|Finding|General Exam|3385,3397|false|false|false|C0427108|General unsteadiness|unsteadiness
Event|Event|General Exam|3400,3409|false|false|false|||Sensation
Finding|Finding|General Exam|3400,3409|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Finding|Organ or Tissue Function|General Exam|3400,3409|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Procedure|Health Care Activity|General Exam|3400,3409|false|false|false|C2229507|sensory exam|Sensation
Event|Event|General Exam|3411,3417|false|false|false|||Intact
Finding|Finding|General Exam|3411,3417|false|false|false|C1554187|Gender Status - Intact|Intact
Drug|Amino Acid, Peptide, or Protein|General Exam|3421,3426|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|General Exam|3421,3426|false|false|false|C1570446|TNFSF14 protein, human|light
Finding|Finding|General Exam|3421,3426|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|General Exam|3421,3426|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|General Exam|3421,3426|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|General Exam|3421,3426|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|General Exam|3421,3426|false|false|false|C0031765|Phototherapy|light
Finding|Physiologic Function|General Exam|3421,3432|false|false|false|C0423553|Light touch|light touch
Event|Event|General Exam|3427,3432|false|false|false|||touch
Finding|Mental Process|General Exam|3427,3432|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Finding|Organ or Tissue Function|General Exam|3427,3432|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Procedure|Therapeutic or Preventive Procedure|General Exam|3427,3432|false|false|false|C0152054|Therapeutic Touch|touch
Event|Event|General Exam|3434,3447|false|false|false|||propioception
Disorder|Injury or Poisoning|General Exam|3462,3471|false|false|false|C0677519|Exposed to vibration|vibration
Event|Event|General Exam|3462,3471|false|false|false|||vibration
Phenomenon|Natural Phenomenon or Process|General Exam|3462,3471|false|false|false|C0459800||vibration
Procedure|Therapeutic or Preventive Procedure|General Exam|3462,3471|false|false|false|C0455941|Vibration - treatment|vibration
Event|Event|General Exam|3486,3494|false|false|false|||Reflexes
Finding|Finding|General Exam|3486,3494|false|false|false|C0034929;C0596002|Observation of reflex;Reflex action|Reflexes
Finding|Organ or Tissue Function|General Exam|3486,3494|false|false|false|C0034929;C0596002|Observation of reflex;Reflex action|Reflexes
Procedure|Diagnostic Procedure|General Exam|3486,3494|false|false|false|C0436145|Examination of reflexes|Reflexes
Finding|Functional Concept|General Exam|3509,3514|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Finding|Functional Concept|General Exam|3528,3532|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|General Exam|3548,3552|false|false|false|C0040357;C4299090|Lower extremity>Toes;Toes|Toes
Event|Event|General Exam|3553,3562|false|false|false|||downgoing
Event|Event|General Exam|3576,3588|false|false|false|||Coordination
Finding|Functional Concept|General Exam|3576,3588|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Finding|Idea or Concept|General Exam|3576,3588|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Finding|Physiologic Function|General Exam|3576,3588|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Anatomy|Body Part, Organ, or Organ Component|General Exam|3590,3594|false|false|false|C0018870|Heel|heel
Anatomy|Body Location or Region|General Exam|3598,3602|false|false|false|C0230444|Shin|shin
Event|Event|General Exam|3603,3609|false|false|false|||intact
Finding|Finding|General Exam|3603,3609|false|false|false|C1554187|Gender Status - Intact|intact
Anatomy|Body Part, Organ, or Organ Component|General Exam|3611,3617|false|false|false|C0016129;C0851278;C4299059|Fingers;Fingers not including thumb;Upper extremity>Finger|finger
Anatomy|Body Part, Organ, or Organ Component|General Exam|3623,3629|false|false|false|C0016129;C0851278;C4299059|Fingers;Fingers not including thumb;Upper extremity>Finger|finger
Event|Event|General Exam|3630,3636|false|false|false|||slowed
Event|Event|General Exam|3641,3653|false|false|false|||overshooting
Anatomy|Body Part, Organ, or Organ Component|General Exam|3659,3665|false|false|false|C0230370|Structure of right hand|R hand
Anatomy|Body Part, Organ, or Organ Component|General Exam|3661,3665|false|false|false|C0018563;C4285005|Hand;Upper extremity>Hand|hand
Finding|Finding|General Exam|3661,3665|false|false|false|C0741992|Hand problem|hand
Event|Event|General Exam|3667,3677|false|false|false|||Difficulty
Finding|Finding|General Exam|3667,3677|false|false|false|C1299586|Has difficulty doing (qualifier value)|Difficulty
Finding|Finding|General Exam|3667,3682|false|false|false|C0332218|Difficult (qualifier value)|Difficulty with
Event|Event|General Exam|3689,3700|false|false|false|||alternating
Finding|Functional Concept|General Exam|3689,3700|false|false|false|C0332270|Alternating|alternating
Event|Event|General Exam|3701,3710|false|false|false|||movements
Finding|Organism Function|General Exam|3701,3710|false|false|false|C0026649|Movement|movements
Anatomy|Body Part, Organ, or Organ Component|General Exam|3716,3722|false|false|false|C0230370|Structure of right hand|R hand
Anatomy|Body Part, Organ, or Organ Component|General Exam|3718,3722|false|false|false|C0018563;C4285005|Hand;Upper extremity>Hand|hand
Finding|Finding|General Exam|3718,3722|false|false|false|C0741992|Hand problem|hand
Event|Event|General Exam|3728,3737|false|false|false|||DISCHARGE
Finding|Body Substance|General Exam|3728,3737|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|3728,3737|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|3728,3737|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|3728,3737|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|General Exam|3746,3749|false|false|false|||VSS
Event|Event|General Exam|3750,3753|false|false|false|||Gen
Finding|Classification|General Exam|3750,3753|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Finding|Gene or Genome|General Exam|3750,3753|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Disorder|Disease or Syndrome|General Exam|3755,3758|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|3755,3758|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|3755,3758|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|3755,3758|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|3755,3758|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|General Exam|3755,3758|false|false|false|||NAD
Finding|Finding|General Exam|3755,3758|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|General Exam|3760,3765|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|General Exam|3767,3773|false|false|false|C0034121|Pupil|Pupils
Event|Event|General Exam|3781,3785|false|false|false|||EOMs
Finding|Functional Concept|General Exam|3781,3785|false|false|false|C0241886|Extraocular|EOMs
Finding|Finding|General Exam|3786,3792|false|false|false|C1554187|Gender Status - Intact|intact
Anatomy|Body Part, Organ, or Organ Component|General Exam|3797,3802|false|false|false|C0024109|Lung|Lungs
Finding|Idea or Concept|General Exam|3804,3809|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Part, Organ, or Organ Component|General Exam|3814,3821|false|false|false|C0018787|Heart|Cardiac
Finding|Intellectual Product|General Exam|3814,3821|false|false|false|C1314974|Cardiac attachment|Cardiac
Finding|Finding|General Exam|3844,3863|false|false|false|C0232258|Pansystolic murmur|holosystolic murmur
Event|Event|General Exam|3857,3863|false|false|false|||murmur
Finding|Finding|General Exam|3857,3863|false|false|false|C0018808|Heart murmur|murmur
Anatomy|Body Location or Region|General Exam|3865,3868|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|Abd
Disorder|Cell or Molecular Dysfunction|General Exam|3865,3868|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|Abd
Attribute|Clinical Attribute|General Exam|3906,3911|true|false|false|C1717255||edema
Event|Event|General Exam|3906,3911|true|false|false|||edema
Finding|Pathologic Function|General Exam|3906,3911|true|false|false|C0013604|Edema|edema
Disorder|Disease or Syndrome|General Exam|3915,3923|true|false|false|C0041834|Erythema|erythema
Event|Event|General Exam|3915,3923|true|false|false|||erythema
Finding|Finding|General Exam|3925,3929|true|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|General Exam|3925,3929|true|false|false|C0687712|warming process|warm
Finding|Finding|General Exam|3930,3934|true|false|false|C5575035|Well (answer to question)|well
Finding|Mental Process|General Exam|3953,3959|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|General Exam|3953,3966|false|false|false|C0488568;C0488569||Mental status
Finding|Finding|General Exam|3953,3966|false|false|false|C0278060|Mental state|Mental status
Attribute|Clinical Attribute|General Exam|3960,3966|false|false|false|C5889824||status
Event|Event|General Exam|3960,3966|false|false|false|||status
Finding|Idea or Concept|General Exam|3960,3966|false|false|false|C1546481|What subject filter - Status|status
Event|Event|General Exam|3968,3973|false|false|false|||Awake
Finding|Finding|General Exam|3968,3973|false|false|false|C0234422|Awake (finding)|Awake
Event|Event|General Exam|3978,3989|false|false|false|||cooperative
Event|Event|General Exam|3995,3999|false|false|false|||exam
Finding|Functional Concept|General Exam|3995,3999|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|General Exam|3995,3999|false|false|false|C0582103|Medical Examination|exam
Event|Event|General Exam|4008,4014|false|false|false|||affect
Finding|Mental Process|General Exam|4008,4014|false|false|false|C0001721|Affect (mental function)|affect
Procedure|Health Care Activity|General Exam|4008,4014|false|false|false|C2237113|assessment of affect|affect
Event|Event|General Exam|4016,4027|false|false|false|||Orientation
Finding|Mental Process|General Exam|4016,4027|false|false|false|C0029266|Mental Orientation|Orientation
Event|Event|General Exam|4029,4037|false|false|false|||Oriented
Finding|Finding|General Exam|4029,4037|false|false|false|C1961028|Oriented to place|Oriented
Finding|Finding|General Exam|4029,4047|false|false|false|C1961030|Oriented to person|Oriented to person
Attribute|Clinical Attribute|General Exam|4041,4047|false|false|false|C5890614||person
Event|Event|General Exam|4041,4047|false|false|false|||person
Finding|Intellectual Product|General Exam|4041,4047|false|false|false|C1522390|Person Info|person
Event|Activity|General Exam|4049,4054|false|false|false|C1882509|put - instruction imperative|place
Event|Event|General Exam|4049,4054|false|false|false|||place
Finding|Functional Concept|General Exam|4049,4054|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|General Exam|4049,4054|false|false|false|C1533810||place
Attribute|Clinical Attribute|General Exam|4066,4074|false|false|false|C2706915||Language
Event|Event|General Exam|4066,4074|false|false|false|||Language
Finding|Intellectual Product|General Exam|4066,4074|false|false|false|C0033348|Programming Languages|Language
Event|Event|General Exam|4076,4082|false|false|false|||Speech
Finding|Organism Function|General Exam|4076,4082|false|false|false|C0037817|Speech|Speech
Procedure|Diagnostic Procedure|General Exam|4076,4082|false|false|false|C0846595|Speech assessment|Speech
Event|Event|General Exam|4086,4092|false|false|false|||fluent
Finding|Idea or Concept|General Exam|4094,4098|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Event|Event|General Exam|4099,4112|false|false|false|||comprehension
Finding|Mental Process|General Exam|4099,4112|false|false|false|C0162340|Comprehension|comprehension
Anatomy|Body Part, Organ, or Organ Component|General Exam|4115,4122|false|false|false|C0037303|Bone structure of cranium|Cranial
Anatomy|Body Part, Organ, or Organ Component|General Exam|4115,4129|false|false|false|C0010268|Cranial Nerves|Cranial Nerves
Disorder|Neoplastic Process|General Exam|4115,4129|false|false|false|C0004992;C0496937|Benign neoplasm of cranial nerves;Neoplasm of uncertain or unknown behavior of cranial nerves|Cranial Nerves
Anatomy|Body Part, Organ, or Organ Component|General Exam|4123,4129|false|false|false|C0027740|Nerve|Nerves
Finding|Functional Concept|General Exam|4138,4144|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|tested
Finding|Intellectual Product|General Exam|4138,4144|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|tested
Event|Event|General Exam|4149,4155|false|false|false|||intact
Finding|Finding|General Exam|4149,4155|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|General Exam|4161,4166|false|false|false|||Motor
Finding|Functional Concept|General Exam|4161,4166|false|false|false|C1513492|motor movement|Motor
Event|Event|General Exam|4172,4180|false|false|false|||strength
Finding|Idea or Concept|General Exam|4172,4180|false|false|false|C0808080|Strength (attribute)|strength
Finding|Pathologic Function|General Exam|4203,4217|true|false|false|C1504476|Pronator drift|pronator drift
Event|Event|General Exam|4212,4217|true|false|false|||drift
Finding|Finding|General Exam|4219,4223|true|false|false|C0016928|Gait|Gait
Event|Event|General Exam|4233,4240|true|false|false|||walking
Finding|Daily or Recreational Activity|General Exam|4233,4240|true|false|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Finding|Finding|General Exam|4233,4240|true|false|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Finding|Sign or Symptom|General Exam|4233,4240|true|false|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Event|Event|General Exam|4249,4259|true|false|false|||assistance
Finding|Social Behavior|General Exam|4249,4259|true|false|false|C0018896|Helping Behavior|assistance
Event|Event|General Exam|4262,4271|false|false|false|||Sensation
Finding|Finding|General Exam|4262,4271|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Finding|Organ or Tissue Function|General Exam|4262,4271|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Procedure|Health Care Activity|General Exam|4262,4271|false|false|false|C2229507|sensory exam|Sensation
Event|Event|General Exam|4281,4287|false|false|false|||intact
Finding|Finding|General Exam|4281,4287|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|General Exam|4294,4302|false|false|false|||Reflexes
Finding|Finding|General Exam|4294,4302|false|false|false|C0034929;C0596002|Observation of reflex;Reflex action|Reflexes
Finding|Organ or Tissue Function|General Exam|4294,4302|false|false|false|C0034929;C0596002|Observation of reflex;Reflex action|Reflexes
Procedure|Diagnostic Procedure|General Exam|4294,4302|false|false|false|C0436145|Examination of reflexes|Reflexes
Finding|Functional Concept|General Exam|4317,4322|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Finding|Functional Concept|General Exam|4336,4340|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|General Exam|4356,4360|false|false|false|C0040357;C4299090|Lower extremity>Toes;Toes|Toes
Event|Event|General Exam|4361,4370|false|false|false|||downgoing
Disorder|Disease or Syndrome|General Exam|4416,4421|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4416,4421|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4416,4421|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|4422,4425|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|4431,4434|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|4431,4434|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|4431,4434|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|4441,4444|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|4441,4444|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|4441,4444|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|4441,4444|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|4451,4454|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|4451,4454|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|4461,4464|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|4461,4464|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|4461,4464|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|4461,4464|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|4461,4464|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|4468,4471|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|4468,4471|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|4468,4471|false|false|false|||MCH
Finding|Gene or Genome|General Exam|4468,4471|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|4468,4471|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|4468,4471|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|4477,4481|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|4477,4481|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|4496,4499|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|4516,4521|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4516,4521|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4516,4521|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|General Exam|4538,4543|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4538,4543|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4538,4543|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|4538,4551|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|4538,4551|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|4538,4551|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|4544,4551|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|4544,4551|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|4544,4551|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|4544,4551|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|4544,4551|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|4544,4551|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|4598,4602|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|4598,4602|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|4598,4602|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|4627,4632|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4627,4632|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4627,4632|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|4627,4640|false|false|false|C0853248|Blood albumin|BLOOD Albumin
Drug|Amino Acid, Peptide, or Protein|General Exam|4633,4640|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Biologically Active Substance|General Exam|4633,4640|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Pharmacologic Substance|General Exam|4633,4640|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Event|Event|General Exam|4633,4640|false|false|false|||Albumin
Finding|Gene or Genome|General Exam|4633,4640|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Finding|Physiologic Function|General Exam|4633,4640|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Procedure|Laboratory Procedure|General Exam|4633,4640|false|false|false|C0201838|Albumin measurement|Albumin
Disorder|Disease or Syndrome|General Exam|4658,4663|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4658,4663|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4658,4663|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|4665,4670|false|false|false|C0019018|Glycosylated hemoglobin A|HbA1c
Drug|Biologically Active Substance|General Exam|4665,4670|false|false|false|C0019018|Glycosylated hemoglobin A|HbA1c
Event|Event|General Exam|4665,4670|false|false|false|||HbA1c
Procedure|Laboratory Procedure|General Exam|4665,4670|false|false|false|C0202054|Glucohemoglobin measurement|HbA1c
Finding|Gene or Genome|General Exam|4676,4679|false|false|false|C1416571|KCNH1 gene|eAG
Disorder|Disease or Syndrome|General Exam|4697,4702|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4697,4702|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4697,4702|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Attribute|Clinical Attribute|General Exam|4717,4724|false|false|false|C0881943||CT Head
Procedure|Diagnostic Procedure|General Exam|4717,4724|false|false|false|C0202691|CAT scan of head|CT Head
Anatomy|Body Location or Region|General Exam|4720,4724|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|Head
Anatomy|Body Part, Organ, or Organ Component|General Exam|4720,4724|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|Head
Disorder|Disease or Syndrome|General Exam|4720,4724|false|false|false|C0362076|Problems with head|Head
Event|Event|General Exam|4720,4724|false|false|false|||Head
Procedure|Therapeutic or Preventive Procedure|General Exam|4720,4724|false|false|false|C0876917|Procedure on head|Head
Event|Event|Impression|4759,4765|false|false|false|||lesion
Finding|Finding|Impression|4759,4765|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|Impression|4759,4765|false|false|false|C0221198;C1546698|Lesion|lesion
Event|Event|Impression|4778,4782|false|false|false|||foci
Finding|Finding|Impression|4778,4782|false|false|false|C4321394|Foci|foci
Event|Event|Impression|4786,4800|false|false|false|||calcifications
Finding|Finding|Impression|4786,4800|false|false|false|C0006660;C2242558|Pathologic calcification, calcified structure;Physiologic calcification|calcifications
Finding|Organ or Tissue Function|Impression|4786,4800|false|false|false|C0006660;C2242558|Pathologic calcification, calcified structure;Physiologic calcification|calcifications
Event|Event|Impression|4802,4811|false|false|false|||measuring
Finding|Finding|Impression|4830,4836|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Impression|4830,4836|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|Impression|4837,4845|false|false|false|||reflects
Event|Event|Impression|4861,4865|false|false|false|||mass
Finding|Finding|Impression|4861,4865|false|true|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|Impression|4861,4865|false|true|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Impression|4861,4865|false|true|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Disorder|Neoplastic Process|Impression|4877,4887|false|false|false|C0025286;C0281784|Benign Meningioma;Meningioma|meningioma
Event|Event|Impression|4877,4887|false|false|false|||meningioma
Event|Event|Impression|4905,4913|false|false|false|||hematoma
Finding|Pathologic Function|Impression|4905,4913|false|false|false|C0018944|Hematoma|hematoma
Event|Event|Impression|4930,4938|false|false|false|||subacute
Event|Event|Impression|4942,4949|false|false|false|||chronic
Finding|Intellectual Product|Impression|4942,4949|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Impression|4942,4949|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Event|Event|Impression|4955,4965|false|false|false|||considered
Event|Event|Impression|4971,4977|false|false|false|||likely
Finding|Finding|Impression|4971,4977|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Impression|4971,4977|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|Impression|4983,4987|false|false|false|||Loss
Finding|Finding|Impression|4983,4987|false|false|false|C5890125|Loss (adaptation)|Loss
Attribute|Clinical Attribute|Impression|5002,5017|false|false|false|C1511938|Cellular Differentiation Qualifier|differentiation
Event|Event|Impression|5002,5017|false|false|false|||differentiation
Finding|Cell Function|Impression|5002,5017|false|false|false|C0007589;C2945687|Cell Differentiation process;Differentiation|differentiation
Finding|Functional Concept|Impression|5002,5017|false|false|false|C0007589;C2945687|Cell Differentiation process;Differentiation|differentiation
Finding|Finding|Impression|5025,5029|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|Impression|5025,5029|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|Impression|5025,5029|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Functional Concept|Impression|5030,5034|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Impression|5051,5055|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|Impression|5051,5055|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Event|Event|Impression|5063,5070|false|false|false|||reflect
Finding|Intellectual Product|Impression|5074,5079|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Pathologic Function|Impression|5074,5087|false|false|false|C0333548|Acute infarct|acute infarct
Event|Event|Impression|5080,5087|false|false|false|||infarct
Finding|Pathologic Function|Impression|5080,5087|false|false|false|C0021308|Infarction|infarct
Event|Event|Impression|5091,5094|false|false|false|||MRI
Finding|Gene or Genome|Impression|5091,5094|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|Impression|5091,5094|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|Impression|5091,5094|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Diagnostic Procedure|Impression|5091,5099|false|false|false|C0412674|MRI of head|MRI Head
Anatomy|Body Location or Region|Impression|5095,5099|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|Head
Anatomy|Body Part, Organ, or Organ Component|Impression|5095,5099|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|Head
Disorder|Disease or Syndrome|Impression|5095,5099|false|false|false|C0362076|Problems with head|Head
Procedure|Therapeutic or Preventive Procedure|Impression|5095,5099|false|false|false|C0876917|Procedure on head|Head
Event|Event|Impression|5105,5110|false|false|false|||Acute
Finding|Intellectual Product|Impression|5105,5110|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Event|Event|Impression|5133,5144|false|false|false|||infarctions
Finding|Pathologic Function|Impression|5133,5144|false|false|false|C0021308|Infarction|infarctions
Event|Event|Impression|5162,5167|false|false|false|||focus
Finding|Functional Concept|Impression|5162,5167|false|false|false|C1285542|Has focus|focus
Finding|Functional Concept|Impression|5176,5180|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Attribute|Clinical Attribute|Impression|5201,5211|false|false|false|C0550215||Appearance
Event|Event|Impression|5201,5211|false|false|false|||Appearance
Procedure|Health Care Activity|Impression|5201,5211|false|false|false|C2051406|patient appearance regarding mental status exam|Appearance
Event|Event|Impression|5231,5237|false|false|false|||lesion
Finding|Finding|Impression|5231,5237|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|Impression|5231,5237|false|false|false|C0221198;C1546698|Lesion|lesion
Event|Event|Impression|5241,5249|false|false|false|||somewhat
Finding|Finding|Impression|5241,5249|false|false|false|C2984079|Somewhat|somewhat
Event|Event|Impression|5277,5286|false|false|false|||recommend
Event|Event|Impression|5287,5296|false|false|false|||attention
Finding|Intellectual Product|Impression|5287,5296|false|false|false|C0004268;C4281780|Attention;Attention - G-code|attention
Finding|Mental Process|Impression|5287,5296|false|false|false|C0004268;C4281780|Attention;Attention - G-code|attention
Event|Event|Impression|5300,5308|true|false|false|||followup
Procedure|Health Care Activity|Impression|5300,5308|true|false|false|C1522577|follow-up|followup
Event|Event|Impression|5310,5317|true|false|false|||imaging
Finding|Finding|Impression|5310,5317|true|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|Impression|5310,5317|true|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Event|Event|Impression|5330,5340|true|false|false|||evaluation
Finding|Idea or Concept|Impression|5330,5340|true|true|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|Impression|5330,5340|true|true|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Event|Event|Impression|5344,5351|false|false|false|||exclude
Event|Event|Impression|5356,5364|true|false|false|||presence
Procedure|Therapeutic or Preventive Procedure|Impression|5356,5364|true|false|false|C0392148|Providing presence (regime/therapy)|presence
Finding|Finding|Impression|5356,5367|true|false|false|C0150312|Present|presence of
Event|Event|Impression|5383,5387|true|false|false|||mass
Finding|Finding|Impression|5383,5387|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|Impression|5383,5387|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Impression|5383,5387|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Disorder|Neoplastic Process|Impression|5393,5404|true|false|false|C0025286|Meningioma|meningiomas
Event|Event|Impression|5393,5404|true|false|false|||meningiomas
Finding|Functional Concept|Impression|5412,5416|true|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|Impression|5417,5431|true|false|false|C0016733;C0162783;C0549224|Frontal region;Prefrontal Cortex;frontal lobe|frontal region
Anatomy|Body Part, Organ, or Organ Component|Impression|5417,5431|true|false|false|C0016733;C0162783;C0549224|Frontal region;Prefrontal Cortex;frontal lobe|frontal region
Drug|Amino Acid Sequence|Impression|5425,5431|true|false|false|C1514562|Protein Domain|region
Finding|Idea or Concept|Impression|5441,5452|true|false|false|C0750502|Significant|significant
Event|Event|Impression|5453,5457|true|false|false|||mass
Finding|Finding|Impression|5453,5457|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|Impression|5453,5457|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Impression|5453,5457|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Finding|Impression|5453,5464|true|false|false|C4086564|Mass Effect|mass effect
Event|Event|Impression|5458,5464|true|false|false|||effect
Event|Event|Impression|5467,5471|false|false|false|||ECHO
Procedure|Health Care Activity|Impression|5467,5471|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Procedure|Therapeutic or Preventive Procedure|Impression|5467,5471|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Finding|Conceptual Entity|Impression|5484,5493|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|Impression|5484,5493|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Functional Concept|Impression|5494,5498|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Attribute|Clinical Attribute|Impression|5494,5522|false|false|false|C3484363||left ventricular hypertrophy
Disorder|Disease or Syndrome|Impression|5494,5522|false|false|false|C0149721|Left Ventricular Hypertrophy|left ventricular hypertrophy
Anatomy|Body Part, Organ, or Organ Component|Impression|5499,5510|false|false|false|C0018827|Heart Ventricle|ventricular
Disorder|Disease or Syndrome|Impression|5499,5522|false|false|false|C0340279|Ventricular hypertrophy|ventricular hypertrophy
Event|Event|Impression|5511,5522|false|false|false|||hypertrophy
Finding|Pathologic Function|Impression|5511,5522|false|false|false|C0020564|Hypertrophy|hypertrophy
Anatomy|Body Space or Junction|Impression|5535,5541|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|Impression|5535,5541|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|Impression|5535,5541|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Finding|Organ or Tissue Function|Impression|5568,5576|false|false|false|C0039155|Systole|systolic
Event|Event|Impression|5577,5585|false|false|false|||function
Finding|Finding|Impression|5577,5585|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|Impression|5577,5585|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|Impression|5577,5585|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|Impression|5577,5585|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|Impression|5587,5591|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Anatomy|Body Part, Organ, or Organ Component|Impression|5592,5598|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|Impression|5592,5604|false|false|false|C0003501;C4533215|Aortic valve structure;Chest>Aortic valve|aortic valve
Anatomy|Body Part, Organ, or Organ Component|Impression|5599,5604|false|false|false|C1186983|Anatomical valve|valve
Event|Event|Impression|5606,5614|false|false|false|||stenosis
Finding|Pathologic Function|Impression|5606,5614|false|false|false|C1261287|Stenosis|stenosis
Finding|Intellectual Product|Impression|5616,5620|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Anatomy|Body Part, Organ, or Organ Component|Impression|5621,5627|false|false|false|C0003483|Aorta|aortic
Disorder|Disease or Syndrome|Impression|5621,5641|false|false|false|C0003504|Aortic Valve Insufficiency|aortic regurgitation
Event|Event|Impression|5628,5641|false|false|false|||regurgitation
Finding|Finding|Impression|5628,5641|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|Impression|5628,5641|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|Impression|5628,5641|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Finding|Functional Concept|Impression|5643,5648|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Part, Organ, or Organ Component|Impression|5643,5670|false|false|false|C4288280|Right Ventricular Free Wall|Right ventricular free wall
Anatomy|Body Part, Organ, or Organ Component|Impression|5649,5660|false|false|false|C0018827|Heart Ventricle|ventricular
Event|Event|Impression|5661,5665|false|false|false|||free
Finding|Functional Concept|Impression|5661,5665|false|false|false|C0332296|Free of (attribute)|free
Event|Event|Impression|5672,5683|false|false|false|||hypertrophy
Finding|Pathologic Function|Impression|5672,5683|false|false|false|C0020564|Hypertrophy|hypertrophy
Anatomy|Body Part, Organ, or Organ Component|Impression|5685,5694|false|false|false|C0024109|Lung|Pulmonary
Attribute|Clinical Attribute|Impression|5685,5694|false|false|false|C2707265||Pulmonary
Finding|Finding|Impression|5685,5694|false|false|false|C4522268|Pulmonary (intended site)|Pulmonary
Anatomy|Body Part, Organ, or Organ Component|Impression|5685,5701|false|false|false|C0034052|Pulmonary artery structure|Pulmonary artery
Anatomy|Body Part, Organ, or Organ Component|Impression|5695,5701|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|Impression|5695,5701|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Finding|Organ or Tissue Function|Impression|5702,5710|false|false|false|C0039155|Systole|systolic
Disorder|Disease or Syndrome|Impression|5702,5723|false|false|false|C0221155|Systolic Hypertension|systolic hypertension
Disorder|Disease or Syndrome|Impression|5711,5723|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|Impression|5711,5723|false|false|false|||hypertension
Finding|Finding|Impression|5725,5732|false|false|false|C0700124|Dilated|Dilated
Finding|Functional Concept|Impression|5734,5743|false|false|false|C1547175;C1962987|Ascend (action);Sequencing - Ascending|ascending
Anatomy|Body Part, Organ, or Organ Component|Impression|5734,5749|false|false|false|C0003956|Ascending aorta structure|ascending aorta
Anatomy|Body Part, Organ, or Organ Component|Impression|5744,5749|false|false|false|C0003483;C4037978|Aorta;Chest+Abdomen>Aorta|aorta
Procedure|Health Care Activity|Impression|5744,5749|false|false|false|C0869784|Procedure on aorta|aorta
Finding|Intellectual Product|Impression|5752,5760|false|false|false|C1315013|Clinical NEC (not elsewhere classified in LNC)|CLINICAL
Finding|Body Substance|Impression|5780,5787|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Impression|5780,5787|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Impression|5780,5787|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|Impression|5780,5791|false|false|false|C0332310|Has patient|patient has
Finding|Intellectual Product|Impression|5792,5796|false|false|false|C1547225|Mild Severity of Illness Code|mild
Anatomy|Body Part, Organ, or Organ Component|Impression|5797,5803|false|false|false|C0003483|Aorta|aortic
Finding|Pathologic Function|Impression|5797,5812|false|false|false|C0003507|Aortic Valve Stenosis|aortic stenosis
Event|Event|Impression|5804,5812|false|false|false|||stenosis
Finding|Pathologic Function|Impression|5804,5812|false|false|false|C1261287|Stenosis|stenosis
Anatomy|Body Part, Organ, or Organ Component|Impression|5827,5830|false|false|false|C0152325;C2954192|Gray matter of anterior cingulate gyrus;Structure of forceps minor|ACC
Anatomy|Tissue|Impression|5827,5830|false|false|false|C0152325;C2954192|Gray matter of anterior cingulate gyrus;Structure of forceps minor|ACC
Disorder|Congenital Abnormality|Impression|5827,5830|false|false|false|C0175754;C0206686;C0282160|Adrenocortical carcinoma;Agenesis of corpus callosum;Aplasia Cutis Congenita|ACC
Disorder|Neoplastic Process|Impression|5827,5830|false|false|false|C0175754;C0206686;C0282160|Adrenocortical carcinoma;Agenesis of corpus callosum;Aplasia Cutis Congenita|ACC
Drug|Amino Acid, Peptide, or Protein|Impression|5827,5830|false|false|false|C3541857;C4724142|Acetyl-CoA Carboxylase 1;Amorphous Calcium Carbonate|ACC
Drug|Enzyme|Impression|5827,5830|false|false|false|C3541857;C4724142|Acetyl-CoA Carboxylase 1;Amorphous Calcium Carbonate|ACC
Drug|Pharmacologic Substance|Impression|5827,5830|false|false|false|C3541857;C4724142|Acetyl-CoA Carboxylase 1;Amorphous Calcium Carbonate|ACC
Event|Event|Impression|5827,5830|false|false|false|||ACC
Finding|Gene or Genome|Impression|5827,5830|false|false|false|C1412104;C3541413|ACACA gene;ACACA wt Allele|ACC
Disorder|Disease or Syndrome|Impression|5831,5834|false|false|false|C0002880;C0272325|Autoimmune hemolytic anemia;Factor 8 deficiency, acquired|AHA
Drug|Organic Chemical|Impression|5831,5834|false|false|false|C0050451|acetohydroxamic acid|AHA
Drug|Pharmacologic Substance|Impression|5831,5834|false|false|false|C0050451|acetohydroxamic acid|AHA
Event|Event|Impression|5831,5834|false|false|false|||AHA
Disorder|Disease or Syndrome|Impression|5836,5858|false|false|false|C0018824|Heart valve disease|Valvular Heart Disease
Anatomy|Body Part, Organ, or Organ Component|Impression|5845,5850|false|false|false|C0018787;C4037974|Chest>Heart;Heart|Heart
Disorder|Neoplastic Process|Impression|5845,5850|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|Heart
Finding|Sign or Symptom|Impression|5845,5850|false|false|false|C0795691|HEART PROBLEM|Heart
Disorder|Disease or Syndrome|Impression|5845,5858|false|false|false|C0018799|Heart Diseases|Heart Disease
Disorder|Disease or Syndrome|Impression|5851,5858|false|false|false|C0012634|Disease|Disease
Event|Event|Impression|5859,5869|false|false|false|||Guidelines
Finding|Intellectual Product|Impression|5859,5869|false|false|false|C0162791;C0220845;C0282423|Guideline (Publication Type);Guidelines;guiding characteristics|Guidelines
Event|Event|Impression|5873,5879|false|false|false|||follow
Finding|Functional Concept|Impression|5873,5879|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|Impression|5873,5879|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|Impression|5873,5882|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|Impression|5873,5882|false|false|false|C1522577|follow-up|follow-up
Event|Event|Impression|5883,5897|false|false|false|||echocardiogram
Procedure|Diagnostic Procedure|Impression|5883,5897|false|false|false|C0013516|Echocardiography|echocardiogram
Event|Event|Impression|5902,5911|false|false|false|||suggested
Disorder|Disease or Syndrome|Impression|5944,5956|false|false|false|C0014118|Endocarditis|endocarditis
Procedure|Therapeutic or Preventive Procedure|Impression|5944,5968|false|false|false|C1396567|Endocarditis prophylaxis|endocarditis prophylaxis
Procedure|Therapeutic or Preventive Procedure|Impression|5957,5968|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Event|Event|Impression|5969,5984|false|false|false|||recommendations
Finding|Idea or Concept|Impression|5969,5984|false|false|false|C0034866|Recommendation|recommendations
Procedure|Health Care Activity|Impression|5991,5995|true|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Procedure|Therapeutic or Preventive Procedure|Impression|5991,5995|true|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Attribute|Clinical Attribute|Impression|5996,6004|true|false|false|C2926606||findings
Event|Event|Impression|5996,6004|true|false|false|||findings
Finding|Functional Concept|Impression|5996,6004|true|false|false|C2607943|findings aspects|findings
Event|Event|Impression|6014,6025|true|false|false|||prophylaxis
Procedure|Therapeutic or Preventive Procedure|Impression|6014,6025|true|false|false|C0199176|Prophylactic treatment|prophylaxis
Event|Event|Impression|6033,6044|true|false|false|||recommended
Finding|Intellectual Product|Impression|6046,6054|false|false|false|C1315013|Clinical NEC (not elsewhere classified in LNC)|Clinical
Event|Event|Impression|6056,6065|false|false|false|||decisions
Finding|Mental Process|Impression|6056,6065|false|false|false|C0679006|Decision|decisions
Event|Event|Impression|6080,6084|false|false|false|||need
Finding|Functional Concept|Impression|6080,6084|false|false|false|C0686904|Patient need for (contextual qualifier)|need
Finding|Functional Concept|Impression|6080,6088|false|false|false|C0686904|Patient need for (contextual qualifier)|need for
Event|Event|Impression|6089,6100|false|false|false|||prophylaxis
Procedure|Therapeutic or Preventive Procedure|Impression|6089,6100|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Event|Event|Impression|6111,6116|false|false|false|||based
Event|Event|Impression|6121,6129|false|false|false|||clinical
Finding|Intellectual Product|Impression|6121,6129|false|false|false|C1315013|Clinical NEC (not elsewhere classified in LNC)|clinical
Event|Event|Impression|6152,6156|false|false|false|||data
Finding|Idea or Concept|Impression|6152,6156|false|false|false|C1511726|Data|data
Drug|Amino Acid, Peptide, or Protein|Impression|6160,6163|false|false|false|C1609165|tocilizumab|MRA
Drug|Immunologic Factor|Impression|6160,6163|false|false|false|C1609165|tocilizumab|MRA
Drug|Pharmacologic Substance|Impression|6160,6163|false|false|false|C1609165|tocilizumab|MRA
Event|Event|Impression|6160,6163|false|false|false|||MRA
Lab|Laboratory or Test Result|Impression|6160,6163|false|false|false|C3891069|MRI-Based Angiogram|MRA
Procedure|Diagnostic Procedure|Impression|6160,6163|false|false|false|C0243032|Magnetic Resonance Angiography|MRA
Procedure|Diagnostic Procedure|Impression|6160,6168|false|false|false|C1636167|Magnetic resonance angiography of vascular structure of head|MRA Head
Anatomy|Body Location or Region|Impression|6164,6168|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|Head
Anatomy|Body Part, Organ, or Organ Component|Impression|6164,6168|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|Head
Disorder|Disease or Syndrome|Impression|6164,6168|false|false|false|C0362076|Problems with head|Head
Event|Event|Impression|6164,6168|false|false|false|||Head
Procedure|Therapeutic or Preventive Procedure|Impression|6164,6168|false|false|false|C0876917|Procedure on head|Head
Anatomy|Body Location or Region|Impression|6169,6173|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|Impression|6169,6173|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|Impression|6169,6173|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Finding|Intellectual Product|Impression|6179,6183|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Finding|Functional Concept|Impression|6184,6199|false|false|false|C0333482|atherosclerotic|atherosclerotic
Disorder|Disease or Syndrome|Impression|6200,6207|false|false|false|C0012634|Disease|disease
Event|Event|Impression|6200,6207|false|false|false|||disease
Anatomy|Body Part, Organ, or Organ Component|Impression|6215,6229|false|false|false|C0004811|Structure of basilar artery|basilar artery
Anatomy|Body Part, Organ, or Organ Component|Impression|6223,6229|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|Impression|6223,6229|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Event|Event|Impression|6244,6252|true|false|false|||evidence
Finding|Idea or Concept|Impression|6244,6252|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Impression|6244,6255|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Finding|Intellectual Product|Impression|6256,6261|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Part, Organ, or Organ Component|Impression|6262,6270|true|false|false|C0005847|Blood Vessel|vascular
Finding|Finding|Impression|6262,6284|true|false|false|C0241657|Abnormality of the vasculature|vascular abnormalities
Disorder|Congenital Abnormality|Impression|6271,6284|true|false|false|C0000768|Congenital Abnormality|abnormalities
Event|Event|Impression|6271,6284|true|false|false|||abnormalities
Finding|Functional Concept|Impression|6271,6284|true|false|false|C0000769|teratologic|abnormalities
Event|Event|Impression|6285,6294|true|false|false|||involving
Anatomy|Body Location or Region|Impression|6300,6312|false|false|false|C0524466|Intracranial|intracranial
Finding|Functional Concept|Impression|6300,6312|false|false|false|C1522213|Intracranial Route of Administration|intracranial
Anatomy|Body Part, Organ, or Organ Component|Impression|6313,6321|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Anatomy|Body System|Impression|6313,6321|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Procedure|Health Care Activity|Impression|6313,6321|false|false|false|C0397581|Procedure on artery|arteries
Event|Event|Hospital Course|6364,6372|false|false|false|||admitted
Event|Occupational Activity|Hospital Course|6394,6401|false|false|false|C0557854|Services|service
Finding|Idea or Concept|Hospital Course|6394,6401|false|false|false|C3245478|ActInformationPrivacyReason - service|service
Event|Event|Hospital Course|6419,6428|false|false|false|||emergency
Finding|Finding|Hospital Course|6419,6428|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Idea or Concept|Hospital Course|6419,6428|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Intellectual Product|Hospital Course|6419,6428|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Pathologic Function|Hospital Course|6419,6428|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Phenomenon|Phenomenon or Process|Hospital Course|6419,6428|false|false|false|C0013956|Emergency Situation|emergency
Procedure|Health Care Activity|Hospital Course|6419,6428|false|false|false|C1553500|emergency encounter|emergency
Finding|Idea or Concept|Hospital Course|6419,6433|false|false|false|C1546435|Encounter Referral Source - emergency room|emergency room
Event|Event|Hospital Course|6449,6455|false|false|false|||series
Disorder|Injury or Poisoning|Hospital Course|6459,6464|false|false|false|C0000921|Accidental Falls|falls
Event|Event|Hospital Course|6459,6464|false|false|false|||falls
Finding|Finding|Hospital Course|6459,6464|false|false|false|C0085639|Falls|falls
Event|Event|Hospital Course|6476,6478|false|false|false|||CT
Anatomy|Body Location or Region|Hospital Course|6486,6490|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6486,6490|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|Hospital Course|6486,6490|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6486,6490|false|false|false|C0876917|Procedure on head|head
Event|Event|Hospital Course|6491,6503|false|false|false|||demonstrated
Finding|Functional Concept|Hospital Course|6506,6510|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Event|Event|Hospital Course|6532,6536|false|false|false|||mass
Finding|Finding|Hospital Course|6532,6536|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|Hospital Course|6532,6536|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Hospital Course|6532,6536|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Finding|Hospital Course|6540,6544|false|false|false|C5575035|Well (answer to question)|well
Finding|Intellectual Product|Hospital Course|6555,6560|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|Hospital Course|6561,6567|false|false|false|||lesion
Finding|Finding|Hospital Course|6561,6567|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|Hospital Course|6561,6567|false|false|false|C0221198;C1546698|Lesion|lesion
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6585,6589|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|Hospital Course|6585,6589|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Finding|Functional Concept|Hospital Course|6597,6601|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Disorder|Injury or Poisoning|Hospital Course|6625,6630|false|false|false|C0000921|Accidental Falls|falls
Event|Event|Hospital Course|6625,6630|false|false|false|||falls
Finding|Finding|Hospital Course|6625,6630|false|false|false|C0085639|Falls|falls
Drug|Organic Chemical|Hospital Course|6636,6644|false|false|false|C0699129|Coumadin|coumadin
Drug|Pharmacologic Substance|Hospital Course|6636,6644|false|false|false|C0699129|Coumadin|coumadin
Event|Event|Hospital Course|6636,6644|false|false|false|||coumadin
Event|Event|Hospital Course|6650,6654|false|false|false|||held
Event|Event|Hospital Course|6666,6672|false|false|false|||placed
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6679,6686|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|Hospital Course|6679,6686|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|Hospital Course|6679,6686|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|Hospital Course|6679,6686|false|false|false|||insulin
Finding|Gene or Genome|Hospital Course|6679,6686|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|Hospital Course|6679,6686|false|false|false|C0202098|Insulin measurement|insulin
Event|Event|Hospital Course|6687,6694|false|false|false|||sliding
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6695,6700|false|false|false|C0222045|Integumentary scale|scale
Event|Activity|Hospital Course|6695,6700|false|false|false|C1947916|Scaling|scale
Finding|Conceptual Entity|Hospital Course|6695,6700|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Finding|Intellectual Product|Hospital Course|6695,6700|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Event|Event|Hospital Course|6720,6727|false|false|false|||concern
Finding|Idea or Concept|Hospital Course|6720,6727|false|false|false|C2699424|Concern|concern
Disorder|Disease or Syndrome|Hospital Course|6732,6744|false|true|false|C0020615|Hypoglycemia|hypoglycemia
Event|Event|Hospital Course|6732,6744|false|false|false|||hypoglycemia
Finding|Finding|Hospital Course|6732,6744|false|true|false|C5767385|Blood glucose below reference range (finding)|hypoglycemia
Event|Event|Hospital Course|6745,6757|false|false|false|||contributing
Event|Event|Hospital Course|6765,6777|false|false|false|||unsteadiness
Finding|Finding|Hospital Course|6765,6777|false|false|false|C0427108|General unsteadiness|unsteadiness
Event|Event|Hospital Course|6784,6787|false|false|false|||MRI
Finding|Gene or Genome|Hospital Course|6784,6787|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|Hospital Course|6784,6787|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|Hospital Course|6784,6787|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Anatomy|Body Location or Region|Hospital Course|6796,6800|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6796,6800|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|Hospital Course|6796,6800|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6796,6800|false|false|false|C0876917|Procedure on head|head
Event|Event|Hospital Course|6805,6813|false|false|false|||obtained
Event|Event|Hospital Course|6820,6829|false|false|false|||confirmed
Disorder|Neoplastic Process|Hospital Course|6832,6842|false|false|false|C0025286;C0281784|Benign Meningioma;Meningioma|meningioma
Event|Event|Hospital Course|6832,6842|false|false|false|||meningioma
Event|Event|Hospital Course|6844,6853|false|false|false|||overlying
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6860,6872|false|false|false|C0016733|frontal lobe|frontal lobe
Disorder|Neoplastic Process|Hospital Course|6860,6872|false|false|false|C0153635|malignant neoplasm of frontal lobe|frontal lobe
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6868,6872|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|Hospital Course|6868,6872|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Event|Event|Hospital Course|6889,6896|false|false|false|||infarct
Finding|Pathologic Function|Hospital Course|6889,6896|false|false|false|C0021308|Infarction|infarct
Event|Event|Hospital Course|6918,6923|false|false|false|||gyrus
Finding|Functional Concept|Hospital Course|6931,6935|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Functional Concept|Hospital Course|6964,6969|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Event|Event|Hospital Course|6977,6985|false|false|false|||weakness
Finding|Sign or Symptom|Hospital Course|6977,6985|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Finding|Finding|Hospital Course|6993,7002|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Idea or Concept|Hospital Course|6993,7002|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Intellectual Product|Hospital Course|6993,7002|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Pathologic Function|Hospital Course|6993,7002|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Phenomenon|Phenomenon or Process|Hospital Course|6993,7002|false|false|false|C0013956|Emergency Situation|emergency
Procedure|Health Care Activity|Hospital Course|6993,7002|false|false|false|C1553500|emergency encounter|emergency
Finding|Idea or Concept|Hospital Course|6993,7007|false|false|false|C1546435|Encounter Referral Source - emergency room|emergency room
Finding|Idea or Concept|Hospital Course|7012,7020|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Idea or Concept|Hospital Course|7021,7024|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|7021,7024|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|7034,7042|false|false|false|||weakness
Finding|Sign or Symptom|Hospital Course|7034,7042|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Finding|Intellectual Product|Hospital Course|7054,7064|false|false|false|C4554154|Completely - dosing instruction fragment|completely
Event|Event|Hospital Course|7065,7073|false|false|false|||resolved
Disorder|Mental or Behavioral Dysfunction|Hospital Course|7082,7091|false|false|false|C0009676|Confusion|confusion
Event|Event|Hospital Course|7082,7091|false|false|false|||confusion
Finding|Finding|Hospital Course|7082,7091|false|false|false|C0683369|Clouded consciousness|confusion
Event|Event|Hospital Course|7102,7108|false|false|false|||better
Finding|Idea or Concept|Hospital Course|7102,7108|false|false|false|C1550462|Observation Interpretation - better|better
Event|Event|Hospital Course|7122,7129|false|false|false|||consult
Procedure|Health Care Activity|Hospital Course|7122,7129|false|false|false|C0009818|Consultation|consult
Event|Event|Hospital Course|7134,7142|false|false|false|||obtained
Event|Event|Hospital Course|7155,7163|false|false|false|||appeared
Disorder|Disease or Syndrome|Hospital Course|7182,7188|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|Hospital Course|7182,7188|false|false|false|||stroke
Finding|Finding|Hospital Course|7182,7188|false|false|false|C5977286|Stroke (heart beat)|stroke
Event|Event|Hospital Course|7196,7199|false|false|false|||MRI
Finding|Gene or Genome|Hospital Course|7196,7199|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|Hospital Course|7196,7199|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|Hospital Course|7196,7199|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Event|Event|Hospital Course|7207,7218|false|false|false|||recommended
Event|Event|Hospital Course|7220,7230|false|false|false|||restarting
Drug|Organic Chemical|Hospital Course|7240,7248|false|false|false|C0699129|Coumadin|coumadin
Drug|Pharmacologic Substance|Hospital Course|7240,7248|false|false|false|C0699129|Coumadin|coumadin
Event|Event|Hospital Course|7240,7248|false|false|false|||coumadin
Event|Event|Hospital Course|7250,7257|false|false|false|||holding
Drug|Organic Chemical|Hospital Course|7262,7270|false|false|false|C0699512|Dilantin|dilantin
Drug|Pharmacologic Substance|Hospital Course|7262,7270|false|false|false|C0699512|Dilantin|dilantin
Event|Event|Hospital Course|7262,7270|false|false|false|||dilantin
Event|Activity|Hospital Course|7275,7283|false|false|false|C1283174||checking
Event|Event|Hospital Course|7275,7283|false|false|false|||checking
Event|Event|Hospital Course|7288,7291|false|false|false|||EEG
Procedure|Diagnostic Procedure|Hospital Course|7288,7291|false|false|false|C0013819|Electroencephalography|EEG
Event|Event|Hospital Course|7325,7334|false|false|false|||inpatient
Finding|Idea or Concept|Hospital Course|7325,7334|false|false|false|C1548438;C1549404|Patient Class - Inpatient;Referral category - Inpatient|inpatient
Procedure|Health Care Activity|Hospital Course|7325,7334|false|false|false|C1555324|inpatient encounter|inpatient
Event|Event|Hospital Course|7365,7369|false|false|false|||echo
Procedure|Health Care Activity|Hospital Course|7365,7369|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7365,7369|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7377,7380|false|false|false|C1609165|tocilizumab|MRA
Drug|Immunologic Factor|Hospital Course|7377,7380|false|false|false|C1609165|tocilizumab|MRA
Drug|Pharmacologic Substance|Hospital Course|7377,7380|false|false|false|C1609165|tocilizumab|MRA
Event|Event|Hospital Course|7377,7380|false|false|false|||MRA
Lab|Laboratory or Test Result|Hospital Course|7377,7380|false|false|false|C3891069|MRI-Based Angiogram|MRA
Procedure|Diagnostic Procedure|Hospital Course|7377,7380|false|false|false|C0243032|Magnetic Resonance Angiography|MRA
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7388,7393|false|false|false|C0006104;C4266577|Brain;Head>Brain|brain
Disorder|Disease or Syndrome|Hospital Course|7388,7393|false|false|false|C0006111|Brain Diseases|brain
Anatomy|Body Location or Region|Hospital Course|7398,7402|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|Hospital Course|7398,7402|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|Hospital Course|7398,7402|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Finding|Finding|Hospital Course|7414,7420|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|7414,7420|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Pathologic Function|Hospital Course|7421,7428|false|true|false|C0013922|Embolism|embolic
Event|Event|Hospital Course|7429,7435|false|false|false|||nature
Finding|Functional Concept|Hospital Course|7429,7435|false|false|false|C0349590;C1262865|Nature;Natures|nature
Finding|Idea or Concept|Hospital Course|7429,7435|false|false|false|C0349590;C1262865|Nature;Natures|nature
Disorder|Disease or Syndrome|Hospital Course|7443,7450|false|false|false|C0038454|Cerebrovascular accident|strokes
Event|Event|Hospital Course|7443,7450|false|false|false|||strokes
Event|Event|Hospital Course|7469,7472|false|false|false|||see
Finding|Functional Concept|Hospital Course|7496,7502|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Anatomy|Body Location or Region|Hospital Course|7503,7507|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7503,7507|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|Hospital Course|7503,7507|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7503,7507|false|false|false|C0876917|Procedure on head|head
Procedure|Diagnostic Procedure|Hospital Course|7503,7511|false|false|false|C0412674|MRI of head|head MRI
Event|Event|Hospital Course|7508,7511|false|false|false|||MRI
Finding|Gene or Genome|Hospital Course|7508,7511|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|Hospital Course|7508,7511|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|Hospital Course|7508,7511|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Event|Event|Hospital Course|7523,7526|false|false|false|||saw
Disorder|Disease or Syndrome|Hospital Course|7539,7547|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|diabetes
Event|Event|Hospital Course|7548,7557|false|false|false|||managment
Event|Event|Hospital Course|7563,7574|false|false|false|||recommended
Event|Event|Hospital Course|7575,7583|false|false|false|||changing
Drug|Organic Chemical|Hospital Course|7588,7597|true|false|false|C0017642|glipizide|glipizide
Drug|Pharmacologic Substance|Hospital Course|7588,7597|true|false|false|C0017642|glipizide|glipizide
Event|Event|Hospital Course|7588,7597|true|false|false|||glipizide
Disorder|Mental or Behavioral Dysfunction|Hospital Course|7604,7607|true|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7604,7607|true|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|7604,7607|true|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|7604,7607|true|false|false|||BID
Finding|Gene or Genome|Hospital Course|7604,7607|true|false|false|C1332410|BID gene|BID
Event|Event|Hospital Course|7618,7626|true|false|false|||starting
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7627,7634|true|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|Hospital Course|7627,7634|true|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|Hospital Course|7627,7634|true|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|Hospital Course|7627,7634|true|false|false|||insulin
Finding|Gene or Genome|Hospital Course|7627,7634|true|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|Hospital Course|7627,7634|true|false|false|C0202098|Insulin measurement|insulin
Drug|Organic Chemical|Hospital Course|7640,7646|false|false|false|C0242209|Sugars|sugars
Drug|Pharmacologic Substance|Hospital Course|7640,7646|false|false|false|C0242209|Sugars|sugars
Event|Event|Hospital Course|7640,7646|false|false|false|||sugars
Procedure|Laboratory Procedure|Hospital Course|7640,7646|false|false|false|C2239291|sugars (lab test)|sugars
Finding|Finding|Hospital Course|7652,7656|false|false|false|C5575035|Well (answer to question)|well
Event|Event|Hospital Course|7657,7667|false|false|false|||controlled
Event|Event|Hospital Course|7708,7716|true|false|false|||episodes
Disorder|Disease or Syndrome|Hospital Course|7720,7732|true|false|false|C0020615|Hypoglycemia|hypoglycemia
Event|Event|Hospital Course|7720,7732|true|false|false|||hypoglycemia
Finding|Finding|Hospital Course|7720,7732|true|false|false|C5767385|Blood glucose below reference range (finding)|hypoglycemia
Event|Event|Hospital Course|7753,7763|false|false|false|||standpoing
Finding|Idea or Concept|Hospital Course|7765,7773|false|false|false|C4288901|In-House|in-house
Event|Event|Hospital Course|7787,7791|false|false|false|||well
Finding|Finding|Hospital Course|7787,7791|false|false|false|C5575035|Well (answer to question)|well
Event|Event|Hospital Course|7797,7806|false|false|false|||resultion
Finding|Functional Concept|Hospital Course|7815,7820|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Finding|Finding|Hospital Course|7815,7835|false|false|false|C0457435|Right hemiparesis|right sided weakness
Event|Event|Hospital Course|7827,7835|false|false|false|||weakness
Finding|Sign or Symptom|Hospital Course|7827,7835|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Finding|Finding|Hospital Course|7849,7861|false|false|false|C0427108|General unsteadiness|unsteadiness
Event|Event|Hospital Course|7862,7871|false|false|false|||continued
Finding|Idea or Concept|Hospital Course|7862,7871|false|false|false|C0549178|Continuous|continued
Event|Event|Hospital Course|7880,7886|false|false|false|||needed
Attribute|Clinical Attribute|Hospital Course|7887,7894|false|false|false|C1317973|Support - dental|support
Drug|Organic Chemical|Hospital Course|7887,7894|false|false|false|C1171411|Support brand of multivitamin|support
Drug|Pharmacologic Substance|Hospital Course|7887,7894|false|false|false|C1171411|Support brand of multivitamin|support
Drug|Vitamin|Hospital Course|7887,7894|false|false|false|C1171411|Support brand of multivitamin|support
Event|Event|Hospital Course|7887,7894|false|false|false|||support
Finding|Conceptual Entity|Hospital Course|7887,7894|false|false|false|C1521721|Supportive assistance|support
Procedure|Health Care Activity|Hospital Course|7887,7894|false|false|false|C0344211|Supportive care|support
Event|Event|Hospital Course|7901,7911|false|false|false|||ambulating
Event|Event|Hospital Course|7919,7930|false|false|false|||recommended
Event|Event|Hospital Course|7934,7936|false|false|false|||go
Finding|Idea or Concept|Hospital Course|7948,7952|false|false|false|C0233324;C1705313|Term (lexical);Term Birth|term
Finding|Organism Function|Hospital Course|7948,7952|false|false|false|C0233324;C1705313|Term (lexical);Term Birth|term
Event|Event|Hospital Course|7953,7958|false|false|false|||rehab
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7953,7958|false|false|false|C0034991|Rehabilitation therapy|rehab
Event|Event|Hospital Course|7972,7978|false|false|false|||better
Finding|Idea or Concept|Hospital Course|7972,7978|false|false|false|C1550462|Observation Interpretation - better|better
Event|Event|Hospital Course|7980,7984|false|false|false|||able
Finding|Finding|Hospital Course|7980,7984|false|false|false|C1299581|Able (qualifier value)|able
Event|Event|Hospital Course|7988,7995|false|false|false|||compete
Event|Event|Hospital Course|7996,8005|false|false|false|||transfers
Finding|Finding|Hospital Course|7996,8005|false|false|false|C0728827|transfers|transfers
Event|Event|Hospital Course|8010,8018|false|false|false|||ambulate
Finding|Finding|Hospital Course|8010,8018|false|false|false|C4036205|Ambulate|ambulate
Event|Event|Hospital Course|8043,8049|false|false|false|||follow
Event|Event|Hospital Course|8058,8067|false|false|false|||neurology
Event|Event|Hospital Course|8072,8084|false|false|false|||neurosurgery
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8072,8084|false|false|false|C0524850|Neurosurgical Procedures|neurosurgery
Event|Event|Hospital Course|8088,8095|false|false|false|||discuss
Disorder|Disease or Syndrome|Hospital Course|8103,8107|false|false|false|C0339510|Vitelliform Macular Dystrophy|best
Event|Event|Hospital Course|8103,8107|false|false|false|||best
Finding|Gene or Genome|Hospital Course|8103,8107|false|false|false|C1826421;C5781213|BEST1 gene;BEST1 wt Allele|best
Event|Event|Hospital Course|8109,8115|false|false|false|||manage
Finding|Functional Concept|Hospital Course|8120,8128|false|false|false|C0475224|Ischemic|ischemic
Disorder|Disease or Syndrome|Hospital Course|8120,8136|false|false|false|C0948008|Ischemic stroke|ischemic strokes
Disorder|Disease or Syndrome|Hospital Course|8129,8136|false|false|false|C0038454|Cerebrovascular accident|strokes
Event|Event|Hospital Course|8129,8136|false|false|false|||strokes
Event|Event|Hospital Course|8141,8148|false|false|false|||address
Disorder|Neoplastic Process|Hospital Course|8153,8163|false|false|false|C0025286;C0281784|Benign Meningioma;Meningioma|meningioma
Event|Event|Hospital Course|8153,8163|false|false|false|||meningioma
Attribute|Clinical Attribute|Hospital Course|8182,8193|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|8182,8193|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|8182,8193|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|8182,8193|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|8182,8206|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|8197,8206|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|8197,8206|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Organic Chemical|Hospital Course|8208,8216|false|false|false|C0699129|Coumadin|Coumadin
Drug|Pharmacologic Substance|Hospital Course|8208,8216|false|false|false|C0699129|Coumadin|Coumadin
Event|Event|Hospital Course|8208,8216|false|false|false|||Coumadin
Event|Event|Hospital Course|8220,8221|false|false|false|||'
Drug|Organic Chemical|Hospital Course|8223,8230|false|false|false|C0722725|Prandin|prandin
Drug|Pharmacologic Substance|Hospital Course|8223,8230|false|false|false|C0722725|Prandin|prandin
Event|Event|Hospital Course|8223,8230|false|false|false|||prandin
Drug|Organic Chemical|Hospital Course|8239,8248|false|false|false|C0017642|glipizide|glipizide
Drug|Pharmacologic Substance|Hospital Course|8239,8248|false|false|false|C0017642|glipizide|glipizide
Event|Event|Hospital Course|8239,8248|false|false|false|||glipizide
Drug|Organic Chemical|Hospital Course|8254,8264|false|false|false|C0022251|isosorbide|isosorbide
Drug|Pharmacologic Substance|Hospital Course|8254,8264|false|false|false|C0022251|isosorbide|isosorbide
Event|Event|Hospital Course|8254,8264|false|false|false|||isosorbide
Event|Event|Hospital Course|8266,8275|false|false|false|||dinitrate
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8282,8292|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|Hospital Course|8282,8292|false|false|false|C0065374|lisinopril|lisinopril
Event|Event|Hospital Course|8282,8292|false|false|false|||lisinopril
Drug|Organic Chemical|Hospital Course|8297,8308|false|false|false|C0002144|allopurinol|allopurinol
Drug|Pharmacologic Substance|Hospital Course|8297,8308|false|false|false|C0002144|allopurinol|allopurinol
Event|Event|Hospital Course|8297,8308|false|false|false|||allopurinol
Drug|Organic Chemical|Hospital Course|8314,8323|false|false|false|C0076840|torsemide|torsemide
Drug|Pharmacologic Substance|Hospital Course|8314,8323|false|false|false|C0076840|torsemide|torsemide
Event|Event|Hospital Course|8314,8323|false|false|false|||torsemide
Drug|Organic Chemical|Hospital Course|8328,8338|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|Hospital Course|8328,8338|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|Hospital Course|8328,8338|false|false|false|||metoprolol
Drug|Organic Chemical|Hospital Course|8346,8353|false|false|false|C0593906|Lipitor|lipitor
Drug|Pharmacologic Substance|Hospital Course|8346,8353|false|false|false|C0593906|Lipitor|lipitor
Event|Event|Hospital Course|8346,8353|false|false|false|||lipitor
Event|Event|Hospital Course|8361,8370|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|8361,8370|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|8361,8370|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|8361,8370|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|8361,8370|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|8361,8382|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|8371,8382|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|8371,8382|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|8371,8382|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|8371,8382|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|8387,8397|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|Hospital Course|8387,8397|false|false|false|C0022251|isosorbide|Isosorbide
Event|Event|Hospital Course|8387,8397|false|false|false|||Isosorbide
Drug|Organic Chemical|Hospital Course|8387,8407|false|false|false|C0022252|isosorbide dinitrate|Isosorbide Dinitrate
Drug|Pharmacologic Substance|Hospital Course|8387,8407|false|false|false|C0022252|isosorbide dinitrate|Isosorbide Dinitrate
Event|Event|Hospital Course|8398,8407|false|false|false|||Dinitrate
Drug|Biomedical or Dental Material|Hospital Course|8414,8420|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|8434,8440|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|8434,8440|false|false|false|||Tablet
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8444,8447|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8444,8447|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8444,8447|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|8444,8447|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|8444,8447|false|false|false|C1332410|BID gene|BID
Finding|Finding|Hospital Course|8450,8457|false|false|false|C4035627|2 times|2 times
Disorder|Disease or Syndrome|Hospital Course|8452,8457|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|Hospital Course|8460,8463|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|8460,8463|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8471,8481|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|Hospital Course|8471,8481|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Biomedical or Dental Material|Hospital Course|8488,8494|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|8508,8514|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|8508,8514|false|false|false|||Tablet
Drug|Organic Chemical|Hospital Course|8539,8549|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|Hospital Course|8539,8549|false|false|false|C0025859|metoprolol|Metoprolol
Event|Event|Hospital Course|8539,8549|false|false|false|||Metoprolol
Drug|Organic Chemical|Hospital Course|8539,8558|false|false|false|C0700548|metoprolol tartrate|Metoprolol Tartrate
Drug|Pharmacologic Substance|Hospital Course|8539,8558|false|false|false|C0700548|metoprolol tartrate|Metoprolol Tartrate
Drug|Organic Chemical|Hospital Course|8550,8558|false|false|false|C0039328;C0144544|Tartrates;tartrate|Tartrate
Drug|Pharmacologic Substance|Hospital Course|8550,8558|false|false|false|C0039328;C0144544|Tartrates;tartrate|Tartrate
Drug|Biomedical or Dental Material|Hospital Course|8565,8571|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|8585,8591|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|8585,8591|false|false|false|||Tablet
Event|Event|Hospital Course|8595,8598|false|false|false|||TID
Finding|Finding|Hospital Course|8601,8608|false|false|false|C4035626|3 times|3 times
Disorder|Disease or Syndrome|Hospital Course|8603,8608|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Event|Event|Hospital Course|8603,8608|false|false|false|||times
Finding|Idea or Concept|Hospital Course|8611,8614|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|8611,8614|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|8622,8633|false|false|false|C0074554|simvastatin|Simvastatin
Drug|Pharmacologic Substance|Hospital Course|8622,8633|false|false|false|C0074554|simvastatin|Simvastatin
Drug|Biomedical or Dental Material|Hospital Course|8640,8646|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|8660,8666|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|8667,8669|false|false|false|||PO
Drug|Organic Chemical|Hospital Course|8691,8702|false|false|false|C0002144|allopurinol|Allopurinol
Drug|Pharmacologic Substance|Hospital Course|8691,8702|false|false|false|C0002144|allopurinol|Allopurinol
Drug|Biomedical or Dental Material|Hospital Course|8710,8716|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|8730,8736|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|8730,8736|false|false|false|||Tablet
Drug|Hazardous or Poisonous Substance|Hospital Course|8761,8769|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|Hospital Course|8761,8769|false|false|false|C0043031|warfarin|Warfarin
Drug|Pharmacologic Substance|Hospital Course|8761,8769|false|false|false|C0043031|warfarin|Warfarin
Drug|Biomedical or Dental Material|Hospital Course|8777,8783|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|8797,8803|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|8804,8806|false|false|false|||PO
Drug|Organic Chemical|Hospital Course|8834,8843|false|false|false|C0076840|torsemide|Torsemide
Drug|Pharmacologic Substance|Hospital Course|8834,8843|false|false|false|C0076840|torsemide|Torsemide
Drug|Biomedical or Dental Material|Hospital Course|8849,8855|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|8869,8875|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|8869,8875|false|false|false|||Tablet
Drug|Organic Chemical|Hospital Course|8899,8908|false|false|false|C0017642|glipizide|Glipizide
Drug|Pharmacologic Substance|Hospital Course|8899,8908|false|false|false|C0017642|glipizide|Glipizide
Drug|Biomedical or Dental Material|Hospital Course|8915,8921|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|8935,8941|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|8935,8941|false|false|false|||Tablet
Event|Event|Hospital Course|8942,8944|false|false|false|||PO
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8945,8948|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8945,8948|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8945,8948|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|8945,8948|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|8945,8948|false|false|false|C1332410|BID gene|BID
Finding|Finding|Hospital Course|8950,8957|false|false|false|C4035627|2 times|2 times
Disorder|Disease or Syndrome|Hospital Course|8952,8957|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Event|Event|Hospital Course|8952,8957|false|false|false|||times
Finding|Idea or Concept|Hospital Course|8961,8964|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|8961,8964|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|8972,8981|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|8972,8981|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|8972,8981|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|8972,8981|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|8972,8981|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|8972,8993|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|8972,8993|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|8982,8993|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|8982,8993|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|8982,8993|false|false|false|C0184758|Patient disposition|Disposition
Finding|Finding|Hospital Course|8995,9003|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|8995,9003|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Procedure|Health Care Activity|Hospital Course|8995,9008|false|false|false|C0023977|long-term care|Extended Care
Event|Activity|Hospital Course|9004,9008|false|false|false|C1947933|care activity|Care
Event|Event|Hospital Course|9004,9008|false|false|false|||Care
Finding|Finding|Hospital Course|9004,9008|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Hospital Course|9004,9008|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Event|Event|Hospital Course|9011,9019|false|false|false|||Facility
Finding|Intellectual Product|Hospital Course|9011,9019|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|Hospital Course|9025,9034|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|9025,9034|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|9025,9034|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|9025,9034|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|9025,9034|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|9025,9044|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|9035,9044|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|9035,9044|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|9035,9044|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|9035,9044|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|9035,9044|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Functional Concept|Hospital Course|9046,9050|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Disorder|Neoplastic Process|Hospital Course|9059,9069|false|false|false|C0025286;C0281784|Benign Meningioma;Meningioma|meningioma
Event|Event|Hospital Course|9059,9069|false|false|false|||meningioma
Finding|Functional Concept|Hospital Course|9071,9075|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Event|Event|Hospital Course|9095,9102|false|false|false|||infarct
Finding|Pathologic Function|Hospital Course|9095,9102|false|false|false|C0021308|Infarction|infarct
Disorder|Disease or Syndrome|Hospital Course|9105,9113|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|Diabetes
Event|Event|Hospital Course|9105,9113|false|false|false|||Diabetes
Finding|Mental Process|Discharge Condition|9138,9144|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|9138,9151|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|9138,9151|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|9145,9151|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|9145,9151|false|false|false|C1546481|What subject filter - Status|Status
Disorder|Mental or Behavioral Dysfunction|Discharge Condition|9153,9161|false|false|false|C0009676|Confusion|Confused
Event|Event|Discharge Condition|9153,9161|false|false|false|||Confused
Finding|Finding|Discharge Condition|9153,9161|false|false|false|C0683369;C1547301|Clouded consciousness;Precaution Code - Confused|Confused
Finding|Intellectual Product|Discharge Condition|9153,9161|false|false|false|C0683369;C1547301|Clouded consciousness;Precaution Code - Confused|Confused
Event|Event|Discharge Condition|9175,9180|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|9175,9197|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|9175,9197|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|9184,9197|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|9184,9197|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|9184,9197|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|9199,9204|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|9199,9204|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|9199,9204|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|9199,9204|false|false|false|||Alert
Finding|Finding|Discharge Condition|9199,9204|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|9199,9204|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|9199,9204|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|9209,9220|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|9209,9220|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|9222,9230|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|9222,9230|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|9222,9230|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|9231,9237|false|false|false|C5889824||Status
Event|Event|Discharge Condition|9231,9237|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|9231,9237|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|Discharge Condition|9239,9249|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|9239,9249|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|9239,9249|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|9239,9249|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|9252,9260|false|false|false|||requires
Event|Event|Discharge Condition|9261,9271|false|false|false|||assistance
Finding|Social Behavior|Discharge Condition|9261,9271|false|false|false|C0018896|Helping Behavior|assistance
Drug|Amino Acid, Peptide, or Protein|Discharge Condition|9275,9278|false|false|false|C1454018|AICDA protein, human|aid
Drug|Enzyme|Discharge Condition|9275,9278|false|false|false|C1454018|AICDA protein, human|aid
Event|Event|Discharge Condition|9275,9278|false|false|false|||aid
Finding|Gene or Genome|Discharge Condition|9275,9278|false|false|false|C1421876;C3540469|AICDA gene;AICDA wt Allele|aid
Procedure|Therapeutic or Preventive Procedure|Discharge Condition|9275,9278|false|false|false|C0021588;C0280108|AID - Artificial insemination by donor;dacarbazine/doxorubicin/ifosfamide protocol|aid
Event|Event|Discharge Condition|9280,9286|false|false|false|||walker
Event|Event|Discharge Instructions|9336,9340|false|false|false|||take
Drug|Organic Chemical|Discharge Instructions|9346,9354|false|false|false|C0699129|Coumadin|coumadin
Drug|Pharmacologic Substance|Discharge Instructions|9346,9354|false|false|false|C0699129|Coumadin|coumadin
Event|Event|Discharge Instructions|9346,9354|false|false|false|||coumadin
Event|Event|Discharge Instructions|9358,9368|false|false|false|||prescribed
Event|Event|Discharge Instructions|9381,9385|true|false|false|||need
Attribute|Clinical Attribute|Discharge Instructions|9399,9410|true|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|9399,9410|true|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|9399,9410|true|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|9399,9410|true|false|false|C4284232|Medications|medications
Event|Event|Discharge Instructions|9434,9440|false|false|false|||follow
Event|Event|Discharge Instructions|9469,9475|false|false|false|||listed
Event|Event|Discharge Instructions|9492,9496|false|false|false|||need
Finding|Functional Concept|Discharge Instructions|9499,9505|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|Discharge Instructions|9499,9505|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|Discharge Instructions|9499,9508|false|false|false|C0589120|Follow-up status|follow up
Procedure|Health Care Activity|Discharge Instructions|9499,9508|false|false|false|C1522577|follow-up|follow up
Event|Event|Discharge Instructions|9509,9512|false|false|false|||MRI
Finding|Gene or Genome|Discharge Instructions|9509,9512|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|Discharge Instructions|9509,9512|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|Discharge Instructions|9509,9512|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Event|Event|Discharge Instructions|9516,9524|false|false|false|||evaluate
Disorder|Disease or Syndrome|Discharge Instructions|9536,9542|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|Discharge Instructions|9536,9542|false|false|false|||stroke
Finding|Finding|Discharge Instructions|9536,9542|false|false|false|C5977286|Stroke (heart beat)|stroke
Finding|Functional Concept|Discharge Instructions|9558,9562|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|9576,9581|false|false|false|C0006104;C4266577|Brain;Head>Brain|brain
Disorder|Disease or Syndrome|Discharge Instructions|9576,9581|false|false|false|C0006111|Brain Diseases|brain
Attribute|Clinical Attribute|Discharge Instructions|9593,9604|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|9593,9604|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|9593,9604|false|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|9593,9604|false|false|false|C4284232|Medications|medications
Event|Event|Discharge Instructions|9608,9618|false|false|false|||prescribed
Event|Event|Discharge Instructions|9623,9629|false|false|false|||follow
Finding|Intellectual Product|Discharge Instructions|9652,9656|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|Discharge Instructions|9660,9665|false|false|false|||check
Finding|Classification|Discharge Instructions|9671,9678|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|Discharge Instructions|9671,9678|false|false|false|C3812897|General medical service|General
Finding|Idea or Concept|Discharge Instructions|9671,9691|false|false|false|C1549999|General Instructions|General Instructions
Attribute|Clinical Attribute|Discharge Instructions|9679,9691|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|9679,9691|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|9679,9691|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Finding|Idea or Concept|Discharge Instructions|9692,9703|false|false|false|C0870705;C1533716;C1561527;C1561528|Acknowledgement Detail Type - Information;Error severity - Information;Information;control act - information|Information
Finding|Intellectual Product|Discharge Instructions|9692,9703|false|false|false|C0870705;C1533716;C1561527;C1561528|Acknowledgement Detail Type - Information;Error severity - Information;Information;control act - information|Information
Event|Event|Discharge Instructions|9705,9709|false|false|false|||Take
Attribute|Clinical Attribute|Discharge Instructions|9715,9719|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|9715,9719|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|9715,9719|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|9715,9719|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Hazardous or Poisonous Substance|Discharge Instructions|9715,9728|false|false|false|C0002771|Analgesics|pain medicine
Drug|Organic Chemical|Discharge Instructions|9715,9728|false|false|false|C0002771|Analgesics|pain medicine
Drug|Pharmacologic Substance|Discharge Instructions|9715,9728|false|false|false|C0002771|Analgesics|pain medicine
Drug|Pharmacologic Substance|Discharge Instructions|9720,9728|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Event|Event|Discharge Instructions|9720,9728|false|false|false|||medicine
Event|Event|Discharge Instructions|9732,9742|false|false|false|||prescribed
Event|Event|Discharge Instructions|9745,9753|false|false|false|||Exercise
Finding|Daily or Recreational Activity|Discharge Instructions|9745,9753|false|false|false|C0015259|Exercise|Exercise
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|9745,9753|false|false|false|C1522704|Exercise Pain Management|Exercise
Event|Event|Discharge Instructions|9764,9771|false|false|false|||limited
Event|Event|Discharge Instructions|9775,9782|false|false|false|||walking
Finding|Daily or Recreational Activity|Discharge Instructions|9775,9782|false|true|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Finding|Finding|Discharge Instructions|9775,9782|false|true|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Finding|Sign or Symptom|Discharge Instructions|9775,9782|false|true|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Event|Activity|Discharge Instructions|9787,9794|true|false|false|C0206244|Lifting|lifting
Event|Event|Discharge Instructions|9787,9794|true|false|false|||lifting
Event|Event|Discharge Instructions|9796,9805|true|false|false|||straining
Finding|Physiologic Function|Discharge Instructions|9796,9805|true|false|false|C0442694|Straining (finding)|straining
Disorder|Disease or Syndrome|Discharge Instructions|9821,9828|false|false|false|C0011119|Decompression Sickness|bending
Event|Event|Discharge Instructions|9821,9828|false|false|false|||bending
Finding|Finding|Discharge Instructions|9821,9828|false|false|false|C0700231;C2584296|Bending - Changing basic body position;Does bend|bending
Finding|Physiologic Function|Discharge Instructions|9821,9828|false|false|false|C0700231;C2584296|Bending - Changing basic body position;Does bend|bending
Event|Event|Discharge Instructions|9831,9839|false|false|false|||Increase
Event|Event|Discharge Instructions|9845,9851|false|false|false|||intake
Finding|Functional Concept|Discharge Instructions|9845,9851|false|false|false|C1512806|Intake|intake
Procedure|Health Care Activity|Discharge Instructions|9845,9851|false|false|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|intake
Drug|Substance|Discharge Instructions|9855,9861|false|false|false|C0302908|Liquid substance|fluids
Event|Event|Discharge Instructions|9855,9861|false|false|false|||fluids
Finding|Body Substance|Discharge Instructions|9855,9861|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|9855,9861|false|false|false|C0016286|Fluid Therapy|fluids
Anatomy|Tissue|Discharge Instructions|9866,9871|false|false|false|C1304649|Tissue fiber|fiber
Drug|Organic Chemical|Discharge Instructions|9866,9871|false|false|false|C0225326;C1321801|Fiber brand of calcium polycarbophil;fiber|fiber
Drug|Pharmacologic Substance|Discharge Instructions|9866,9871|false|false|false|C0225326;C1321801|Fiber brand of calcium polycarbophil;fiber|fiber
Drug|Hazardous or Poisonous Substance|Discharge Instructions|9876,9884|false|false|false|C0027415|Narcotics|narcotic
Drug|Pharmacologic Substance|Discharge Instructions|9876,9884|false|false|false|C0027415|Narcotics|narcotic
Attribute|Clinical Attribute|Discharge Instructions|9885,9889|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|9885,9889|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|9885,9889|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|9885,9889|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Pharmacologic Substance|Discharge Instructions|9891,9899|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Event|Event|Discharge Instructions|9891,9899|false|false|false|||medicine
Event|Event|Discharge Instructions|9904,9909|false|false|false|||cause
Event|Event|Discharge Instructions|9910,9922|false|false|false|||constipation
Finding|Sign or Symptom|Discharge Instructions|9910,9922|false|false|false|C0009806|Constipation|constipation
Event|Event|Discharge Instructions|9937,9946|false|false|false|||recommend
Event|Event|Discharge Instructions|9947,9953|false|false|false|||taking
Drug|Pharmacologic Substance|Discharge Instructions|9958,9974|false|false|false|C0013231|Drugs, Non-Prescription|over the counter
Drug|Hazardous or Poisonous Substance|Discharge Instructions|9967,9974|false|false|false|C0702263|Counter brand of Terbufos|counter
Drug|Organic Chemical|Discharge Instructions|9967,9974|false|false|false|C0702263|Counter brand of Terbufos|counter
Finding|Body Substance|Discharge Instructions|9975,9980|false|false|false|C0015733|Feces|stool
Drug|Organic Chemical|Discharge Instructions|9975,9989|false|false|false|C0301470;C1154263|Stool Softener;Stool Softener brand of docusate sodium|stool softener
Drug|Pharmacologic Substance|Discharge Instructions|9975,9989|false|false|false|C0301470;C1154263|Stool Softener;Stool Softener brand of docusate sodium|stool softener
Event|Event|Discharge Instructions|9981,9989|false|false|false|||softener
Drug|Organic Chemical|Discharge Instructions|9999,10007|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Discharge Instructions|9999,10007|false|false|false|C1692318|docusate|Docusate
Drug|Organic Chemical|Discharge Instructions|10009,10015|false|false|false|C0282139|Colace|Colace
Drug|Pharmacologic Substance|Discharge Instructions|10009,10015|false|false|false|C0282139|Colace|Colace
Drug|Hazardous or Poisonous Substance|Discharge Instructions|10031,10039|false|false|false|C0027415|Narcotics|narcotic
Drug|Pharmacologic Substance|Discharge Instructions|10031,10039|false|false|false|C0027415|Narcotics|narcotic
Attribute|Clinical Attribute|Discharge Instructions|10040,10044|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|10040,10044|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|10040,10044|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|10040,10044|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Pharmacologic Substance|Discharge Instructions|10045,10055|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Discharge Instructions|10045,10055|false|false|false|||medication
Finding|Intellectual Product|Discharge Instructions|10045,10055|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Discharge Instructions|10065,10073|true|false|false|||directed
Event|Event|Discharge Instructions|10082,10088|true|false|false|||doctor
Finding|Intellectual Product|Discharge Instructions|10082,10088|true|false|false|C2348314|Doctor - Title|doctor
Event|Event|Discharge Instructions|10097,10101|true|false|false|||take
Drug|Pharmacologic Substance|Discharge Instructions|10107,10124|true|false|false|C0003209|Anti-Inflammatory Agents|anti-inflammatory
Drug|Pharmacologic Substance|Discharge Instructions|10125,10134|true|false|false|C0013227|Pharmaceutical Preparations|medicines
Event|Event|Discharge Instructions|10125,10134|true|false|false|||medicines
Drug|Organic Chemical|Discharge Instructions|10143,10149|true|false|false|C0699203|Motrin|Motrin
Drug|Pharmacologic Substance|Discharge Instructions|10143,10149|true|false|false|C0699203|Motrin|Motrin
Drug|Organic Chemical|Discharge Instructions|10151,10158|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Discharge Instructions|10151,10158|false|false|false|C0004057|aspirin|Aspirin
Event|Event|Discharge Instructions|10151,10158|false|false|false|||Aspirin
Drug|Organic Chemical|Discharge Instructions|10160,10165|false|false|false|C0593507|Advil|Advil
Drug|Pharmacologic Substance|Discharge Instructions|10160,10165|false|false|false|C0593507|Advil|Advil
Event|Event|Discharge Instructions|10160,10165|false|false|false|||Advil
Finding|Gene or Genome|Discharge Instructions|10160,10165|false|false|false|C1422473|AVIL gene|Advil
Drug|Organic Chemical|Discharge Instructions|10172,10181|false|false|false|C0020740|ibuprofen|Ibuprofen
Drug|Pharmacologic Substance|Discharge Instructions|10172,10181|false|false|false|C0020740|ibuprofen|Ibuprofen
Finding|Idea or Concept|Discharge Instructions|10182,10185|false|false|false|C1548556|Etc.|etc
Event|Event|Discharge Instructions|10208,10212|false|false|false|||sent
Event|Event|Discharge Instructions|10213,10217|false|false|false|||home
Finding|Idea or Concept|Discharge Instructions|10213,10217|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Discharge Instructions|10213,10217|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Discharge Instructions|10213,10217|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Discharge Instructions|10221,10228|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Drug|Pharmacologic Substance|Discharge Instructions|10221,10228|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Drug|Pharmacologic Substance|Discharge Instructions|10229,10239|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Discharge Instructions|10229,10239|false|false|false|||medication
Finding|Intellectual Product|Discharge Instructions|10229,10239|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Discharge Instructions|10246,10250|false|false|false|||sure
Finding|Intellectual Product|Discharge Instructions|10246,10250|false|false|false|C4724437|SURE Test|sure
Event|Event|Discharge Instructions|10260,10266|false|false|false|||taking
Drug|Pharmacologic Substance|Discharge Instructions|10269,10279|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Discharge Instructions|10269,10279|false|false|false|||medication
Finding|Intellectual Product|Discharge Instructions|10269,10279|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Discharge Instructions|10283,10290|false|false|false|||protect
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|10296,10303|false|false|false|C0038351;C3714551;C4266636|Abdomen>Stomach;Stomach;Stomach structure|stomach
Disorder|Disease or Syndrome|Discharge Instructions|10296,10303|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Disorder|Neoplastic Process|Discharge Instructions|10296,10303|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Event|Event|Discharge Instructions|10296,10303|false|false|false|||stomach
Finding|Finding|Discharge Instructions|10296,10303|false|false|false|C0577027|Stomach problem|stomach
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10296,10303|false|false|false|C0872393|Procedure on stomach|stomach
Drug|Organic Chemical|Discharge Instructions|10305,10313|false|false|false|C0700777|Prilosec|Prilosec
Drug|Pharmacologic Substance|Discharge Instructions|10305,10313|false|false|false|C0700777|Prilosec|Prilosec
Drug|Organic Chemical|Discharge Instructions|10316,10324|false|false|false|C0876139|Protonix|Protonix
Drug|Pharmacologic Substance|Discharge Instructions|10316,10324|false|false|false|C0876139|Protonix|Protonix
Drug|Organic Chemical|Discharge Instructions|10329,10335|false|false|false|C0678119|Pepcid|Pepcid
Drug|Pharmacologic Substance|Discharge Instructions|10329,10335|false|false|false|C0678119|Pepcid|Pepcid
Event|Event|Discharge Instructions|10329,10335|false|false|false|||Pepcid
Attribute|Clinical Attribute|Discharge Instructions|10347,10358|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|10347,10358|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|10347,10358|false|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|10347,10358|false|false|false|C4284232|Medications|medications
Event|Event|Discharge Instructions|10363,10368|false|false|false|||cause
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|10369,10376|false|false|false|C0038351;C3714551;C4266636|Abdomen>Stomach;Stomach;Stomach structure|stomach
Disorder|Disease or Syndrome|Discharge Instructions|10369,10376|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Disorder|Neoplastic Process|Discharge Instructions|10369,10376|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Event|Event|Discharge Instructions|10369,10376|false|false|false|||stomach
Finding|Finding|Discharge Instructions|10369,10376|false|false|false|C0577027|Stomach problem|stomach
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10369,10376|false|false|false|C0872393|Procedure on stomach|stomach
Event|Event|Discharge Instructions|10378,10388|false|false|false|||irritation
Finding|Intellectual Product|Discharge Instructions|10378,10388|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Finding|Mental Process|Discharge Instructions|10378,10388|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Finding|Pathologic Function|Discharge Instructions|10378,10388|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Phenomenon|Phenomenon or Process|Discharge Instructions|10378,10388|false|false|false|C0441723|Irritation|irritation
Finding|Functional Concept|Discharge Instructions|10391,10395|false|false|false|C0947322;C1881534|Make - Instruction Imperative;Manufacturer Name|Make
Finding|Intellectual Product|Discharge Instructions|10391,10395|false|false|false|C0947322;C1881534|Make - Instruction Imperative;Manufacturer Name|Make
Event|Event|Discharge Instructions|10396,10400|false|false|false|||sure
Finding|Intellectual Product|Discharge Instructions|10396,10400|false|false|false|C4724437|SURE Test|sure
Event|Event|Discharge Instructions|10404,10408|false|false|false|||take
Drug|Organic Chemical|Discharge Instructions|10414,10421|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Drug|Pharmacologic Substance|Discharge Instructions|10414,10421|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Drug|Pharmacologic Substance|Discharge Instructions|10422,10432|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Discharge Instructions|10422,10432|false|false|false|||medication
Finding|Intellectual Product|Discharge Instructions|10422,10432|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Discharge Instructions|10439,10444|false|false|false|||meals
Finding|Daily or Recreational Activity|Discharge Instructions|10439,10444|false|false|false|C1998602|Meal (occasion for eating)|meals
Disorder|Disease or Syndrome|Discharge Instructions|10451,10456|false|false|false|C2676739|Chromosome 2q32-Q33 Deletion Syndrome|glass
Drug|Hazardous or Poisonous Substance|Discharge Instructions|10451,10456|false|false|false|C0025611|methamphetamine|glass
Drug|Organic Chemical|Discharge Instructions|10451,10456|false|false|false|C0025611|methamphetamine|glass
Drug|Pharmacologic Substance|Discharge Instructions|10451,10456|false|false|false|C0025611|methamphetamine|glass
Event|Event|Discharge Instructions|10451,10456|false|false|false|||glass
Drug|Food|Discharge Instructions|10460,10464|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|milk
Drug|Immunologic Factor|Discharge Instructions|10460,10464|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|milk
Drug|Pharmacologic Substance|Discharge Instructions|10460,10464|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|milk
Drug|Substance|Discharge Instructions|10460,10464|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|milk
Event|Event|Discharge Instructions|10460,10464|false|false|false|||milk
Finding|Body Substance|Discharge Instructions|10460,10464|false|false|false|C0026131;C1546713|Milk (body substance);Milk Specimen Code|milk
Finding|Intellectual Product|Discharge Instructions|10460,10464|false|false|false|C0026131;C1546713|Milk (body substance);Milk Specimen Code|milk
Event|Event|Discharge Instructions|10467,10468|false|false|false|||
Attribute|Clinical Attribute|Discharge Instructions|10468,10477|false|false|false|C1382187|Clearance of substance|Clearance
Event|Event|Discharge Instructions|10468,10477|false|false|false|||Clearance
Phenomenon|Natural Phenomenon or Process|Discharge Instructions|10468,10477|false|false|false|C2825073|Clearance [PK]|Clearance
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10468,10477|false|false|false|C4554548|Clearance procedure|Clearance
Event|Event|Discharge Instructions|10481,10486|false|false|false|||drive
Event|Event|Discharge Instructions|10491,10497|false|false|false|||return
Event|Occupational Activity|Discharge Instructions|10501,10505|false|false|false|C0043227|Work|work
Event|Event|Discharge Instructions|10514,10523|false|false|false|||addressed
Event|Event|Discharge Instructions|10548,10554|false|false|false|||office
Finding|Idea or Concept|Discharge Instructions|10548,10554|false|false|false|C1549636|Address type - Office|office
Procedure|Health Care Activity|Discharge Instructions|10548,10560|false|false|false|C0028900|Office Visits|office visit
Event|Event|Discharge Instructions|10555,10560|false|false|false|||visit
Finding|Social Behavior|Discharge Instructions|10555,10560|false|false|false|C0545082|Visit|visit
Event|Event|Discharge Instructions|10563,10567|false|false|false|||Make
Finding|Functional Concept|Discharge Instructions|10563,10567|false|false|false|C0947322;C1881534|Make - Instruction Imperative;Manufacturer Name|Make
Finding|Intellectual Product|Discharge Instructions|10563,10567|false|false|false|C0947322;C1881534|Make - Instruction Imperative;Manufacturer Name|Make
Event|Event|Discharge Instructions|10568,10572|false|false|false|||sure
Finding|Intellectual Product|Discharge Instructions|10568,10572|false|false|false|C4724437|SURE Test|sure
Event|Event|Discharge Instructions|10576,10584|false|false|false|||continue
Finding|Idea or Concept|Discharge Instructions|10576,10584|false|false|false|C0549178|Continuous|continue
Event|Event|Discharge Instructions|10588,10591|false|false|false|||use
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10597,10617|false|false|false|C0454512|Incentive spirometry|incentive spirometer
Finding|Finding|Discharge Instructions|10625,10632|false|false|false|C4534363|At home|at home
Event|Event|Discharge Instructions|10628,10632|false|false|false|||home
Finding|Idea or Concept|Discharge Instructions|10628,10632|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Discharge Instructions|10628,10632|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Discharge Instructions|10628,10632|false|false|false|C1553498|home health encounter|home
Event|Event|Discharge Instructions|10634,10638|false|false|false|||CALL
Finding|Functional Concept|Discharge Instructions|10634,10638|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|CALL
Finding|Gene or Genome|Discharge Instructions|10634,10638|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|CALL
Finding|Intellectual Product|Discharge Instructions|10634,10638|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|CALL
Finding|Mental Process|Discharge Instructions|10634,10638|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|CALL
Attribute|Clinical Attribute|Discharge Instructions|10644,10651|false|false|false|C5444295||SURGEON
Event|Event|Discharge Instructions|10644,10651|false|false|false|||SURGEON
Event|Event|Discharge Instructions|10671,10681|true|false|false|||EXPERIENCE
Finding|Mental Process|Discharge Instructions|10671,10681|true|false|false|C0237607;C0596545|Experience;Experience (Practice)|EXPERIENCE
Event|Event|Discharge Instructions|10682,10685|false|false|false|||ANY
Finding|Finding|Discharge Instructions|10706,10709|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Finding|Idea or Concept|Discharge Instructions|10706,10709|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Finding|Finding|Discharge Instructions|10706,10715|false|false|false|C0746890|new onset|New onset
Event|Event|Discharge Instructions|10710,10715|false|false|false|||onset
Event|Event|Discharge Instructions|10719,10726|false|false|false|||tremors
Finding|Sign or Symptom|Discharge Instructions|10719,10726|false|false|false|C0040822|Tremor|tremors
Event|Event|Discharge Instructions|10730,10738|false|false|false|||seizures
Finding|Sign or Symptom|Discharge Instructions|10730,10738|false|false|false|C0036572|Seizures|seizures
Disorder|Mental or Behavioral Dysfunction|Discharge Instructions|10745,10754|true|false|false|C0009676|Confusion|confusion
Event|Event|Discharge Instructions|10745,10754|true|false|false|||confusion
Finding|Finding|Discharge Instructions|10745,10754|true|false|false|C0683369|Clouded consciousness|confusion
Event|Event|Discharge Instructions|10758,10764|true|false|false|||change
Finding|Functional Concept|Discharge Instructions|10758,10764|true|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10758,10764|true|false|false|C4319952|Change - procedure|change
Finding|Functional Concept|Discharge Instructions|10758,10767|true|false|false|C0392747|Changing|change in
Attribute|Clinical Attribute|Discharge Instructions|10758,10781|true|false|false|C5774124||change in mental status
Finding|Finding|Discharge Instructions|10758,10781|true|false|false|C0856054|Mental status changes|change in mental status
Finding|Mental Process|Discharge Instructions|10768,10774|true|false|false|C0229992|Psyche structure|mental
Attribute|Clinical Attribute|Discharge Instructions|10768,10781|true|false|false|C0488568;C0488569||mental status
Finding|Finding|Discharge Instructions|10768,10781|true|false|false|C0278060|Mental state|mental status
Attribute|Clinical Attribute|Discharge Instructions|10775,10781|true|false|false|C5889824||status
Event|Event|Discharge Instructions|10775,10781|true|false|false|||status
Finding|Idea or Concept|Discharge Instructions|10775,10781|true|false|false|C1546481|What subject filter - Status|status
Event|Event|Discharge Instructions|10789,10797|true|false|false|||numbness
Finding|Finding|Discharge Instructions|10789,10797|true|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|Discharge Instructions|10789,10797|true|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Disorder|Disease or Syndrome|Discharge Instructions|10799,10807|true|false|false|C0030554|Paresthesia|tingling
Event|Event|Discharge Instructions|10799,10807|true|false|false|||tingling
Finding|Sign or Symptom|Discharge Instructions|10799,10807|true|false|false|C2242996|Has tingling sensation|tingling
Event|Event|Discharge Instructions|10809,10817|true|false|false|||weakness
Finding|Sign or Symptom|Discharge Instructions|10809,10817|true|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|10826,10837|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Attribute|Clinical Attribute|Discharge Instructions|10840,10844|false|false|false|C2598155||Pain
Event|Event|Discharge Instructions|10840,10844|false|false|false|||Pain
Finding|Functional Concept|Discharge Instructions|10840,10844|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Discharge Instructions|10840,10844|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Event|Event|Discharge Instructions|10848,10856|true|false|false|||headache
Finding|Sign or Symptom|Discharge Instructions|10848,10856|true|false|false|C0018681|Headache|headache
Event|Event|Discharge Instructions|10877,10887|true|false|false|||increasing
Event|Event|Discharge Instructions|10897,10905|true|false|false|||relieved
Attribute|Clinical Attribute|Discharge Instructions|10909,10913|true|false|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|10909,10913|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|10909,10913|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Pharmacologic Substance|Discharge Instructions|10914,10924|true|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Discharge Instructions|10914,10924|true|false|false|||medication
Finding|Intellectual Product|Discharge Instructions|10914,10924|true|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Finding|Finding|Discharge Instructions|10927,10932|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Finding|Sign or Symptom|Discharge Instructions|10927,10932|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Event|Event|Discharge Instructions|10949,10954|false|false|false|||equal
Finding|Intellectual Product|Discharge Instructions|10949,10954|false|false|false|C1549782|Relational Operator - Equal|equal
Procedure|Health Care Activity|Discharge Instructions|10969,10977|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|10978,10990|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|10978,10990|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|10978,10990|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

