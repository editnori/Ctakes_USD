 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|25,29
No|30,32
:|32,33
_|36,37
_|37,38
_|38,39
<EOL>|39,40
<EOL>|41,42
Admission|42,51
Date|52,56
:|56,57
_|59,60
_|60,61
_|61,62
Discharge|76,85
Date|86,90
:|90,91
_|94,95
_|95,96
_|96,97
<EOL>|97,98
<EOL>|99,100
Date|100,104
of|105,107
Birth|108,113
:|113,114
_|116,117
_|117,118
_|118,119
Sex|132,135
:|135,136
F|139,140
<EOL>|140,141
<EOL>|142,143
Service|143,150
:|150,151
MEDICINE|152,160
<EOL>|160,161
<EOL>|162,163
IV|175,177
Dye|178,181
,|181,182
Iodine|183,189
Containing|190,200
Contrast|201,209
Media|210,215
/|216,217
Oxycodone|218,227
/|228,229
<EOL>|230,231
cilostazol|231,241
/|242,243
Varenicline|244,255
<EOL>|255,256
<EOL>|257,258
Attending|258,267
:|267,268
_|269,270
_|270,271
_|271,272
.|272,273
<EOL>|273,274
<EOL>|275,276
Anemia|293,299
,|299,300
Melena|301,307
,|307,308
SOB|309,312
<EOL>|312,313
<EOL>|314,315
Major|315,320
Surgical|321,329
or|330,332
Invasive|333,341
Procedure|342,351
:|351,352
<EOL>|352,353
Upper|353,358
endoscopy|359,368
_|369,370
_|370,371
_|371,372
<EOL>|372,373
<EOL>|373,374
<EOL>|375,376
_|404,405
_|405,406
_|406,407
yo|408,410
female|411,417
with|418,422
history|423,430
of|431,433
Afib|434,438
on|439,441
Xarelto|442,449
,|449,450
COPD|451,455
,|455,456
HTN|457,460
,|460,461
PAD|462,465
who|466,469
<EOL>|470,471
presents|471,479
for|480,483
abnormal|484,492
labs|493,497
.|497,498
She|499,502
noted|503,508
dark|509,513
,|513,514
tarry|515,520
,|520,521
stool|522,527
on|528,530
<EOL>|531,532
_|532,533
_|533,534
_|534,535
and|536,539
presented|540,549
to|550,552
PCP|553,556
_|557,558
_|558,559
_|559,560
_|561,562
_|562,563
_|563,564
,|564,565
where|566,571
H|572,573
/|573,574
H|574,575
was|576,579
noted|580,585
<EOL>|586,587
to|587,589
be|590,592
8.8|593,596
/|596,597
28.6|597,601
from|602,606
prior|607,612
11.|613,616
_|616,617
_|617,618
_|618,619
.6|619,621
(|622,623
baseline|623,631
Hct|632,635
about|636,641
38|642,644
)|644,645
.|645,646
She|647,650
<EOL>|651,652
has|652,655
also|656,660
been|661,665
experiencing|666,678
bright|679,685
red|686,689
blood|690,695
with|696,700
wiping|701,707
,|707,708
she|709,712
<EOL>|713,714
believes|714,722
from|723,727
her|728,731
hemorrhoids|732,743
.|743,744
PCP|745,748
called|749,755
pt|756,758
who|759,762
agreed|763,769
to|770,772
come|773,777
<EOL>|778,779
to|779,781
ED|782,784
.|784,785
She|786,789
had|790,793
colonoscopy|794,805
in|806,808
_|809,810
_|810,811
_|811,812
with|813,817
showed|818,824
a|825,826
benign|827,833
polyp|834,839
,|839,840
<EOL>|841,842
internal|842,850
hemorrhoids|851,862
,|862,863
and|864,867
diverticulosis|868,882
.|882,883
Her|884,887
last|888,892
BM|893,895
was|896,899
_|900,901
_|901,902
_|902,903
,|903,904
<EOL>|905,906
was|906,909
reportedly|910,920
"|921,922
regular|922,929
.|929,930
"|930,931
She|932,935
currently|936,945
complains|946,955
of|956,958
increased|959,968
<EOL>|969,970
exertional|970,980
fatigue|981,988
and|989,992
has|993,996
been|997,1001
feeling|1002,1009
more|1010,1014
SOB|1015,1018
than|1019,1023
her|1024,1027
<EOL>|1028,1029
baseline|1029,1037
.|1037,1038
Over|1040,1044
the|1045,1048
last|1049,1053
6|1054,1055
months|1056,1062
she|1063,1066
has|1067,1070
noticed|1071,1078
she|1079,1082
becomes|1083,1090
<EOL>|1091,1092
increasingly|1092,1104
out|1105,1108
of|1109,1111
breath|1112,1118
,|1118,1119
walking|1120,1127
or|1128,1130
climbing|1131,1139
stairs|1140,1146
.|1146,1147
She|1149,1152
<EOL>|1153,1154
becomes|1154,1161
SOB|1162,1165
after|1166,1171
6|1172,1173
stairs|1174,1180
or|1181,1183
less|1184,1188
than|1189,1193
1|1194,1195
block|1196,1201
,|1201,1202
requiring|1203,1212
her|1213,1216
<EOL>|1217,1218
to|1218,1220
stop|1221,1225
,|1225,1226
and|1227,1230
at|1231,1233
times|1234,1239
use|1240,1243
albuterol|1244,1253
inhaler|1254,1261
.|1261,1262
She|1263,1266
used|1267,1271
to|1272,1274
use|1275,1278
her|1279,1282
<EOL>|1283,1284
only|1284,1288
use|1289,1292
her|1293,1296
inhaler|1297,1304
_|1305,1306
_|1306,1307
_|1307,1308
times|1309,1314
per|1315,1318
day|1319,1322
,|1322,1323
now|1324,1327
she|1328,1331
uses|1332,1336
it|1337,1339
over|1340,1344
<EOL>|1345,1346
four|1346,1350
times|1351,1356
a|1357,1358
day|1359,1362
and|1363,1366
nebulizers|1367,1377
twice|1378,1383
a|1384,1385
day|1386,1389
.|1389,1390
<EOL>|1391,1392
<EOL>|1392,1393
She|1393,1396
denies|1397,1403
any|1404,1407
fevers|1408,1414
,|1414,1415
chills|1416,1422
,|1422,1423
nausea|1424,1430
/|1430,1431
vomit|1431,1436
,|1436,1437
diarrhea|1438,1446
,|1446,1447
dysuria|1448,1455
,|1455,1456
<EOL>|1457,1458
rash|1458,1462
,|1462,1463
unintentional|1464,1477
weight|1478,1484
loss|1485,1489
.|1489,1490
<EOL>|1492,1493
<EOL>|1494,1495
<EOL>|1496,1497
In|1497,1499
the|1500,1503
ED|1504,1506
,|1506,1507
initial|1508,1515
vitals|1516,1522
:|1522,1523
0|1524,1525
98|1526,1528
64|1529,1531
149|1532,1535
/|1535,1536
85|1536,1538
20|1539,1541
98|1542,1544
%|1544,1545
RA|1546,1548
<EOL>|1549,1550
Labs|1550,1554
significant|1555,1566
for|1567,1570
:|1570,1571
<EOL>|1571,1572
WBC|1572,1575
5.0|1576,1579
HGB|1580,1583
8.8|1584,1587
HCT|1588,1591
28|1592,1594
.|1594,1595
4|1595,1596
(|1596,1597
Last|1598,1602
baseline|1603,1611
of|1612,1614
11.|1615,1618
_|1618,1619
_|1619,1620
_|1620,1621
/|1621,1622
34.6|1622,1626
in|1627,1629
<EOL>|1630,1631
_|1631,1632
_|1632,1633
_|1633,1634
MCV|1635,1638
PLT|1639,1642
240|1643,1646
<EOL>|1647,1648
_|1648,1649
_|1649,1650
_|1650,1651
16.7|1652,1656
INR|1657,1660
1.5|1661,1664
PTT|1665,1668
38.8|1669,1673
<EOL>|1673,1674
Chem|1674,1678
7|1679,1680
was|1681,1684
normal|1685,1691
<EOL>|1691,1692
<EOL>|1692,1693
She|1693,1696
was|1697,1700
given|1701,1706
albuterol|1707,1716
nebs|1717,1721
and|1722,1725
started|1726,1733
on|1734,1736
IV|1737,1739
normal|1740,1746
saline|1747,1753
<EOL>|1753,1754
<EOL>|1755,1756
On|1756,1758
transfer|1759,1767
,|1767,1768
vitals|1769,1775
were|1776,1780
:|1780,1781
T|1783,1784
:|1784,1785
98.4|1785,1789
BP|1791,1793
:|1793,1794
152|1795,1798
/|1798,1799
60|1799,1801
P|1802,1803
:|1803,1804
68|1804,1806
R|1807,1808
:|1808,1809
18|1809,1811
18|1812,1814
<EOL>|1815,1816
O2|1816,1818
:|1818,1819
97|1819,1821
%|1821,1822
RA|1822,1824
<EOL>|1826,1827
On|1827,1829
arrival|1830,1837
to|1838,1840
the|1841,1844
floor|1845,1850
patient|1851,1858
was|1859,1862
stable|1863,1869
and|1870,1873
in|1874,1876
good|1877,1881
spirits|1882,1889
.|1889,1890
<EOL>|1891,1892
She|1892,1895
notes|1896,1901
that|1902,1906
she|1907,1910
had|1911,1914
some|1915,1919
blood|1920,1925
per|1926,1929
rectum|1930,1936
on|1937,1939
her|1940,1943
underwear|1944,1953
.|1953,1954
<EOL>|1956,1957
<EOL>|1957,1958
<EOL>|1959,1960
ASTHMA|1982,1988
/|1988,1989
COPD|1989,1993
/|1993,1994
Tobacco|1994,2001
use|2002,2005
,|2005,2006
Peripheral|2007,2017
Arterial|2018,2026
disease|2027,2034
s|2035,2036
/|2036,2037
p|2037,2038
recent|2039,2045
<EOL>|2046,2047
common|2047,2053
iliac|2054,2059
stenting|2060,2068
,|2068,2069
ATRIAL|2070,2076
TACHYCARDIA|2077,2088
,|2088,2089
ATYPICAL|2090,2098
CHEST|2099,2104
PAIN|2105,2109
,|2109,2110
<EOL>|2111,2112
CERVICAL|2112,2120
RADICULITIS|2121,2132
,|2132,2133
CERVICAL|2134,2142
SPONDYLOSIS|2143,2154
,|2154,2155
CORONARY|2156,2164
ARTERY|2165,2171
<EOL>|2172,2173
DISEASE|2173,2180
<EOL>|2182,2183
HEADACHE|2183,2191
,|2191,2192
HIP|2193,2196
REPLACEMENT|2197,2208
,|2208,2209
HYPERLIPIDEMIA|2210,2224
,|2224,2225
HYPERTENSION|2226,2238
,|2238,2239
<EOL>|2240,2241
OSTEOARTHRITIS|2241,2255
,|2255,2256
HERPES|2257,2263
ZOSTER|2264,2270
,|2270,2271
TOBACCO|2272,2279
ABUSE|2280,2285
,|2285,2286
ATRIAL|2287,2293
<EOL>|2294,2295
FIBRILLATION|2295,2307
<EOL>|2309,2310
ANXIETY|2310,2317
,|2317,2318
GASTROINTESTINAL|2318,2334
BLEEDING|2335,2343
,|2343,2344
OSTEOARTHRITIS|2345,2359
,|2359,2360
<EOL>|2361,2362
ATHEROSCLEROTIC|2362,2377
CARDIOVASCULAR|2378,2392
DISEASE|2393,2400
,|2400,2401
PERIPHERAL|2402,2412
VASCULAR|2413,2421
<EOL>|2422,2423
DISEASE|2423,2430
,|2430,2431
CATARACT|2432,2440
SURGERY|2441,2448
_|2449,2450
_|2450,2451
_|2451,2452
<EOL>|2454,2455
Surgery|2455,2462
:|2462,2463
<EOL>|2465,2466
BILATERAL|2466,2475
COMMON|2476,2482
ILIAC|2483,2488
ARTERY|2489,2495
STENTING|2496,2504
_|2505,2506
_|2506,2507
_|2507,2508
<EOL>|2510,2511
BUNIONECTOMY|2511,2523
<EOL>|2525,2526
HIP|2526,2529
REPLACEMENT|2530,2541
<EOL>|2543,2544
PRIOR|2544,2549
CESAREAN|2550,2558
SECTION|2559,2566
<EOL>|2568,2569
GANGLION|2569,2577
CYST|2578,2582
<EOL>|2582,2583
<EOL>|2584,2585
:|2599,2600
<EOL>|2600,2601
_|2601,2602
_|2602,2603
_|2603,2604
<EOL>|2604,2605
:|2619,2620
<EOL>|2620,2621
Mother|2621,2627
:|2627,2628
_|2629,2630
_|2630,2631
_|2631,2632
,|2632,2633
HTN|2634,2637
<EOL>|2639,2640
Father|2640,2646
:|2646,2647
_|2648,2649
_|2649,2650
_|2650,2651
CA|2652,2654
<EOL>|2656,2657
Brother|2657,2664
:|2664,2665
CA|2666,2668
?|2668,2669
<EOL>|2671,2672
Brother|2672,2679
:|2679,2680
_|2681,2682
_|2682,2683
_|2683,2684
<EOL>|2685,2686
<EOL>|2687,2688
Physical|2688,2696
_|2697,2698
_|2698,2699
_|2699,2700
:|2700,2701
<EOL>|2701,2702
ADMISSION|2702,2711
PHYSICAL|2712,2720
EXAM|2721,2725
:|2725,2726
<EOL>|2726,2727
Vitals|2727,2733
:|2733,2734
T|2735,2736
:|2736,2737
98.4|2737,2741
BP|2743,2745
:|2745,2746
152|2747,2750
/|2750,2751
60|2751,2753
P|2754,2755
:|2755,2756
68|2756,2758
R|2759,2760
:|2760,2761
18|2761,2763
18|2764,2766
O2|2767,2769
:|2769,2770
97|2770,2772
%|2772,2773
RA|2773,2775
<EOL>|2777,2778
GENERAL|2778,2785
:|2785,2786
Well|2787,2791
nourished|2792,2801
,|2801,2802
well|2803,2807
appearing|2808,2817
AA|2818,2820
female|2821,2827
,|2827,2828
sitting|2829,2836
up|2837,2839
in|2840,2842
<EOL>|2843,2844
bed|2844,2847
Alert|2848,2853
,|2853,2854
oriented|2855,2863
,|2863,2864
no|2865,2867
acute|2868,2873
distress|2874,2882
<EOL>|2884,2885
HEENT|2885,2890
:|2890,2891
Sclera|2892,2898
anicteric|2899,2908
,|2908,2909
MMM|2910,2913
,|2913,2914
oropharynx|2915,2925
clear|2926,2931
<EOL>|2933,2934
NECK|2934,2938
:|2938,2939
supple|2940,2946
,|2946,2947
JVP|2948,2951
not|2952,2955
elevated|2956,2964
,|2964,2965
no|2966,2968
LAD|2969,2972
<EOL>|2974,2975
LUNGS|2975,2980
:|2980,2981
Clear|2982,2987
to|2988,2990
auscultation|2991,3003
bilaterally|3004,3015
though|3016,3022
decreased|3023,3032
air|3033,3036
<EOL>|3037,3038
movement|3038,3046
.|3046,3047
No|3048,3050
no|3051,3053
wheezes|3054,3061
,|3061,3062
rales|3063,3068
,|3068,3069
rhonchi|3070,3077
<EOL>|3079,3080
CV|3080,3082
:|3082,3083
Irregularly|3084,3095
irregular|3096,3105
rate|3106,3110
and|3111,3114
rhythm|3115,3121
,|3121,3122
normal|3123,3129
S1|3130,3132
S2|3133,3135
,|3135,3136
_|3137,3138
_|3138,3139
_|3139,3140
<EOL>|3141,3142
systolic|3142,3150
murmur|3151,3157
heard|3158,3163
best|3164,3168
at|3169,3171
RUSB|3172,3176
,|3176,3177
no|3178,3180
rubs|3181,3185
or|3186,3188
gallops|3189,3196
<EOL>|3198,3199
ABD|3199,3202
:|3202,3203
soft|3204,3208
,|3208,3209
non-tender|3210,3220
,|3220,3221
non-distended|3222,3235
,|3235,3236
bowel|3237,3242
sounds|3243,3249
present|3250,3257
,|3257,3258
no|3259,3261
<EOL>|3262,3263
rebound|3263,3270
tenderness|3271,3281
or|3282,3284
guarding|3285,3293
,|3293,3294
no|3295,3297
organomegaly|3298,3310
<EOL>|3311,3312
Rectum|3312,3318
:|3318,3319
No|3320,3322
obvious|3323,3330
hemorrhoids|3331,3342
<EOL>|3344,3345
EXT|3345,3348
:|3348,3349
Warm|3350,3354
,|3354,3355
well|3356,3360
perfused|3361,3369
,|3369,3370
2|3371,3372
+|3372,3373
pulses|3374,3380
,|3380,3381
no|3382,3384
clubbing|3385,3393
,|3393,3394
cyanosis|3395,3403
or|3404,3406
<EOL>|3407,3408
edema|3408,3413
<EOL>|3415,3416
SKIN|3416,3420
:|3420,3421
clear|3422,3427
<EOL>|3427,3428
NEURO|3428,3433
:|3433,3434
No|3435,3437
gross|3438,3443
deficits|3444,3452
.|3452,3453
<EOL>|3453,3454
<EOL>|3454,3455
DISCHARGE|3455,3464
PHYSICAL|3465,3473
EXAM|3474,3478
:|3478,3479
<EOL>|3479,3480
Vitals|3480,3486
:|3486,3487
T|3488,3489
:|3489,3490
98.2|3491,3495
,|3495,3496
BP|3497,3499
:|3499,3500
146|3501,3504
-|3504,3505
152|3505,3508
/|3508,3509
67|3509,3511
-|3511,3512
78|3512,3514
,|3514,3515
P|3516,3517
:|3517,3518
57|3518,3520
-|3520,3521
60|3521,3523
,|3523,3524
_|3525,3526
_|3526,3527
_|3527,3528
,|3528,3529
O2|3530,3532
:|3532,3533
97|3533,3535
%|3535,3536
RA|3536,3538
<EOL>|3540,3541
GENERAL|3541,3548
:|3548,3549
Well|3550,3554
nourished|3555,3564
,|3564,3565
well|3566,3570
appearing|3571,3580
,|3580,3581
sitting|3582,3589
up|3590,3592
in|3593,3595
bed|3596,3599
,|3599,3600
NAD|3601,3604
<EOL>|3604,3605
HEENT|3605,3610
:|3610,3611
Sclera|3612,3618
anicteric|3619,3628
,|3628,3629
MMM|3630,3633
,|3633,3634
oropharynx|3635,3645
clear|3646,3651
<EOL>|3653,3654
NECK|3654,3658
:|3658,3659
supple|3660,3666
,|3666,3667
JVP|3668,3671
not|3672,3675
elevated|3676,3684
,|3684,3685
no|3686,3688
LAD|3689,3692
<EOL>|3694,3695
LUNGS|3695,3700
:|3700,3701
Scattered|3702,3711
wheezes|3712,3719
bilaterally|3720,3731
but|3732,3735
no|3736,3738
resp|3739,3743
distress|3744,3752
<EOL>|3753,3754
CV|3754,3756
:|3756,3757
Irregularly|3758,3769
irregular|3770,3779
rate|3780,3784
and|3785,3788
rhythm|3789,3795
,|3795,3796
normal|3797,3803
S1|3804,3806
S2|3807,3809
,|3809,3810
_|3811,3812
_|3812,3813
_|3813,3814
<EOL>|3815,3816
systolic|3816,3824
murmur|3825,3831
heard|3832,3837
best|3838,3842
at|3843,3845
RUSB|3846,3850
,|3850,3851
no|3852,3854
rubs|3855,3859
or|3860,3862
gallops|3863,3870
<EOL>|3870,3871
ABD|3871,3874
:|3874,3875
soft|3876,3880
,|3880,3881
non-tender|3882,3892
,|3892,3893
non-distended|3894,3907
,|3907,3908
bowel|3909,3914
sounds|3915,3921
present|3922,3929
,|3929,3930
no|3931,3933
<EOL>|3934,3935
rebound|3935,3942
tenderness|3943,3953
or|3954,3956
guarding|3957,3965
,|3965,3966
no|3967,3969
organomegaly|3970,3982
<EOL>|3982,3983
EXT|3983,3986
:|3986,3987
Warm|3988,3992
,|3992,3993
well|3994,3998
perfused|3999,4007
,|4007,4008
2|4009,4010
+|4010,4011
pulses|4012,4018
,|4018,4019
no|4020,4022
clubbing|4023,4031
,|4031,4032
cyanosis|4033,4041
or|4042,4044
<EOL>|4045,4046
edema|4046,4051
<EOL>|4053,4054
SKIN|4054,4058
:|4058,4059
clear|4060,4065
<EOL>|4065,4066
NEURO|4066,4071
:|4071,4072
No|4073,4075
gross|4076,4081
deficits|4082,4090
.|4090,4091
<EOL>|4092,4093
<EOL>|4094,4095
Pertinent|4095,4104
Results|4105,4112
:|4112,4113
<EOL>|4113,4114
ADMISSION|4114,4123
LABS|4124,4128
:|4128,4129
<EOL>|4129,4130
=|4130,4131
=|4131,4132
=|4132,4133
=|4133,4134
=|4134,4135
=|4135,4136
=|4136,4137
=|4137,4138
=|4138,4139
=|4139,4140
=|4140,4141
=|4141,4142
=|4142,4143
=|4143,4144
=|4144,4145
=|4145,4146
<EOL>|4146,4147
_|4147,4148
_|4148,4149
_|4149,4150
12|4151,4153
:|4153,4154
28PM|4154,4158
BLOOD|4159,4164
WBC|4165,4168
-|4168,4169
5.0|4169,4172
RBC|4173,4176
-|4176,4177
3|4177,4178
.|4178,4179
28|4179,4181
*|4181,4182
Hgb|4183,4186
-|4186,4187
8|4187,4188
.|4188,4189
8|4189,4190
*|4190,4191
Hct|4192,4195
-|4195,4196
28|4196,4198
.|4198,4199
4|4199,4200
*|4200,4201
<EOL>|4202,4203
MCV|4203,4206
-|4206,4207
87|4207,4209
MCH|4210,4213
-|4213,4214
26.8|4214,4218
MCHC|4219,4223
-|4223,4224
31|4224,4226
.|4226,4227
0|4227,4228
*|4228,4229
RDW|4230,4233
-|4233,4234
16|4234,4236
.|4236,4237
1|4237,4238
*|4238,4239
RDWSD|4240,4245
-|4245,4246
50|4246,4248
.|4248,4249
4|4249,4250
*|4250,4251
Plt|4252,4255
_|4256,4257
_|4257,4258
_|4258,4259
<EOL>|4259,4260
_|4260,4261
_|4261,4262
_|4262,4263
02|4264,4266
:|4266,4267
28PM|4267,4271
BLOOD|4272,4277
_|4278,4279
_|4279,4280
_|4280,4281
PTT|4282,4285
-|4285,4286
38|4286,4288
.|4288,4289
8|4289,4290
*|4290,4291
_|4292,4293
_|4293,4294
_|4294,4295
<EOL>|4295,4296
_|4296,4297
_|4297,4298
_|4298,4299
12|4300,4302
:|4302,4303
28PM|4303,4307
BLOOD|4308,4313
Glucose|4314,4321
-|4321,4322
96|4322,4324
UreaN|4325,4330
-|4330,4331
18|4331,4333
Creat|4334,4339
-|4339,4340
1.0|4340,4343
Na|4344,4346
-|4346,4347
137|4347,4350
<EOL>|4351,4352
K|4352,4353
-|4353,4354
3.6|4354,4357
Cl|4358,4360
-|4360,4361
98|4361,4363
HCO3|4364,4368
-|4368,4369
28|4369,4371
AnGap|4372,4377
-|4377,4378
15|4378,4380
<EOL>|4380,4381
<EOL>|4381,4382
PERTINENT|4382,4391
FINDINGS|4392,4400
:|4400,4401
<EOL>|4401,4402
=|4402,4403
=|4403,4404
=|4404,4405
=|4405,4406
=|4406,4407
=|4407,4408
=|4408,4409
=|4409,4410
=|4410,4411
=|4411,4412
=|4412,4413
=|4413,4414
=|4414,4415
=|4415,4416
=|4416,4417
=|4417,4418
=|4418,4419
=|4419,4420
=|4420,4421
=|4421,4422
<EOL>|4422,4423
EGD|4423,4426
negative|4427,4435
for|4436,4439
evidence|4440,4448
of|4449,4451
bleeding|4452,4460
<EOL>|4460,4461
<EOL>|4461,4462
DISCHARGE|4462,4471
LABS|4472,4476
:|4476,4477
<EOL>|4477,4478
=|4478,4479
=|4479,4480
=|4480,4481
=|4481,4482
=|4482,4483
=|4483,4484
=|4484,4485
=|4485,4486
=|4486,4487
=|4487,4488
=|4488,4489
=|4489,4490
=|4490,4491
=|4491,4492
=|4492,4493
=|4493,4494
<EOL>|4494,4495
_|4495,4496
_|4496,4497
_|4497,4498
06|4499,4501
:|4501,4502
35AM|4502,4506
BLOOD|4507,4512
WBC|4513,4516
-|4516,4517
4.7|4517,4520
RBC|4521,4524
-|4524,4525
3|4525,4526
.|4526,4527
38|4527,4529
*|4529,4530
Hgb|4531,4534
-|4534,4535
9|4535,4536
.|4536,4537
1|4537,4538
*|4538,4539
Hct|4540,4543
-|4543,4544
29|4544,4546
.|4546,4547
1|4547,4548
*|4548,4549
<EOL>|4550,4551
MCV|4551,4554
-|4554,4555
86|4555,4557
MCH|4558,4561
-|4561,4562
26.9|4562,4566
MCHC|4567,4571
-|4571,4572
31|4572,4574
.|4574,4575
3|4575,4576
*|4576,4577
RDW|4578,4581
-|4581,4582
16|4582,4584
.|4584,4585
1|4585,4586
*|4586,4587
RDWSD|4588,4593
-|4593,4594
50|4594,4596
.|4596,4597
5|4597,4598
*|4598,4599
Plt|4600,4603
_|4604,4605
_|4605,4606
_|4606,4607
<EOL>|4607,4608
_|4608,4609
_|4609,4610
_|4610,4611
06|4612,4614
:|4614,4615
35AM|4615,4619
BLOOD|4620,4625
_|4626,4627
_|4627,4628
_|4628,4629
PTT|4630,4633
-|4633,4634
37|4634,4636
.|4636,4637
1|4637,4638
*|4638,4639
_|4640,4641
_|4641,4642
_|4642,4643
<EOL>|4643,4644
_|4644,4645
_|4645,4646
_|4646,4647
06|4648,4650
:|4650,4651
35AM|4651,4655
BLOOD|4656,4661
Glucose|4662,4669
-|4669,4670
99|4670,4672
UreaN|4673,4678
-|4678,4679
8|4679,4680
Creat|4681,4686
-|4686,4687
0.9|4687,4690
Na|4691,4693
-|4693,4694
137|4694,4697
<EOL>|4698,4699
K|4699,4700
-|4700,4701
3|4701,4702
.|4702,4703
2|4703,4704
*|4704,4705
Cl|4706,4708
-|4708,4709
98|4709,4711
HCO3|4712,4716
-|4716,4717
30|4717,4719
AnGap|4720,4725
-|4725,4726
12|4726,4728
<EOL>|4728,4729
_|4729,4730
_|4730,4731
_|4731,4732
06|4733,4735
:|4735,4736
35AM|4736,4740
BLOOD|4741,4746
Calcium|4747,4754
-|4754,4755
9.5|4755,4758
Phos|4759,4763
-|4763,4764
3.3|4764,4767
Mg|4768,4770
-|4770,4771
2|4771,4772
.|4772,4773
_|4773,4774
_|4774,4775
_|4775,4776
PMH|4777,4780
of|4781,4783
CAD|4784,4787
,|4787,4788
PVD|4789,4792
,|4792,4793
and|4794,4797
COPD|4798,4802
and|4803,4806
history|4807,4814
of|4815,4817
recurrent|4818,4827
chest|4828,4833
<EOL>|4834,4835
pain|4835,4839
present|4840,4847
with|4848,4852
drop|4853,4857
in|4858,4860
HCT|4861,4864
and|4865,4868
progressive|4869,4880
SOB|4881,4884
.|4884,4885
<EOL>|4886,4887
<EOL>|4887,4888
ACTIVE|4888,4894
PROBLEMS|4895,4903
<EOL>|4903,4904
#|4904,4905
GI|4905,4907
Bleed|4908,4913
:|4913,4914
Presented|4915,4924
to|4925,4927
PCP|4928,4931
with|4932,4936
melena|4937,4943
and|4944,4947
wiping|4948,4954
BRBPR|4955,4960
.|4960,4961
CBC|4962,4965
<EOL>|4966,4967
was|4967,4970
taken|4971,4976
and|4977,4980
Hgb|4981,4984
found|4985,4990
to|4991,4993
drop|4994,4998
from|4999,5003
11.3|5004,5008
-|5008,5009
>|5009,5010
8.8|5010,5013
.|5013,5014
Two|5015,5018
large|5019,5024
bore|5025,5029
<EOL>|5030,5031
IVs|5031,5034
were|5035,5039
placed|5040,5046
,|5046,5047
started|5048,5055
on|5056,5058
IV|5059,5061
PPI|5062,5065
,|5065,5066
and|5067,5070
she|5071,5074
was|5075,5078
type|5079,5083
and|5084,5087
<EOL>|5088,5089
screened|5089,5097
.|5097,5098
Vitals|5099,5105
remained|5106,5114
stable|5115,5121
,|5121,5122
so|5123,5125
patient|5126,5133
was|5134,5137
continued|5138,5147
on|5148,5150
<EOL>|5151,5152
home|5152,5156
rivaroxaban|5157,5168
.|5168,5169
She|5170,5173
was|5174,5177
evaluated|5178,5187
by|5188,5190
GI|5191,5193
who|5194,5197
recommended|5198,5209
upper|5210,5215
<EOL>|5216,5217
GI|5217,5219
endoscopy|5220,5229
,|5229,5230
which|5231,5236
showed|5237,5243
no|5244,5246
evidence|5247,5255
of|5256,5258
bleeding|5259,5267
.|5267,5268
She|5269,5272
remained|5273,5281
<EOL>|5282,5283
hemodynamically|5283,5298
stable|5299,5305
throughout|5306,5316
the|5317,5320
admission|5321,5330
.|5330,5331
Hgb|5332,5335
9.1|5336,5339
on|5340,5342
day|5343,5346
<EOL>|5347,5348
of|5348,5350
discharge|5351,5360
.|5360,5361
She|5362,5365
was|5366,5369
discharged|5370,5380
home|5381,5385
on|5386,5388
both|5389,5393
her|5394,5397
Xarelto|5398,5405
and|5406,5409
<EOL>|5410,5411
ASA|5411,5414
.|5414,5415
<EOL>|5415,5416
<EOL>|5416,5417
#|5417,5418
SOB|5418,5421
:|5421,5422
Long|5423,5427
standing|5428,5436
history|5437,5444
of|5445,5447
smoking|5448,5455
and|5456,5459
COPD|5460,5464
.|5464,5465
Progressive|5466,5477
<EOL>|5478,5479
exertional|5479,5489
dyspnea|5490,5497
despite|5498,5505
use|5506,5509
of|5510,5512
Spiriva|5513,5520
,|5520,5521
advair|5522,5528
,|5528,5529
fluticasone|5530,5541
<EOL>|5542,5543
nasal|5543,5548
spray|5549,5554
,|5554,5555
theophylline|5556,5568
,|5568,5569
and|5570,5573
albuterol|5574,5583
nebulizers|5584,5594
.|5594,5595
Has|5596,5599
<EOL>|5600,5601
increased|5601,5610
rescue|5611,5617
inhaler|5618,5625
use|5626,5629
.|5629,5630
Etiology|5632,5640
unclear|5641,5648
,|5648,5649
does|5650,5654
not|5655,5658
appear|5659,5665
<EOL>|5666,5667
to|5667,5669
be|5670,5672
infectious|5673,5683
given|5684,5689
chronicity|5690,5700
.|5700,5701
Most|5702,5706
likely|5707,5713
is|5714,5716
progression|5717,5728
of|5729,5731
<EOL>|5732,5733
underlying|5733,5743
COPD|5744,5748
.|5748,5749
PFT|5750,5753
's|5753,5755
were|5756,5760
obtained|5761,5769
while|5770,5775
in|5776,5778
-|5778,5779
house|5779,5784
.|5784,5785
Smoking|5786,5793
<EOL>|5794,5795
cessation|5795,5804
was|5805,5808
also|5809,5813
discussed|5814,5823
.|5823,5824
Will|5825,5829
need|5830,5834
continued|5835,5844
outpatient|5845,5855
f|5856,5857
/|5857,5858
u|5858,5859
<EOL>|5860,5861
re|5861,5863
:|5863,5864
her|5865,5868
COPD|5869,5873
.|5873,5874
<EOL>|5874,5875
<EOL>|5875,5876
CHRONIC|5876,5883
PROBLEMS|5884,5892
<EOL>|5892,5893
#|5893,5894
Afib|5894,5898
:|5898,5899
Continued|5900,5909
home|5910,5914
amiodarone|5915,5925
and|5926,5929
diltiazem|5930,5939
.|5939,5940
Continued|5941,5950
<EOL>|5951,5952
rivaroxaban|5952,5963
for|5964,5967
anticoagulation|5968,5983
,|5983,5984
as|5985,5987
discussed|5988,5997
above|5998,6003
.|6003,6004
<EOL>|6004,6005
<EOL>|6005,6006
#|6006,6007
HTN|6007,6010
:|6010,6011
Stable|6012,6018
,|6018,6019
continued|6020,6029
on|6030,6032
home|6033,6037
diltiazem|6038,6047
,|6047,6048
Imdur|6049,6054
,|6054,6055
HCTZ|6056,6060
<EOL>|6060,6061
<EOL>|6061,6062
#|6062,6063
Anxiety|6063,6070
/|6070,6071
insomnia|6071,6079
:|6079,6080
stable|6081,6087
,|6087,6088
continued|6089,6098
home|6099,6103
lorazepam|6104,6113
QHS|6114,6117
PRN|6118,6121
for|6122,6125
<EOL>|6126,6127
insomnia|6127,6135
/|6135,6136
anxiety|6136,6143
.|6143,6144
<EOL>|6144,6145
<EOL>|6145,6146
#|6146,6147
Dry|6147,6150
eyes|6151,6155
:|6155,6156
History|6157,6164
of|6165,6167
glaucoma|6168,6176
.|6176,6177
Continued|6178,6187
home|6188,6192
latanoprost|6193,6204
<EOL>|6205,6206
ophthalmic|6206,6216
drops|6217,6222
.|6222,6223
<EOL>|6223,6224
<EOL>|6224,6225
#|6225,6226
PAD|6226,6229
:|6229,6230
Stable|6231,6237
,|6237,6238
continued|6239,6248
on|6249,6251
home|6252,6256
atorvastatin|6257,6269
,|6269,6270
s|6271,6272
/|6272,6273
p|6273,6274
iliac|6275,6280
stent|6281,6286
.|6286,6287
<EOL>|6288,6289
OK|6289,6291
to|6292,6294
continue|6295,6303
aspirin|6304,6311
as|6312,6314
well|6315,6319
.|6319,6320
<EOL>|6320,6321
<EOL>|6321,6322
TRANSITIONAL|6322,6334
ISSUES|6335,6341
:|6341,6342
<EOL>|6342,6343
-|6343,6344
Should|6345,6351
consider|6352,6360
outpatient|6361,6371
colonoscopy|6372,6383
to|6384,6386
potentially|6387,6398
identify|6399,6407
<EOL>|6408,6409
any|6409,6412
source|6413,6419
of|6420,6422
lower|6423,6428
GI|6429,6431
Bleed|6432,6437
.|6437,6438
<EOL>|6438,6439
-|6439,6440
Given|6441,6446
stable|6447,6453
hemoglobin|6454,6464
/|6464,6465
hematocrit|6465,6475
while|6476,6481
inpatient|6482,6491
as|6492,6494
well|6495,6499
as|6500,6502
<EOL>|6503,6504
no|6504,6506
evidence|6507,6515
of|6516,6518
bleeding|6519,6527
on|6528,6530
EGD|6531,6534
,|6534,6535
her|6536,6539
Xarelto|6540,6547
and|6548,6551
Aspirin|6552,6559
were|6560,6564
<EOL>|6565,6566
continued|6566,6575
on|6576,6578
discharge|6579,6588
<EOL>|6588,6589
-|6589,6590
Was|6591,6594
treated|6595,6602
with|6603,6607
IV|6608,6610
PPI|6611,6614
while|6615,6620
inpatient|6621,6630
,|6630,6631
but|6632,6635
given|6636,6641
no|6642,6644
evidence|6645,6653
<EOL>|6654,6655
of|6655,6657
active|6658,6664
bleeding|6665,6673
,|6673,6674
was|6675,6678
discharged|6679,6689
on|6690,6692
home|6693,6697
Ranitidine|6698,6708
300mg|6709,6714
PO|6715,6717
<EOL>|6718,6719
daily|6719,6724
<EOL>|6724,6725
-|6725,6726
Continue|6727,6735
to|6736,6738
encourage|6739,6748
smoking|6749,6756
cessation|6757,6766
<EOL>|6766,6767
<EOL>|6767,6768
<EOL>|6769,6770
Medications|6770,6781
on|6782,6784
Admission|6785,6794
:|6794,6795
<EOL>|6795,6796
The|6796,6799
Preadmission|6800,6812
Medication|6813,6823
list|6824,6828
is|6829,6831
accurate|6832,6840
and|6841,6844
complete|6845,6853
.|6853,6854
<EOL>|6854,6855
1.|6855,6857
Rivaroxaban|6858,6869
20|6870,6872
mg|6873,6875
PO|6876,6878
QPM|6879,6882
<EOL>|6883,6884
2.|6884,6886
Acetaminophen|6887,6900
325|6901,6904
mg|6905,6907
PO|6908,6910
Q6H|6911,6914
:|6914,6915
PRN|6915,6918
pain|6919,6923
<EOL>|6924,6925
3.|6925,6927
Albuterol|6928,6937
0.083|6938,6943
%|6943,6944
Neb|6945,6948
Soln|6949,6953
1|6954,6955
NEB|6956,6959
IH|6960,6962
Q6H|6963,6966
:|6966,6967
PRN|6967,6970
SOB|6971,6974
<EOL>|6975,6976
4.|6976,6978
Aspirin|6979,6986
81|6987,6989
mg|6990,6992
PO|6993,6995
DAILY|6996,7001
<EOL>|7002,7003
5.|7003,7005
Atorvastatin|7006,7018
10|7019,7021
mg|7022,7024
PO|7025,7027
QPM|7028,7031
<EOL>|7032,7033
6.|7033,7035
Diltiazem|7036,7045
Extended|7046,7054
-|7054,7055
Release|7055,7062
180|7063,7066
mg|7067,7069
PO|7070,7072
BID|7073,7076
<EOL>|7077,7078
7.|7078,7080
Fluticasone|7081,7092
Propionate|7093,7103
NASAL|7104,7109
2|7110,7111
SPRY|7112,7116
NU|7117,7119
BID|7120,7123
nasal|7124,7129
congestion|7130,7140
<EOL>|7141,7142
8.|7142,7144
Fluticasone|7145,7156
-|7156,7157
Salmeterol|7157,7167
Diskus|7168,7174
(|7175,7176
250|7176,7179
/|7179,7180
50|7180,7182
)|7182,7183
1|7185,7186
INH|7187,7190
IH|7191,7193
BID|7194,7197
<EOL>|7198,7199
9.|7199,7201
Hydrochlorothiazide|7202,7221
50|7222,7224
mg|7225,7227
PO|7228,7230
DAILY|7231,7236
<EOL>|7237,7238
10.|7238,7241
Isosorbide|7242,7252
Mononitrate|7253,7264
(|7265,7266
Extended|7266,7274
Release|7275,7282
)|7282,7283
240|7284,7287
mg|7288,7290
PO|7291,7293
DAILY|7294,7299
<EOL>|7300,7301
11.|7301,7304
Latanoprost|7305,7316
0.005|7317,7322
%|7322,7323
Ophth|7324,7329
.|7329,7330
Soln.|7331,7336
1|7337,7338
DROP|7339,7343
LEFT|7344,7348
EYE|7349,7352
QHS|7353,7356
<EOL>|7357,7358
12.|7358,7361
Lorazepam|7362,7371
0.5|7372,7375
mg|7376,7378
PO|7379,7381
QHS|7382,7385
:|7385,7386
PRN|7386,7389
insomnia|7390,7398
<EOL>|7399,7400
13.|7400,7403
Multivitamins|7404,7417
W|7418,7419
/|7419,7420
minerals|7420,7428
1|7429,7430
TAB|7431,7434
PO|7435,7437
DAILY|7438,7443
<EOL>|7444,7445
14.|7445,7448
Ranitidine|7449,7459
300|7460,7463
mg|7464,7466
PO|7467,7469
DAILY|7470,7475
<EOL>|7476,7477
15.|7477,7480
Theophylline|7481,7493
ER|7494,7496
300|7497,7500
mg|7501,7503
PO|7504,7506
BID|7507,7510
<EOL>|7511,7512
16|7512,7514
.|7514,7515
Tiotropium|7516,7526
Bromide|7527,7534
1|7535,7536
CAP|7537,7540
IH|7541,7543
BID|7544,7547
<EOL>|7548,7549
17.|7549,7552
TraMADOL|7553,7561
(|7562,7563
Ultram|7563,7569
)|7569,7570
50|7571,7573
mg|7574,7576
PO|7577,7579
BID|7580,7583
pain|7584,7588
<EOL>|7589,7590
18.|7590,7593
Artificial|7594,7604
Tears|7605,7610
Preserv|7611,7618
.|7618,7619
Free|7620,7624
_|7625,7626
_|7626,7627
_|7627,7628
DROP|7629,7633
BOTH|7634,7638
EYES|7639,7643
PRN|7644,7647
<EOL>|7648,7649
irritation|7649,7659
<EOL>|7660,7661
19|7661,7663
.|7663,7664
Amiodarone|7665,7675
200|7676,7679
mg|7680,7682
PO|7683,7685
DAILY|7686,7691
<EOL>|7692,7693
<EOL>|7693,7694
<EOL>|7695,7696
Discharge|7696,7705
Medications|7706,7717
:|7717,7718
<EOL>|7718,7719
1.|7719,7721
Acetaminophen|7722,7735
325|7736,7739
mg|7740,7742
PO|7743,7745
Q6H|7746,7749
:|7749,7750
PRN|7750,7753
pain|7754,7758
<EOL>|7759,7760
2.|7760,7762
Albuterol|7763,7772
0.083|7773,7778
%|7778,7779
Neb|7780,7783
Soln|7784,7788
1|7789,7790
NEB|7791,7794
IH|7795,7797
Q6H|7798,7801
:|7801,7802
PRN|7802,7805
SOB|7806,7809
<EOL>|7810,7811
3.|7811,7813
Amiodarone|7814,7824
200|7825,7828
mg|7829,7831
PO|7832,7834
DAILY|7835,7840
<EOL>|7841,7842
4.|7842,7844
Atorvastatin|7845,7857
10|7858,7860
mg|7861,7863
PO|7864,7866
QPM|7867,7870
<EOL>|7871,7872
5.|7872,7874
Artificial|7875,7885
Tears|7886,7891
Preserv|7892,7899
.|7899,7900
Free|7901,7905
_|7906,7907
_|7907,7908
_|7908,7909
DROP|7910,7914
BOTH|7915,7919
EYES|7920,7924
PRN|7925,7928
<EOL>|7929,7930
irritation|7930,7940
<EOL>|7941,7942
6.|7942,7944
Diltiazem|7945,7954
Extended|7955,7963
-|7963,7964
Release|7964,7971
180|7972,7975
mg|7976,7978
PO|7979,7981
BID|7982,7985
<EOL>|7986,7987
7.|7987,7989
Fluticasone|7990,8001
Propionate|8002,8012
NASAL|8013,8018
2|8019,8020
SPRY|8021,8025
NU|8026,8028
BID|8029,8032
nasal|8033,8038
congestion|8039,8049
<EOL>|8050,8051
8.|8051,8053
Fluticasone|8054,8065
-|8065,8066
Salmeterol|8066,8076
Diskus|8077,8083
(|8084,8085
250|8085,8088
/|8088,8089
50|8089,8091
)|8091,8092
1|8094,8095
INH|8096,8099
IH|8100,8102
BID|8103,8106
<EOL>|8107,8108
9.|8108,8110
Hydrochlorothiazide|8111,8130
50|8131,8133
mg|8134,8136
PO|8137,8139
DAILY|8140,8145
<EOL>|8146,8147
10.|8147,8150
Isosorbide|8151,8161
Mononitrate|8162,8173
(|8174,8175
Extended|8175,8183
Release|8184,8191
)|8191,8192
240|8193,8196
mg|8197,8199
PO|8200,8202
DAILY|8203,8208
<EOL>|8209,8210
11.|8210,8213
Latanoprost|8214,8225
0.005|8226,8231
%|8231,8232
Ophth|8233,8238
.|8238,8239
Soln.|8240,8245
1|8246,8247
DROP|8248,8252
LEFT|8253,8257
EYE|8258,8261
QHS|8262,8265
<EOL>|8266,8267
12.|8267,8270
Lorazepam|8271,8280
0.5|8281,8284
mg|8285,8287
PO|8288,8290
QHS|8291,8294
:|8294,8295
PRN|8295,8298
insomnia|8299,8307
<EOL>|8308,8309
13.|8309,8312
Rivaroxaban|8313,8324
20|8325,8327
mg|8328,8330
PO|8331,8333
QPM|8334,8337
<EOL>|8338,8339
14.|8339,8342
Theophylline|8343,8355
ER|8356,8358
300|8359,8362
mg|8363,8365
PO|8366,8368
BID|8369,8372
<EOL>|8373,8374
15.|8374,8377
Ranitidine|8378,8388
300|8389,8392
mg|8393,8395
PO|8396,8398
DAILY|8399,8404
<EOL>|8405,8406
16|8406,8408
.|8408,8409
TraMADOL|8410,8418
(|8419,8420
Ultram|8420,8426
)|8426,8427
50|8428,8430
mg|8431,8433
PO|8434,8436
BID|8437,8440
pain|8441,8445
<EOL>|8446,8447
17|8447,8449
.|8449,8450
Tiotropium|8451,8461
Bromide|8462,8469
1|8470,8471
CAP|8472,8475
IH|8476,8478
BID|8479,8482
<EOL>|8483,8484
18.|8484,8487
Multivitamins|8488,8501
W|8502,8503
/|8503,8504
minerals|8504,8512
1|8513,8514
TAB|8515,8518
PO|8519,8521
DAILY|8522,8527
<EOL>|8528,8529
19|8529,8531
.|8531,8532
Aspirin|8533,8540
81|8541,8543
mg|8544,8546
PO|8547,8549
DAILY|8550,8555
<EOL>|8556,8557
<EOL>|8557,8558
<EOL>|8559,8560
Discharge|8560,8569
Disposition|8570,8581
:|8581,8582
<EOL>|8582,8583
Home|8583,8587
<EOL>|8587,8588
<EOL>|8589,8590
Discharge|8590,8599
Diagnosis|8600,8609
:|8609,8610
<EOL>|8610,8611
Primary|8611,8618
:|8618,8619
<EOL>|8619,8620
-|8620,8621
Anemia|8622,8628
<EOL>|8628,8629
<EOL>|8629,8630
Secondary|8630,8639
:|8639,8640
<EOL>|8640,8641
-|8641,8642
Afib|8643,8647
<EOL>|8647,8648
-|8648,8649
CAD|8650,8653
<EOL>|8653,8654
-|8654,8655
HTN|8656,8659
<EOL>|8659,8660
-|8660,8661
COPD|8662,8666
<EOL>|8666,8667
<EOL>|8667,8668
<EOL>|8669,8670
Mental|8691,8697
Status|8698,8704
:|8704,8705
Clear|8706,8711
and|8712,8715
coherent|8716,8724
.|8724,8725
<EOL>|8725,8726
Level|8726,8731
of|8732,8734
Consciousness|8735,8748
:|8748,8749
Alert|8750,8755
and|8756,8759
interactive|8760,8771
.|8771,8772
<EOL>|8772,8773
Activity|8773,8781
Status|8782,8788
:|8788,8789
Ambulatory|8790,8800
-|8801,8802
Independent|8803,8814
.|8814,8815
<EOL>|8815,8816
<EOL>|8816,8817
<EOL>|8818,8819
Ms.|8843,8846
_|8847,8848
_|8848,8849
_|8849,8850
,|8850,8851
<EOL>|8851,8852
<EOL>|8852,8853
You|8853,8856
were|8857,8861
admitted|8862,8870
to|8871,8873
_|8874,8875
_|8875,8876
_|8876,8877
due|8878,8881
to|8882,8884
<EOL>|8885,8886
a|8886,8887
decrease|8888,8896
in|8897,8899
blood|8900,8905
count|8906,8911
on|8912,8914
laboratory|8915,8925
testing|8926,8933
.|8933,8934
Because|8935,8942
we|8943,8945
were|8946,8950
<EOL>|8951,8952
concerned|8952,8961
for|8962,8965
a|8966,8967
bleed|8968,8973
in|8974,8976
your|8977,8981
GI|8982,8984
tract|8985,8990
,|8990,8991
you|8992,8995
underwent|8996,9005
an|9006,9008
upper|9009,9014
<EOL>|9015,9016
endoscopy|9016,9025
.|9025,9026
Fortunately|9027,9038
,|9038,9039
this|9040,9044
did|9045,9048
not|9049,9052
show|9053,9057
any|9058,9061
evidence|9062,9070
of|9071,9073
<EOL>|9074,9075
bleeding|9075,9083
.|9083,9084
Your|9085,9089
blood|9090,9095
counts|9096,9102
remained|9103,9111
stable|9112,9118
while|9119,9124
in|9125,9127
the|9128,9131
<EOL>|9132,9133
hospital|9133,9141
.|9141,9142
You|9143,9146
were|9147,9151
discharged|9152,9162
with|9163,9167
plan|9168,9172
for|9173,9176
outpatient|9177,9187
follow|9188,9194
up|9195,9197
<EOL>|9198,9199
with|9199,9203
GI|9204,9206
for|9207,9210
colonoscopy|9211,9222
in|9223,9225
the|9226,9229
future|9230,9236
.|9236,9237
Pulmonary|9238,9247
function|9248,9256
<EOL>|9257,9258
testing|9258,9265
was|9266,9269
done|9270,9274
as|9275,9277
well|9278,9282
while|9283,9288
you|9289,9292
were|9293,9297
here|9298,9302
.|9302,9303
You|9304,9307
will|9308,9312
also|9313,9317
<EOL>|9318,9319
follow|9319,9325
up|9326,9328
with|9329,9333
Dr.|9334,9337
_|9338,9339
_|9339,9340
_|9340,9341
in|9342,9344
his|9345,9348
clinic|9349,9355
.|9355,9356
<EOL>|9356,9357
<EOL>|9357,9358
It|9358,9360
was|9361,9364
a|9365,9366
pleasure|9367,9375
taking|9376,9382
care|9383,9387
of|9388,9390
your|9391,9395
at|9396,9398
_|9399,9400
_|9400,9401
_|9401,9402
.|9402,9403
If|9404,9406
you|9407,9410
have|9411,9415
any|9416,9419
<EOL>|9420,9421
questions|9421,9430
about|9431,9436
the|9437,9440
care|9441,9445
you|9446,9449
received|9450,9458
,|9458,9459
please|9460,9466
do|9467,9469
not|9470,9473
hesitate|9474,9482
to|9483,9485
<EOL>|9486,9487
ask|9487,9490
.|9490,9491
<EOL>|9491,9492
<EOL>|9492,9493
Sincerely|9493,9502
,|9502,9503
<EOL>|9503,9504
Your|9504,9508
Inpatient|9509,9518
_|9519,9520
_|9520,9521
_|9521,9522
Care|9523,9527
Team|9528,9532
<EOL>|9532,9533
<EOL>|9533,9534
<EOL>|9535,9536
Followup|9536,9544
Instructions|9545,9557
:|9557,9558
<EOL>|9558,9559
_|9559,9560
_|9560,9561
_|9561,9562
<EOL>|9562,9563

