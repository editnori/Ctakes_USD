CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Known|Modifier|false|false||Knownnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Adverse reaction to drug|Finding|true|false||Adverse Drug Reactionsnull|Adverse reaction to drug|Finding|true|false||Drug Reactionsnull|Pharmaceutical Preparations|Drug|false|false||Drug
null|Pharmacologic Substance|Drug|false|false||Drugnull|Drug problem|Finding|false|false||Drugnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Chief complaint (finding)|Finding|false|false||Chief Complaintnull|Complaint (finding)|Finding|false|false||Complaintnull|null|Attribute|false|false||Complaintnull|Deep thrombophlebitis|Disorder|false|false|C5239664|DVT
null|Deep Vein Thrombosis|Disorder|false|false|C5239664|DVTnull|area DVT|Anatomy|false|false|C0149871;C0151950;C2926618|DVTnull|null|Attribute|false|false|C5239664|DVTnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Esophagogastroduodenoscopy|Procedure|false|false||EGDnull|History of present illness (finding)|Finding|false|false||History of Present Illnessnull|null|Attribute|false|false||History of Present Illnessnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Present illness|Finding|false|false||Present Illnessnull|Present|Finding|false|false||Present
null|Presentation|Finding|false|false||Presentnull|Illness (finding)|Finding|false|false||Illnessnull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Hypertensive disease|Disorder|false|false||HTNnull|Chronic Kidney Diseases|Disorder|false|false||CKDnull|Stage level 4|Finding|false|false||stage IVnull|Tumor stage|Attribute|false|false||stagenull|Stage|Time|false|false||stage
null|Phase|Time|false|false||stagenull|Peripheral Vascular Diseases|Disorder|false|false||PVDnull|Pomalidomide/Bortezomib/Dexamethasone Regimen|Procedure|false|false||PVDnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Superficial|Modifier|false|false||superficialnull|Femur|Anatomy|false|false||femoralnull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Structure of left lower leg|Anatomy|false|false||lower Left legnull|Body Site Modifier - Lower|Anatomy|false|false|C2003888|lowernull|Lower (action)|Event|false|false|C1548802|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|numbness of left leg|Finding|false|false|C1140621;C0023216;C0230443;C0230416|Left leg numbnessnull|Structure of left lower leg|Anatomy|false|false|C2219779|Left leg
null|Left lower extremity|Anatomy|false|false|C2219779|Left legnull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Numbness in leg|Finding|false|false|C1140621;C0023216|leg numbnessnull|Lower Extremity|Anatomy|false|false|C0857160;C2219779|leg
null|Leg|Anatomy|false|false|C0857160;C2219779|legnull|Numbness|Finding|false|false||numbness
null|Hypesthesia|Finding|false|false||numbnessnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Evening|Time|false|false||eveningnull|Numbness|Finding|false|false||numbness
null|Hypesthesia|Finding|false|false||numbnessnull|Last|Modifier|false|false||lastnull|Night time|Time|false|false||nightnull|BORNHOLM EYE DISEASE|Disorder|false|false||bednull|Bachelor of Education|Finding|false|false||bednull|Beds|Device|false|false||bednull|Patient Location - Bed|Modifier|false|false||bednull|Onset of (contextual qualifier)|Modifier|false|false||onsetnull|Age of Onset|LabModifier|false|false||onsetnull|Gradual|Modifier|false|false||gradualnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Muscle Cramp|Finding|false|false||crampingnull|Cramping sensation quality|Modifier|false|false||crampingnull|Lateral|Modifier|false|false||lateralnull|Structure of calf of leg|Anatomy|false|false|C0555980|calf
null|null|Anatomy|false|false|C0555980|calfnull|Cattle calf (organism)|Entity|false|false||calfnull|Foot problem|Finding|false|false|C4299097;C0016504;C0230445;C1305418|footnull|Lower extremity>Foot|Anatomy|false|false|C0555980|foot
null|Foot|Anatomy|false|false|C0555980|footnull|Foot Unit of Length|LabModifier|false|false||footnull|Usually|Finding|false|false||usuallynull|Usual|Modifier|false|false||usuallynull|BORNHOLM EYE DISEASE|Disorder|false|false||bednull|Bachelor of Education|Finding|false|false||bednull|Beds|Device|false|false||bednull|Patient Location - Bed|Modifier|false|false||bednull|Exertion|Finding|false|false||exertionnull|Muscle Weakness Lower Limb|Finding|true|false|C1140621;C0023216|leg weakness
null|Monoparesis of lower limb|Finding|true|false|C1140621;C0023216|leg weaknessnull|Leg|Anatomy|false|false|C3714552;C0004093;C1836296;C0427068|leg
null|Lower Extremity|Anatomy|false|false|C3714552;C0004093;C1836296;C0427068|legnull|Weakness|Finding|true|false|C1140621;C0023216|weakness
null|Asthenia|Finding|true|false|C1140621;C0023216|weaknessnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|Helping Behavior|Finding|true|false||assistancenull|Assisted (qualifier value)|Modifier|false|false||assistancenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Numbness|Finding|false|false||numbness
null|Hypesthesia|Finding|false|false||numbnessnull|Residual|Modifier|false|false||residualnull|Numbness|Finding|false|false|C0230445;C1305418|numbness
null|Hypesthesia|Finding|false|false|C0230445;C1305418|numbnessnull|Lateral|Modifier|false|false||lateralnull|Structure of calf of leg|Anatomy|false|false|C0028643;C0020580|calf
null|null|Anatomy|false|false|C0028643;C0020580|calfnull|Cattle calf (organism)|Entity|false|false||calfnull|Deep thrombophlebitis|Disorder|true|false|C5239664|DVT
null|Deep Vein Thrombosis|Disorder|true|false|C5239664|DVTnull|area DVT|Anatomy|false|false|C0149871;C0151950;C2926618|DVTnull|null|Attribute|true|false|C5239664|DVTnull|Spine Problem|Finding|false|false|C2752558;C0037949|spinenull|Neuron spine|Anatomy|false|false|C0150920|spine
null|Vertebral column|Anatomy|false|false|C0150920|spinenull|Physical trauma|Disorder|true|false||trauma
null|Traumatic injury|Disorder|true|false||trauma
null|Trauma|Disorder|true|false||traumanull|Trauma assessment and care|Procedure|true|false||traumanull|Trauma, nursing specialty|Title|false|false||traumanull|trauma qualifier|Modifier|false|false||traumanull|Back Pain|Finding|true|false||back painnull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Incontinence|Disorder|true|false||incontinencenull|Fever|Finding|false|false||feversnull|Chills|Finding|false|false||chillsnull|Numbness|Finding|true|false||numbness
null|Hypesthesia|Finding|true|false||numbnessnull|Headache|Finding|false|false||headachenull|Visual changes|Finding|false|false||visual changesnull|Visual|Finding|false|false||visualnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0741025;C2926613;C0008031|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025;C2926613;C0008031|chestnull|Chest Pain|Finding|false|false|C1527391;C0817096|pain, chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Chest pressure|Finding|false|false|C1527391;C0817096|chest pressurenull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0438716;C0741025;C0008031|chest
null|Anterior thoracic region|Anatomy|false|false|C0438716;C0741025;C0008031|chestnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0741025|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025|chestnull|Palpitations|Finding|false|false||palpitationsnull|Dyspnea|Finding|false|false||shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false||breathnull|Abdominal Pain|Finding|false|false|C0000726|abdominal painnull|Abdomen|Anatomy|false|false|C0000737;C1549543;C0030193|abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Administration Method - Pain|Finding|false|false|C0000726|pain
null|Pain|Finding|false|false|C0000726|painnull|null|Attribute|false|false||painnull|Dysuria|Finding|false|false||dysurianull|rectal discharge diarrhea (physical finding)|Finding|false|false||diarrhea
null|Diarrhea|Finding|false|false||diarrheanull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Hypertensive disease|Disorder|false|false||hypertensionnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||diabetes
null|Diabetes|Disorder|false|false||diabetes
null|Diabetes Mellitus|Disorder|false|false||diabetesnull|Cyclophosphamide/Doxorubicin/Vincristine|Drug|false|false||CVAnull|Acute ill-defined cerebrovascular disease|Disorder|false|false||CVA
null|Cerebrovascular accident|Disorder|false|false||CVAnull|Cerebellum|Anatomy|false|false||cerebellarnull|Medullary - body parts|Anatomy|false|false|C0038454;C5977286|medullary
null|Medulla Oblongata|Anatomy|false|false|C0038454;C5977286|medullary
null|Adrenal Medulla|Anatomy|false|false|C0038454;C5977286|medullarynull|Cerebrovascular accident|Disorder|false|false|C1550278;C0025148;C0001629|strokenull|Stroke (heart beat)|Finding|false|false|C1550278;C0025148;C0001629|strokenull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Burning Mouth Syndrome|Disorder|false|false||BMSnull|Circumflex|Modifier|false|false||circumflexnull|Peripheral Arterial Diseases|Disorder|false|false|C0003842|peripheral arterial disease
null|Peripheral Vascular Diseases|Disorder|false|false|C0003842|peripheral arterial diseasenull|Peripheral|Modifier|false|false||peripheralnull|Arteriopathic disease|Disorder|false|false|C0003842|arterial diseasenull|Arteries|Anatomy|false|false|C0021775;C1704436;C0085096;C0012634;C1456822;C0311395;C0852949|arterialnull|Arterial|Modifier|false|false||arterialnull|Disease|Disorder|false|false|C0003842|diseasenull|Intermittent Claudication|Disorder|false|false|C0003842|claudicationnull|Claudication (finding)|Finding|false|false|C0003842|claudication
null|Lameness|Finding|false|false|C0003842|claudicationnull|Blood Vessel|Anatomy|false|false||vascularnull|Vascular|Modifier|false|false||vascularnull|Stage level 4|Finding|false|false||stage IVnull|Tumor stage|Attribute|false|false||stagenull|Stage|Time|false|false||stage
null|Phase|Time|false|false||stagenull|Chronic Kidney Diseases|Disorder|false|false||CKDnull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Gastroesophageal reflux disease|Disorder|false|false||GERDnull|Terminal esophageal web|Disorder|false|false||esophageal ringsnull|Esophageal Diseases|Disorder|false|false||esophagealnull|Esophageal|Modifier|false|false||esophagealnull|Ring device|Device|false|false||ringsnull|ring form of protozoa|Entity|false|false||ringsnull|Social and personal history|Finding|false|false||Social History
null|Social History|Finding|false|false||Social Historynull|Social|Finding|false|false||Socialnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Family Medical History|Finding|false|false||Family Historynull|Entity Name Part Type - family|Finding|false|false||Family
null|Last Name|Finding|false|false||Family
null|Living Arrangement - Family|Finding|false|false||Family
null|Family (taxonomic)|Finding|false|false||Family
null|Family Collection|Finding|false|false||Familynull|Family|Subject|false|false||Familynull|History of present illness (finding)|Finding|false|true||History
null|History of previous events|Finding|false|true||History
null|Historical aspects qualifier|Finding|false|true||History
null|Medical History|Finding|false|true||History
null|Concept History|Finding|false|true||Historynull|History|Subject|false|false||Historynull|Niece|Subject|false|false||Niecenull|Sorting - Cell Movement|Finding|false|false||sort
null|Sorting (Cognition)|Finding|false|false||sortnull|Sorting|Event|false|false||sortnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Indirect exposure mechanism - Father|Finding|false|false||Father
null|Relationship - Father|Finding|false|false||Father
null|Father - courtesy title|Finding|false|false||Fathernull|Father (person)|Subject|false|false||Fathernull|Lung diseases|Disorder|false|false|C4037972;C0024109|lung diseasenull|Lung diseases|Disorder|false|false|C4037972;C0024109|lungnull|Lung Problem|Finding|false|false|C4037972;C0024109|lungnull|Chest>Lung|Anatomy|false|false|C0012634;C0024115;C0740941;C0024115|lung
null|Lung|Anatomy|false|false|C0012634;C0024115;C0740941;C0024115|lungnull|Disease|Disorder|false|false|C4037972;C0024109|diseasenull|Relationship - Mother|Finding|false|false||Mothernull|Mother (person)|Subject|false|false||Mothernull|unknown vaccine or immune globulin|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|unknown vaccine or immune globulin|Drug|false|false||unknownnull|Unknown - Patient_s Relationship to Insured|Finding|false|false||unknown
null|Unknown - Special Program Code|Finding|false|false||unknown
null|Unknown - Production Class Code|Finding|false|false||unknown
null|Unknown - Patient Outcome|Finding|false|false||unknown
null|Unknown - Recreational Drug Use Code|Finding|false|false||unknown
null|Unknown - Escort Required|Finding|false|false||unknown
null|Unknown - Transport Arranged|Finding|false|false||unknown
null|Unknown - Living Arrangement|Finding|false|false||unknown
null|Unknown - Employment Status|Finding|false|false||unknown
null|Unknown - Relationship|Finding|false|false||unknown
null|Unknown - publishing section|Finding|false|false||unknown
null|Unknown Publicity Code|Finding|false|false||unknown
null|Unknown - Event reason|Finding|false|false||unknown
null|Unknown - Religion|Finding|false|false||unknown
null|Unknown - Organ Donor Code|Finding|false|false||unknown
null|unknown - NullFlavor|Finding|false|false||unknown
null|Unknown - Notify Clergy Code|Finding|false|false||unknown
null|Unknown - Administrative Gender|Finding|false|false||unknown
null|Unknown - Patient Condition Code|Finding|false|false||unknown
null|Unknown - Living Will Code|Finding|false|false||unknown
null|Marital Status - Unknown|Finding|false|false||unknown
null|Unknown - mode of arrival code|Finding|false|false||unknown
null|Unknown - Patient Class|Finding|false|false||unknown
null|Unknown - Event Expected|Finding|false|false||unknown
null|Unknown - Expanded yes/no indicator|Finding|false|false||unknown
null|Unknown - Immunization Registry Status|Finding|false|false||unknown
null|Unknown - Container status|Finding|false|false||unknown
null|Unknown - CWE statuses|Finding|false|false||unknown
null|Unknown - Job Status|Finding|false|false||unknown
null|Unknown - Precaution Code|Finding|false|false||unknown
null|Unknown - Contact Role|Finding|false|false||unknown
null|Unknown - Living Dependency|Finding|false|false||unknownnull|Ethnic group unknown|Subject|false|false||unknownnull|Unknown - Allergy Severity|Modifier|false|false||unknown
null|Unknown - HL7 update mode|Modifier|false|false||unknown
null|Unknown|Modifier|false|false||unknownnull|Science of Etiology|Finding|false|false||cause
null|Etiology aspects|Finding|false|false||causenull|Early|Time|false|false||earlynull|DFFB protein, human|Drug|true|false||CAD
null|DFFB protein, human|Drug|true|false||CADnull|Cold Hemagglutinin Disease|Disorder|true|false||CAD
null|Coronary heart disease|Disorder|true|false||CAD
null|Coronary Artery Disease|Disorder|true|false||CADnull|CAD gene|Finding|true|false||CAD
null|CALD1 wt Allele|Finding|true|false||CAD
null|B4GALNT2 gene|Finding|true|false||CAD
null|DFFB wt Allele|Finding|true|false||CAD
null|ACOD1 gene|Finding|true|false||CAD
null|DFFB gene|Finding|true|false||CADnull|cytarabine/daunorubicin protocol|Procedure|true|false||CAD
null|Computer Assisted Diagnosis|Procedure|true|false||CAD
null|Collision-Induced Dissociation|Procedure|true|false||CAD
null|CyADIC regimen|Procedure|true|false||CADnull|Caddo language|Entity|true|false||CADnull|Sudden Cardiac Death|Finding|true|false|C0018787|sudden cardiac deathnull|Sudden (qualifier value)|Modifier|false|false||suddennull|Cardiac Death|Finding|true|false|C0018787|cardiac deathnull|Cardiac attachment|Finding|false|false|C0018787|cardiacnull|Heart|Anatomy|false|false|C0376297;C1314974;C0085298|cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||cardiacnull|Event Consequence - Death|Finding|false|false||death
null|Death (finding)|Finding|false|false||death
null|Cessation of life|Finding|false|false||deathnull|Known|Modifier|false|false||knownnull|Medical History|Finding|true|false||history ofnull|History of present illness (finding)|Finding|true|false||history
null|History of previous events|Finding|true|false||history
null|Historical aspects qualifier|Finding|true|false||history
null|Medical History|Finding|true|false||history
null|Concept History|Finding|true|false||historynull|History|Subject|false|false||historynull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|physical examination (physical finding)|Finding|false|false||PHYSICAL EXAMnull|Physical Examination|Procedure|false|false||PHYSICAL EXAMnull|physical examination (physical finding)|Finding|false|false||PHYSICAL
null|Physical|Finding|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||PHYSICALnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Generalnull|General medical service|Procedure|false|false||Generalnull|Generalized|Modifier|false|false||Generalnull|Pleasant|Finding|false|false||Pleasantnull|Affect (mental function)|Finding|false|false||affectnull|assessment of affect|Procedure|false|false||affectnull|BORNHOLM EYE DISEASE|Disorder|false|false||bednull|Bachelor of Education|Finding|false|false||bednull|Beds|Device|false|false||bednull|Patient Location - Bed|Modifier|false|false||bednull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|HEENT|Anatomy|false|false||HEENTnull|Scleral Diseases|Disorder|false|false|C0036410|Scleranull|examination of sclera|Procedure|false|false|C0036410|Scleranull|Sclera|Anatomy|false|false|C0036412;C0026987;C0205180;C2228481|Scleranull|Anicteric|Finding|false|false|C0036410|anictericnull|Myelofibrosis|Disorder|false|false|C0694605;C0036410|MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false|C0026987|MMMnull|Oropharyngeal|Anatomy|false|false|C1550016|oropharynxnull|Remote control command - Clear|Finding|false|false|C0521367|clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Pupil equal round and reacting to light|Finding|false|false||PERRLnull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|Neck
null|Neck problem|Finding|false|false|C0027530;C3159206|Necknull|dendritic spine neck|Anatomy|false|false|C0812434;C0684335|Neck
null|Neck|Anatomy|false|false|C0812434;C0684335|Necknull|Supple|Finding|false|false||Supplenull|Jugular venous pressure|Finding|false|false||JVPnull|Regular|Modifier|false|false||Regularnull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Rhythm|Finding|false|false||rhythm
null|rhythmic process (biological)|Finding|false|false||rhythmnull|Heart murmur|Finding|true|false||murmursnull|Pericardial friction rub|Finding|true|false||rubsnull|Lung|Anatomy|false|false||Lungsnull|Minimal|Modifier|false|false||Minimal
null|Mild (qualifier value)|Modifier|false|false||Minimal
null|Minimum|Modifier|false|false||Minimalnull|Basilar Rales|Finding|false|false||crackles
null|Rales|Finding|false|false||cracklesnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|Abdomennull|Abdomen problem|Finding|false|false|C0230168;C0000726|Abdomennull|Abdomen|Anatomy|false|false|C0941288;C0153662|Abdomen
null|Abdominal Cavity|Anatomy|false|false|C0941288;C0153662|Abdomennull|Obese abdomen|Finding|false|false|C0230168;C0000726|obese abdomennull|Obesity|Disorder|false|false|C0230168;C0000726|obesenull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|abdomennull|Abdomen problem|Finding|false|false|C0230168;C0000726|abdomennull|Abdomen|Anatomy|false|false|C0426650;C0153662;C0941288;C0028754|abdomen
null|Abdominal Cavity|Anatomy|false|false|C0426650;C0153662;C0941288;C0028754|abdomennull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|Protective muscle spasm|Finding|false|false||guardingnull|Hereditary Multiple Exostoses|Disorder|false|false||Extnull|EXT1 wt Allele|Finding|false|false||Ext
null|EXT1 gene|Finding|false|false||Extnull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Posterior part of right leg|Anatomy|false|false|C0013604;C0038999|right calfnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Swollen calf|Finding|false|false|C0230445;C1305418|calf swellingnull|Structure of calf of leg|Anatomy|false|false|C0238882|calf
null|null|Anatomy|false|false|C0238882|calfnull|Cattle calf (organism)|Entity|false|false||calfnull|Swelling|Finding|false|false|C0489801|swelling
null|Edema|Finding|false|false|C0489801|swellingnull|Greater|LabModifier|false|false||greaternull|Posterior part of left leg|Anatomy|false|false|C0238882;C1552822;C0013604;C0038999|left calfnull|Table Cell Horizontal Align - left|Finding|false|false|C0489800|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Swollen calf|Finding|false|false|C0230445;C1305418;C0489800|calf swellingnull|Structure of calf of leg|Anatomy|false|false|C0238882|calf
null|null|Anatomy|false|false|C0238882|calfnull|Cattle calf (organism)|Entity|false|false||calfnull|Swelling|Finding|false|false|C0489800|swelling
null|Edema|Finding|false|false|C0489800|swellingnull|CALF TENDERNESS|Finding|true|false|C0230445;C1305418|calf tendernessnull|Structure of calf of leg|Anatomy|false|false|C0684239;C0234233;C0238883|calf
null|null|Anatomy|false|false|C0684239;C0234233;C0238883|calfnull|Cattle calf (organism)|Entity|true|false||calfnull|Emotional tenderness|Finding|true|false|C0230445;C1305418|tenderness
null|Sore to touch|Finding|true|false|C0230445;C1305418|tendernessnull|Palpation|Procedure|false|false||palpationnull|Thick|Modifier|false|false||Thicknull|Structure of nail of toe|Anatomy|false|false|C1546781;C0444099;C0151908;C0043345;C0178298;C0496955|toenailsnull|Dry Skin brand of emollient|Drug|false|false|C1123023;C4520765|dry skinnull|Xeroderma|Disorder|false|false|C0040357;C4299090;C1123023;C4520765;C0222007|dry skinnull|Dry skin|Finding|false|false|C1123023;C4520765;C0040357;C4299090;C0222007|dry skinnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C0040357;C4299090;C1123023;C4520765;C0222007|skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C0040357;C4299090;C1123023;C4520765;C0222007|skinnull|Skin Specimen Source Code|Finding|false|false|C0222007;C0040357;C4299090;C1123023;C4520765|skin
null|Skin Specimen|Finding|false|false|C0222007;C0040357;C4299090;C1123023;C4520765|skinnull|Skin, Human|Anatomy|false|false|C0151908;C0043345;C0720057;C1546781;C0444099;C0178298;C0496955|skin
null|Skin|Anatomy|false|false|C0151908;C0043345;C0720057;C1546781;C0444099;C0178298;C0496955|skinnull|Lower extremity>Toes|Anatomy|false|false|C0151908;C0043345;C1546781;C0444099;C0178298;C0496955|toes
null|Toes|Anatomy|false|false|C0151908;C0043345;C1546781;C0444099;C0178298;C0496955|toesnull|Congenital hallux valgus|Disorder|false|false|C0018534|Hallux valgus
null|Hallux Valgus|Disorder|false|false|C0018534|Hallux valgus
null|Acquired hallux valgus|Disorder|false|false|C0018534|Hallux valgusnull|Hallux structure|Anatomy|false|false|C0018536;C0158458;C0265656;C0042282|Halluxnull|Valgus deformity|Disorder|false|false|C0018534|valgusnull|Valgus <Valginae>|Entity|false|false||valgusnull|Valgus position|Modifier|false|false||valgusnull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Strength (attribute)|Finding|false|false|C0278454;C0015385;C0023216|strengthnull|Pharmaceutical Strength|LabModifier|false|false||strength
null|Physical Strength|LabModifier|false|false||strengthnull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Lower Extremity|Anatomy|false|false|C0808080|lower extremitiesnull|Body Site Modifier - Lower|Anatomy|false|false|C2003888|lowernull|Lower (action)|Event|false|false|C1548802;C0278454;C0015385|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|All extremities|Anatomy|false|false|C2003888;C0808080|extremities
null|Limb structure|Anatomy|false|false|C2003888;C0808080|extremitiesnull|Observation of Sensation|Finding|false|false||sensation
null|Sensory perception|Finding|false|false||sensationnull|sensory exam|Procedure|false|false||sensationnull|Sensation quality|Modifier|false|false||sensationnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|physical examination (physical finding)|Finding|false|false||PHYSICAL EXAMnull|Physical Examination|Procedure|false|false||PHYSICAL EXAMnull|physical examination (physical finding)|Finding|false|false||PHYSICAL
null|Physical|Finding|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||PHYSICALnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|Tmax|LabModifier|false|false||Tmaxnull|Saturation of Peripheral Oxygen|Attribute|false|false||SpO2null|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Generalnull|General medical service|Procedure|false|false||Generalnull|Generalized|Modifier|false|false||Generalnull|Pleasant|Finding|false|false||Pleasantnull|Affect (mental function)|Finding|false|false||affectnull|assessment of affect|Procedure|false|false||affectnull|BORNHOLM EYE DISEASE|Disorder|false|false||bednull|Bachelor of Education|Finding|false|false||bednull|Beds|Device|false|false||bednull|Patient Location - Bed|Modifier|false|false||bednull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|HEENT|Anatomy|false|false||HEENTnull|Scleral Diseases|Disorder|false|false|C0036410|Scleranull|examination of sclera|Procedure|false|false|C0036410|Scleranull|Sclera|Anatomy|false|false|C2228481;C0205180;C0036412;C0026987|Scleranull|Anicteric|Finding|false|false|C0036410|anictericnull|Myelofibrosis|Disorder|false|false|C0694605;C0036410|MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false|C0026987|MMMnull|Oropharyngeal|Anatomy|false|false|C1550016|oropharynxnull|Remote control command - Clear|Finding|false|false|C0521367|clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Pupil equal round and reacting to light|Finding|false|false||PERRLnull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|Neck
null|Neck problem|Finding|false|false|C0027530;C3159206|Necknull|dendritic spine neck|Anatomy|false|false|C0812434;C0684335|Neck
null|Neck|Anatomy|false|false|C0812434;C0684335|Necknull|Supple|Finding|false|false||Supplenull|Jugular venous pressure|Finding|false|false||JVPnull|Regular|Modifier|false|false||Regularnull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Rhythm|Finding|false|false||rhythm
null|rhythmic process (biological)|Finding|false|false||rhythmnull|Heart murmur|Finding|true|false||murmursnull|Pericardial friction rub|Finding|true|false||rubsnull|Lung|Anatomy|false|false||Lungsnull|Remote control command - Clear|Finding|false|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Auscultation|Procedure|false|false||auscultationnull|Wheezing|Finding|true|false||wheezesnull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|Abdomennull|Abdomen problem|Finding|false|false|C0230168;C0000726|Abdomennull|Abdomen|Anatomy|false|false|C0941288;C0153662|Abdomen
null|Abdominal Cavity|Anatomy|false|false|C0941288;C0153662|Abdomennull|Obese abdomen|Finding|false|false|C0230168;C0000726|obese abdomennull|Obesity|Disorder|false|false|C0230168;C0000726|obesenull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|abdomennull|Abdomen problem|Finding|false|false|C0230168;C0000726|abdomennull|Abdomen|Anatomy|false|false|C0941288;C0028754;C0426650;C0153662|abdomen
null|Abdominal Cavity|Anatomy|false|false|C0941288;C0028754;C0426650;C0153662|abdomennull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|Protective muscle spasm|Finding|false|false||guardingnull|Hereditary Multiple Exostoses|Disorder|false|false||Extnull|EXT1 wt Allele|Finding|false|false||Ext
null|EXT1 gene|Finding|false|false||Extnull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsenull|Pulse taking|Procedure|false|false||pulsenull|Pulse Rate|Attribute|false|false||pulsenull|Pulse phenomenon|Phenomenon|false|false||pulsenull|Physiologic pulse|Finding|false|false||pulsenull|Pulse taking|Procedure|false|false||pulsenull|Pulse Rate|Attribute|false|false||pulsenull|Pulse phenomenon|Phenomenon|false|false||pulsenull|null|Finding|false|false||radial pulsenull|examination of radial pulses|Procedure|false|false||radial pulsenull|Radial|Finding|false|false||radial
null|Circumpennate|Finding|false|false||radialnull|Pulse Wave Normal|Finding|false|false||pulse 2+null|Physiologic pulse|Finding|false|false||pulsenull|Pulse taking|Procedure|false|false||pulsenull|Pulse Rate|Attribute|false|false||pulsenull|Pulse phenomenon|Phenomenon|false|false||pulsenull|null|Finding|false|false||radial pulsenull|examination of radial pulses|Procedure|false|false||radial pulsenull|Radial|Finding|false|false||radial
null|Circumpennate|Finding|false|false||radialnull|Pulse Wave Decreased|Finding|false|false||pulse 1+null|Physiologic pulse|Finding|false|false||pulsenull|Pulse taking|Procedure|false|false||pulsenull|Pulse Rate|Attribute|false|false||pulsenull|Pulse phenomenon|Phenomenon|false|false||pulsenull|Mild Severity of Illness Code|Finding|false|false|C0230445;C1305418;C0489801|mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Posterior part of right leg|Anatomy|false|false|C1552823;C0238882;C0013604;C0038999;C1547225|right calfnull|Table Cell Horizontal Align - right|Finding|false|false|C0489801;C0230445;C1305418|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Swollen calf|Finding|false|false|C0230445;C1305418;C0489801|calf swellingnull|Structure of calf of leg|Anatomy|false|false|C0238882;C0013604;C0038999;C1547225;C1552823|calf
null|null|Anatomy|false|false|C0238882;C0013604;C0038999;C1547225;C1552823|calfnull|Cattle calf (organism)|Entity|false|false||calfnull|Swelling|Finding|false|false|C0230445;C1305418;C0489801|swelling
null|Edema|Finding|false|false|C0230445;C1305418;C0489801|swellingnull|Greater Than|LabModifier|false|false||greater thannull|Greater|LabModifier|false|false||greaternull|Posterior part of left leg|Anatomy|false|false|C1552822|left calfnull|Table Cell Horizontal Align - left|Finding|false|false|C0230445;C1305418;C0489800|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Swollen calf|Finding|false|false|C0230445;C1305418|calf swellingnull|Structure of calf of leg|Anatomy|false|false|C0238882;C1552822|calf
null|null|Anatomy|false|false|C0238882;C1552822|calfnull|Cattle calf (organism)|Entity|false|false||calfnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|CALF TENDERNESS|Finding|true|false|C0230445;C1305418|calf tendernessnull|Structure of calf of leg|Anatomy|false|false|C0684239;C0234233;C0238883|calf
null|null|Anatomy|false|false|C0684239;C0234233;C0238883|calfnull|Cattle calf (organism)|Entity|false|false||calfnull|Emotional tenderness|Finding|true|false|C0230445;C1305418|tenderness
null|Sore to touch|Finding|true|false|C0230445;C1305418|tendernessnull|Palpation|Procedure|false|false||palpationnull|Administration Method - Pain|Finding|true|false|C4299097;C0016504|pain
null|Pain|Finding|true|false|C4299097;C0016504|painnull|null|Attribute|true|false||painnull|Palpation|Procedure|false|false||palpationnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Dorsal|Modifier|false|false||dorsalnull|Lateral|Modifier|false|false||lateralnull|Foot problem|Finding|false|false|C4299097;C0016504|footnull|Lower extremity>Foot|Anatomy|false|false|C0555980;C1549543;C0030193|foot
null|Foot|Anatomy|false|false|C0555980;C1549543;C0030193|footnull|Foot Unit of Length|LabModifier|false|false||footnull|Skin callus|Disorder|false|false|C4299097;C0016504|callousnull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Lateral to the left|Modifier|false|false||left lateralnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Lateral|Modifier|false|false||lateralnull|Foot problem|Finding|false|false|C4299097;C0016504|footnull|Lower extremity>Foot|Anatomy|false|false|C0555980;C0376154|foot
null|Foot|Anatomy|false|false|C0555980;C0376154|footnull|Foot Unit of Length|LabModifier|false|false||footnull|Thick toenails|Finding|false|false|C0222007|Thick toenailsnull|Thick|Modifier|false|false||Thicknull|Structure of nail of toe|Anatomy|false|false|C1546781;C0444099;C0178298;C0496955;C4540337|toenailsnull|Dry Skin brand of emollient|Drug|false|false|C1123023;C4520765|dry skinnull|Xeroderma|Disorder|false|false|C1123023;C4520765|dry skinnull|Dry skin|Finding|false|false|C1123023;C4520765|dry skinnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C0222007;C1123023;C4520765|skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C0222007;C1123023;C4520765|skinnull|Skin Specimen Source Code|Finding|false|false|C0222007;C1123023;C4520765|skin
null|Skin Specimen|Finding|false|false|C0222007;C1123023;C4520765|skinnull|Skin, Human|Anatomy|false|false|C0043345;C0151908;C0178298;C0496955;C0720057;C1546781;C0444099|skin
null|Skin|Anatomy|false|false|C0043345;C0151908;C0178298;C0496955;C0720057;C1546781;C0444099|skinnull|Lower extremity>Toes|Anatomy|false|false||toes
null|Toes|Anatomy|false|false||toesnull|indurated|Finding|false|false|C0446523;C0694648;C1550235|induratednull|Cone-Rod Dystrophy 2|Disorder|false|false|C1550235;C0694648;C1549091;C0836913;C0446523|cordnull|Cord - Body Parts|Anatomy|false|false|C3489532;C0702114;C1552822|cordnull|Cord Device|Device|false|false||cordnull|left antecubital fossa|Anatomy|false|false|C3489532;C0702114;C1552822|left antecubital fossanull|Table Cell Horizontal Align - left|Finding|false|false|C0446523;C0836913;C0694648;C1550235|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Antecubital Fossa|Anatomy|false|false|C1552822;C0702114;C3489532|antecubital fossanull|Antecubital|Anatomy|false|false|C3489532|antecubitalnull|Fossa|Anatomy|false|false|C1552822;C3489532|fossanull|Fossa <Euplerinae>|Entity|false|false||fossa
null|Cryptoprocta ferox|Entity|false|false||fossanull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|Alert brand of caffeine|Drug|false|false||alert
null|Alert brand of caffeine|Drug|false|false||alertnull|Mentally alert|Finding|false|false||alert
null|Consciousness clear|Finding|false|false||alert
null|Alert note|Finding|false|false||alert
null|Alert|Finding|false|false||alertnull|null|Attribute|false|false||alertnull|Oriented to place|Finding|false|false||orientednull|Orientation, Spatial|Modifier|false|false||orientednull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Ruta graveolens preparation|Drug|false|false||RUE
null|Ruta graveolens preparation|Drug|false|false||RUEnull|Ruta graveolens|Entity|false|false||RUE
null|Ruta|Entity|false|false||RUEnull|Strength (attribute)|Finding|false|false||strengthnull|Pharmaceutical Strength|LabModifier|false|false||strength
null|Physical Strength|LabModifier|false|false||strengthnull|heme iron polypeptide|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|ST13 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|ST13 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|RPL29 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|RPL29 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|HHIP protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|HHIP protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|heme iron polypeptide|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hipnull|RPL29 wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C1879367|hip
null|REG3A gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C1879367|hip
null|RPL29 gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C1879367|hip
null|ST13 wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C1879367|hip
null|ST13 gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C1879367|hip
null|HHIP gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C1879367|hip
null|HHIP wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C1879367|hip
null|REG3A wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C1879367|hipnull|Procedure on hip|Procedure|false|false|C1879367;C0022122;C0228391;C0019552;C4299095|hipnull|Lower extremity>Hip|Anatomy|false|false|C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1430701;C0529134;C1505163;C1654726;C1292890;C0808080|hip
null|Hip structure|Anatomy|false|false|C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1430701;C0529134;C1505163;C1654726;C1292890;C0808080|hip
null|Structure of habenulopeduncular tract|Anatomy|false|false|C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1430701;C0529134;C1505163;C1654726;C1292890;C0808080|hip
null|Bone structure of ischium|Anatomy|false|false|C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1430701;C0529134;C1505163;C1654726;C1292890;C0808080|hipnull|Flexor (Anatomical coordinate)|Anatomy|false|false|C1292890;C0808080;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725|flexornull|Flexor <Diplocrepinae>|Entity|false|false||flexornull|Strength (attribute)|Finding|false|false|C1879367;C0022122;C0228391;C0019552;C4299095|strengthnull|Pharmaceutical Strength|LabModifier|false|false||strength
null|Physical Strength|LabModifier|false|false||strengthnull|Plantar (qualifier value)|Anatomy|false|false||plantar
null|Sole of Foot|Anatomy|false|false||plantarnull|null|Finding|false|false|C1548802;C0023216;C0278454;C0015385|flexionnull|W flexion|Attribute|false|false|C0023216;C1548802|flexionnull|Bilateral|Modifier|false|false||bilateralnull|Lower Extremity|Anatomy|false|false|C1552823;C2003888;C1525443;C0231452|lower extremitiesnull|Body Site Modifier - Lower|Anatomy|false|false|C2003888;C0231452;C1525443|lowernull|Lower (action)|Event|false|false|C1548802;C0023216;C0278454;C0015385|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|All extremities|Anatomy|false|false|C2003888;C0231452|extremities
null|Limb structure|Anatomy|false|false|C2003888;C0231452|extremitiesnull|Table Cell Horizontal Align - right|Finding|false|false|C0023216|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Body Site Modifier - Lower|Anatomy|false|false|C2003888|lowernull|Lower (action)|Event|false|false|C1548802|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Limb structure|Anatomy|false|false||extremitynull|Legal fine|Entity|false|false||finenull|Fine (qualifier value)|Modifier|false|false||finenull|Touch sensation|Finding|false|false||touch sensationnull|Touch sensation|Finding|false|false||touch
null|Touch Perception|Finding|false|false||touchnull|Therapeutic Touch|Procedure|false|false||touchnull|Tactile|Modifier|false|false||touchnull|Observation of Sensation|Finding|false|false|C0278454;C0015385|sensation
null|Sensory perception|Finding|false|false|C0278454;C0015385|sensationnull|sensory exam|Procedure|false|false|C0278454;C0015385|sensationnull|Sensation quality|Modifier|false|false||sensationnull|All extremities|Anatomy|false|false|C0036658;C0542538;C2229507|extremities
null|Limb structure|Anatomy|false|false|C0036658;C0542538;C2229507|extremitiesnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0851353;C0005768;C0229664;C0005767|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Lymph|Finding|false|false||Lymphsnull|Monos|Drug|false|false||Monos
null|Mono-S|Drug|false|false||Monos
null|Monos|Drug|false|false||Monosnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||Eos
null|Familial eosinophilia|Disorder|false|false||Eosnull|PRSS33 gene|Finding|false|false||Eos
null|IKZF4 gene|Finding|false|false||Eosnull|Eos <Loriini>|Entity|false|false||Eosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Thyrotropin-Releasing Hormone, human|Drug|false|false||TRF
null|IL5 protein, human|Drug|false|false||TRF
null|IL5 protein, human|Drug|false|false||TRF
null|thyrotropin-releasing hormone|Drug|false|false||TRF
null|thyrotropin-releasing hormone|Drug|false|false||TRF
null|thyrotropin-releasing hormone|Drug|false|false||TRF
null|Tocotrienol-rich Fraction|Drug|false|false||TRF
null|Thyrotropin-Releasing Hormone, human|Drug|false|false||TRFnull|TERF1 wt Allele|Finding|false|false||TRF
null|TERF1 gene|Finding|false|false||TRF
null|IL5 gene|Finding|false|false||TRFnull|Laboratory test finding|Lab|false|false||LABSnull|Imaging problem|Finding|false|false||IMAGINGnull|Diagnostic Imaging|Procedure|false|false||IMAGING
null|Imaging Techniques|Procedure|false|false||IMAGINGnull|Imaging Technology|Title|false|false||IMAGINGnull|Packed red blood cells|Drug|false|false||pRBCs
null|Packed red blood cells|Drug|false|false||pRBCsnull|On admission|Time|false|false||on admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0851353;C0005768;C0229664;C0005767|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|Episode of|Time|false|false||episode ofnull|Episode of|Time|false|false||episodenull|Coffee ground vomiting|Finding|false|false||coffee ground emesis
null|Vomit contains coffee grounds (finding)|Finding|false|false||coffee ground emesisnull|Coffee|Drug|false|false||coffeenull|Coffea <Coffeeae>|Entity|false|false||coffeenull|Emesis [PE]|Finding|false|false||emesis
null|Vomiting|Finding|false|false||emesis
null|Vomitus|Finding|false|false||emesisnull|Emesis <Emesidini>|Entity|false|false||emesis
null|Emesis <subgenus>|Entity|false|false||emesisnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0005768;C0229664;C0005767;C0851353|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0851353;C0005768;C0229664;C0005767|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C0014792;C1114281|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Bilateral|Modifier|false|false||bilateralnull|Lower Extremity|Anatomy|false|false|C0554756|lower extremitynull|Body Site Modifier - Lower|Anatomy|false|false|C2003888|lowernull|Lower (action)|Event|false|false|C1548802|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Limb structure|Anatomy|false|false|C0554756|extremitynull|Doppler studies|Procedure|false|false|C0015385;C0023216|dopplernull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Deep Vein Thrombosis|Disorder|false|false|C0042449;C0040184|Deep venous thrombosisnull|Deep Resection Margin|Attribute|false|false||Deepnull|Deep (qualifier value)|Modifier|false|false||Deepnull|Venous thrombosis after immobility|Finding|false|false|C0040184;C0042449|venous thrombosis
null|Venous Thrombosis|Finding|false|false|C0040184;C0042449|venous thrombosisnull|Veins|Anatomy|false|false|C0149871;C0517555;C0042487|venousnull|Venous|Modifier|false|false||venousnull|Thrombosis|Finding|false|false|C0040184|thrombosisnull|Bilateral|Modifier|false|false||bilateralnull|Posterior pituitary disease|Disorder|false|false|C0040184|posteriornull|Dorsal|Modifier|false|false||posteriornull|Bone structure of tibia|Anatomy|false|false|C0517555;C0042487;C0751438;C0040053;C0149871|tibialnull|Procedure on vein|Procedure|false|false|C0042449|veinsnull|Veins|Anatomy|false|false|C0398102|veinsnull|Right sided|Modifier|false|false||right-sidednull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Cyst|Disorder|false|false||cystnull|SpecimenType - Cyst|Finding|false|false||cyst
null|null|Finding|false|false||cystnull|Cyst form of protozoa|Entity|false|false||cystnull|Esophagogastroduodenoscopy|Procedure|false|false||EGDnull|Small amount|LabModifier|false|false||Small amountnull|Small|LabModifier|false|false||Smallnull|Amount class - Amount|Finding|false|false||amountnull|Quantity|LabModifier|false|false||amountnull|Hematin|Drug|false|false||hematin
null|Hematin|Drug|false|false||hematinnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Ulceration|Finding|true|false||ulceration
null|Ulcer|Finding|true|false||ulcerationnull|Hemorrhage|Finding|false|false||bleedingnull|Junction Device|Device|false|false||junctionnull|Junctional|Modifier|false|false||junctionnull|Neoplasm of uncertain or unknown behavior of stomach|Disorder|false|false|C3714551;C0038351;C4266636|stomach
null|Stomach Diseases|Disorder|false|false|C3714551;C0038351;C4266636|stomach
null|Benign neoplasm of stomach|Disorder|false|false|C3714551;C0038351;C4266636|stomach
null|Carcinoma in situ of stomach|Disorder|false|false|C3714551;C0038351;C4266636|stomachnull|Stomach problem|Finding|false|false|C3714551;C0038351;C4266636|stomachnull|Procedure on stomach|Procedure|false|false|C3714551;C0038351;C4266636|stomachnull|Stomach structure|Anatomy|false|false|C0038354;C0496905;C0153943;C0154060;C0577027;C0872393|stomach
null|Abdomen>Stomach|Anatomy|false|false|C0038354;C0496905;C0153943;C0154060;C0577027;C0872393|stomach
null|Stomach|Anatomy|false|false|C0038354;C0496905;C0153943;C0154060;C0577027;C0872393|stomachnull|Diffuse|Modifier|false|false||Diffusenull|Erythema|Disorder|false|false||erythemanull|Superficial|Modifier|false|false||superficialnull|Ulcer|Finding|false|false||ulcerationsnull|Carcinoma in situ of stomach|Disorder|false|false|C3714551;C0038351;C4266636|stomach
null|Stomach Diseases|Disorder|false|false|C3714551;C0038351;C4266636|stomach
null|Benign neoplasm of stomach|Disorder|false|false|C3714551;C0038351;C4266636|stomach
null|Neoplasm of uncertain or unknown behavior of stomach|Disorder|false|false|C3714551;C0038351;C4266636|stomachnull|Stomach problem|Finding|false|false|C3714551;C0038351;C4266636|stomachnull|Procedure on stomach|Procedure|false|false|C3714551;C0038351;C4266636|stomachnull|Stomach structure|Anatomy|false|false|C0872393;C0332290;C0038354;C0496905;C0153943;C0154060;C0577027|stomach
null|Abdomen>Stomach|Anatomy|false|false|C0872393;C0332290;C0038354;C0496905;C0153943;C0154060;C0577027|stomach
null|Stomach|Anatomy|false|false|C0872393;C0332290;C0038354;C0496905;C0153943;C0154060;C0577027|stomachnull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false|C3714551;C0038351;C4266636|consistentnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Gastritis|Disorder|false|false||gastritisnull|Hemorrhage|Finding|true|false||bleedingnull|Medium (Substance)|Drug|false|false||Medium
null|Culture Media|Drug|false|false||Mediumnull|A Medium Amount of Time|Finding|false|false||Medium
null|Communications Media|Finding|false|false||Medium
null|A Medium Amount|Finding|false|false||Mediumnull|Message Waiting Priority - Medium|Modifier|false|false||Medium
null|medium exposure|Modifier|false|false||Mediumnull|Medium|LabModifier|false|false||Mediumnull|Hiatal Hernia|Disorder|false|false||hiatal hernianull|Hernia|Disorder|false|false||hernianull|Erythema|Disorder|false|false|C1947952;C0025148;C0013303;C0227300|Erythemanull|Superficial|Modifier|false|false||superficialnull|Ulcer|Finding|false|false|C0227300;C1947952;C0025148|ulcerationsnull|Duodenal ampulla|Anatomy|false|false|C0041582;C0041834|duodenal bulbnull|Duodenum|Anatomy|false|false|C0041834|duodenalnull|anatomical bulb|Anatomy|false|false|C0041834;C0041582|bulb
null|Medulla Oblongata|Anatomy|false|false|C0041834;C0041582|bulbnull|plant bulb|Entity|false|false||bulbnull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|Duodenitis|Disorder|false|false||duodenitis
null|Acute Enteritis of the Mouse Intestinal Tract|Disorder|false|false||duodenitisnull|Esophagogastroduodenoscopy|Procedure|false|false|C0013303|EGDnull|III (suffix)|Modifier|false|false||thirdnull|Third|LabModifier|false|false||thirdnull|part of|Modifier|false|false||part ofnull|Role Class - part|Finding|false|false|C0013303|partnull|Part|Modifier|false|false||partnull|Part Dosing Unit|LabModifier|false|false||partnull|Malignant neoplasm of duodenum|Disorder|false|false|C0013303|duodenum
null|Benign neoplasm of duodenum|Disorder|false|false|C0013303|duodenumnull|Duodenum|Anatomy|false|false|C0496869;C0153426;C0079304;C1552020|duodenumnull|Left upper extremity|Anatomy|false|false|C0041621;C1456803;C1315081;C0041618;C0220934;C1552822|Left upper extremitynull|Table Cell Horizontal Align - left|Finding|false|false|C0230330;C1140618|Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Upper Extremity|Anatomy|false|false|C0220934;C1315081;C0041618;C1552822;C0041621;C1456803|upper extremitynull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Limb structure|Anatomy|false|false|C1315081;C0041618;C0041621;C1456803;C0220934|extremitynull|Ultrasonic|Finding|false|false|C1140618;C0015385;C0230330|ultrasoundnull|Urological ultrasound|Procedure|false|false|C0230330;C0015385;C1140618|ultrasound
null|Ultrasonography|Procedure|false|false|C0230330;C0015385;C1140618|ultrasoundnull|ultrasound device|Device|false|false||ultrasoundnull|Ultrasonic Shockwave|Phenomenon|false|false|C0230330;C0015385;C1140618|ultrasound
null|Ultrasonics (sound)|Phenomenon|false|false|C0230330;C0015385;C1140618|ultrasoundnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false|C0226514;C0042449|evidencenull|Deep vein thrombosis of lower limb|Disorder|true|false|C0226514;C0042449|deep vein thrombosis
null|Deep Vein Thrombosis|Disorder|true|false|C0226514;C0042449|deep vein thrombosisnull|Structure of deep vein|Anatomy|false|false|C0040053;C0042487;C3887511;C0149871;C0340708|deep veinnull|Deep Resection Margin|Attribute|true|false||deepnull|Deep (qualifier value)|Modifier|false|false||deepnull|Venous Thrombosis|Finding|true|false|C0226514;C0042449|vein thrombosisnull|Veins|Anatomy|false|false|C0040053;C3887511;C0042487;C0149871;C0340708|veinnull|Thrombosis|Finding|true|false|C0226514;C0042449|thrombosisnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Limb structure|Anatomy|false|false||extremitynull|Probable diagnosis|Finding|false|false|C0446523;C0694648;C0836913|Likely
null|Probably|Finding|false|false|C0446523;C0694648;C0836913|Likelynull|Evolving|Finding|false|false|C0836913;C0694648;C0446523|evolvingnull|Hematoma|Finding|false|false|C0694648;C0446523;C0836913|hematomanull|left antecubital fossa|Anatomy|false|false|C1552822;C0332148;C0750492;C0018944;C0332253|left antecubital fossanull|Table Cell Horizontal Align - left|Finding|false|false|C0694648;C0446523|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Antecubital Fossa|Anatomy|false|false|C0332148;C0750492;C1552822;C0018944;C0332253|antecubital fossanull|Antecubital|Anatomy|false|false||antecubitalnull|Fossa|Anatomy|false|false|C0332253;C0332148;C0750492;C0018944|fossanull|Fossa <Euplerinae>|Entity|false|false||fossa
null|Cryptoprocta ferox|Entity|false|false||fossanull|CAT scan of head|Procedure|false|false|C0018670;C0152336|CT headnull|null|Attribute|false|false|C0018670;C0152336|CT headnull|Problems with head|Disorder|false|false|C0018670;C0152336|headnull|Procedure on head|Procedure|false|false|C0018670;C0152336|headnull|Structure of head of caudate nucleus|Anatomy|false|false|C0362076;C0202691;C0876917;C0881943|head
null|Head|Anatomy|false|false|C0362076;C0202691;C0876917;C0881943|headnull|Head Device|Device|false|false||headnull|Contrast Media|Drug|false|false||contrastnull|Contrast|Modifier|false|false||contrastnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|false|false||acutenull|Infarction|Finding|true|false||infarctionnull|Hemorrhage|Finding|false|false||hemorrhagenull|Fracture|Disorder|false|false||fracturesnull|Fractured|Finding|false|false||fracturesnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Laboratory test finding|Lab|false|false||LABSnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0851353;C0005768;C0229664;C0005767|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C0014792;C1114281|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|edetic acid|Drug|false|false||EDTA
null|edetic acid|Drug|false|false||EDTAnull|BRIEF Health Literacy Screening Tool|Finding|false|false||Brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||Briefnull|Brief|Time|false|false||Briefnull|Shortened|Modifier|false|false||Briefnull|Hospital course|Finding|false|false||Hospital Coursenull|null|Attribute|false|false||Hospital Coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||Coursenull|Referral category - Outpatient|Finding|false|false||Outpatient
null|Patient Class - Outpatient|Finding|false|false||Outpatientnull|Outpatients|Subject|false|false||Outpatientnull|Provider|Finding|false|false||Providersnull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Hypertensive disease|Disorder|false|false||HTNnull|Chronic Kidney Diseases|Disorder|false|false||CKDnull|Stage level 4|Finding|false|false||stage IVnull|Tumor stage|Attribute|false|false||stagenull|Stage|Time|false|false||stage
null|Phase|Time|false|false||stagenull|Peripheral Vascular Diseases|Disorder|false|false||PVDnull|Pomalidomide/Bortezomib/Dexamethasone Regimen|Procedure|false|false||PVDnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Superficial|Modifier|false|false||superficialnull|Lower extremity>Femoral artery|Anatomy|false|false|C0857160;C2003888;C2219779;C1552822|femoral artery
null|Structure of femoral artery|Anatomy|false|false|C0857160;C2003888;C2219779;C1552822|femoral arterynull|Femur|Anatomy|false|false||femoralnull|Arterial system|Anatomy|false|false|C1552822;C0857160;C2003888;C2219779|artery
null|Arteries|Anatomy|false|false|C1552822;C0857160;C2003888;C2219779|arterynull|Structure of left lower leg|Anatomy|false|false||lower left legnull|Body Site Modifier - Lower|Anatomy|false|false|C2003888|lowernull|Lower (action)|Event|false|false|C0226004;C0003842;C4299099;C0015801;C1548802|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|numbness of left leg|Finding|false|false|C1140621;C0023216;C0226004;C0003842;C4299099;C0015801;C0230443;C0230416|left leg numbnessnull|Structure of left lower leg|Anatomy|false|false|C2219779|left leg
null|Left lower extremity|Anatomy|false|false|C2219779|left legnull|Table Cell Horizontal Align - left|Finding|false|false|C0226004;C0003842;C4299099;C0015801|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Numbness in leg|Finding|false|false|C0226004;C0003842;C4299099;C0015801;C1140621;C0023216|leg numbnessnull|Lower Extremity|Anatomy|false|false|C2219779;C0857160|leg
null|Leg|Anatomy|false|false|C2219779;C0857160|legnull|Numbness|Finding|false|false||numbness
null|Hypesthesia|Finding|false|false||numbnessnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Bilateral|Modifier|false|false||bilateralnull|Deep thrombophlebitis|Disorder|false|false|C5239664|DVT
null|Deep Vein Thrombosis|Disorder|false|false|C5239664|DVTnull|area DVT|Anatomy|false|false|C2926618;C0149871;C0151950|DVTnull|null|Attribute|false|false|C5239664|DVTnull|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|Hemorrhage|Finding|false|false||bleedingnull|Event|Event|false|false||eventsnull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Esophagogastroduodenoscopy|Procedure|false|false||EGDnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Coffee|Drug|false|false||coffeenull|Coffea <Coffeeae>|Entity|false|false||coffeenull|Emesis [PE]|Finding|false|false||emesis
null|Vomiting|Finding|false|false||emesis
null|Vomitus|Finding|false|false||emesisnull|Emesis <Emesidini>|Entity|false|false||emesis
null|Emesis <subgenus>|Entity|false|false||emesisnull|Feces|Finding|false|false||stoolsnull|null|Attribute|false|false||stoolsnull|Stool seat|Device|false|false||stoolsnull|BRAF Gene Rearrangement|Disorder|false|false||positivenull|Rh Positive Blood Group|Finding|false|false||positive
null|Positive Finding|Finding|false|false||positive
null|Positive|Finding|false|false||positivenull|Positive Charge|Modifier|false|false||positivenull|Positive Number|LabModifier|false|false||positivenull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Rectal Dosage Form|Drug|false|false||rectalnull|Rectal Route of Administration|Finding|false|false||rectal
null|Rectal (intended site)|Finding|false|false||rectalnull|TUBE,RECTAL,24FR,PLASTIC B#6510|Device|false|false||rectalnull|rectal|Modifier|false|false||rectalnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Consent Type - Colonoscopy|Procedure|false|false||colonoscopy
null|colonoscopy|Procedure|false|false||colonoscopynull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Left upper arm structure|Anatomy|false|false|C0018944;C3495676;C1552822;C1824218;C3715044;C1522541;C5400986;C4761640|left arm
null|Left arm|Anatomy|false|false|C0018944;C3495676;C1552822;C1824218;C3715044;C1522541;C5400986;C4761640|left armnull|Table Cell Horizontal Align - left|Finding|false|false|C0230347;C5779993|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Anorectal Malformations|Disorder|false|false|C0230347;C5779993;C0446516;C1140618;C1269078|armnull|AKR1A1 wt Allele|Finding|false|false|C0446516;C1140618;C1269078;C0230347;C5779993|arm
null|ARMC9 gene|Finding|false|false|C0446516;C1140618;C1269078;C0230347;C5779993|armnull|Protocol Treatment Arm|Procedure|false|false|C0446516;C1140618;C1269078;C0230347;C5779993|arm
null|Axillary Reverse Mapping|Procedure|false|false|C0446516;C1140618;C1269078;C0230347;C5779993|arm
null|Study Arm|Procedure|false|false|C0446516;C1140618;C1269078;C0230347;C5779993|armnull|Upper arm|Anatomy|false|false|C1824218;C3715044;C3495676;C1522541;C5400986;C4761640|arm
null|null|Anatomy|false|false|C1824218;C3715044;C3495676;C1522541;C5400986;C4761640|arm
null|Upper Extremity|Anatomy|false|false|C1824218;C3715044;C3495676;C1522541;C5400986;C4761640|armnull|Hematoma|Finding|false|false|C0230347;C5779993|hematomanull|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Hematoma|Finding|false|false||hematomanull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Radial|Finding|false|false||radial
null|Circumpennate|Finding|false|false||radialnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Bilateral|Modifier|false|false||bilateralnull|Lower Extremity|Anatomy|false|false||lower extremitynull|Body Site Modifier - Lower|Anatomy|false|false|C2003888|lowernull|Lower (action)|Event|false|false|C1548802|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Limb structure|Anatomy|false|false||extremitynull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Diagnostic Service Section ID - Hematology|Finding|false|false||Hematologynull|diagnostic service sources hematology (procedure)|Procedure|false|false||Hematology
null|Hematology procedure|Procedure|false|false||Hematology
null|Hematologic Tests|Procedure|false|false||Hematologynull|hematology (field)|Title|false|false||Hematologynull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Left upper arm structure|Anatomy|false|false|C3495676;C1824218;C3715044;C1522541;C5400986;C4761640|left arm
null|Left arm|Anatomy|false|false|C3495676;C1824218;C3715044;C1522541;C5400986;C4761640|left armnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Anorectal Malformations|Disorder|false|false|C0230347;C5779993;C0446516;C1140618;C1269078|armnull|AKR1A1 wt Allele|Finding|false|false|C0230347;C5779993;C0446516;C1140618;C1269078|arm
null|ARMC9 gene|Finding|false|false|C0230347;C5779993;C0446516;C1140618;C1269078|armnull|Protocol Treatment Arm|Procedure|false|false|C0446516;C1140618;C1269078;C0230347;C5779993|arm
null|Axillary Reverse Mapping|Procedure|false|false|C0446516;C1140618;C1269078;C0230347;C5779993|arm
null|Study Arm|Procedure|false|false|C0446516;C1140618;C1269078;C0230347;C5779993|armnull|Upper arm|Anatomy|false|false|C1522541;C5400986;C4761640;C3495676;C1824218;C3715044|arm
null|null|Anatomy|false|false|C1522541;C5400986;C4761640;C3495676;C1824218;C3715044|arm
null|Upper Extremity|Anatomy|false|false|C1522541;C5400986;C4761640;C3495676;C1824218;C3715044|armnull|Hematoma|Finding|false|false||hematomanull|Slow|Modifier|false|false||slowlynull|Recommendation|Finding|false|false||recommendationsnull|Coumadin|Drug|false|false||coumadin
null|Coumadin|Drug|false|false||coumadinnull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|On discharge|Time|false|false||on dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Rehabilitation therapy|Procedure|false|false||rehabnull|More|LabModifier|false|false||morenull|Problem|Finding|false|false||problemnull|null|Attribute|false|false||problemnull|summary - ActRelationshipSubset|Finding|false|false||summary
null|Summary (document)|Finding|false|false||summarynull|Marketing basis - Transitional|Finding|false|false||transitionalnull|Transitional cell morphology|Modifier|false|false||transitionalnull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Hypertensive disease|Disorder|false|false||HTNnull|Chronic Kidney Diseases|Disorder|false|false||CKDnull|Stage level 4|Finding|false|false||stage IVnull|Tumor stage|Attribute|false|false||stagenull|Stage|Time|false|false||stage
null|Phase|Time|false|false||stagenull|Peripheral Vascular Diseases|Disorder|false|false||PVDnull|Pomalidomide/Bortezomib/Dexamethasone Regimen|Procedure|false|false||PVDnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Superficial femoral artery|Anatomy|false|false||superficial femoral arterynull|Superficial|Modifier|false|false||superficialnull|Lower extremity>Femoral artery|Anatomy|false|false||femoral artery
null|Structure of femoral artery|Anatomy|false|false||femoral arterynull|Femur|Anatomy|false|false||femoralnull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Structure of left lower leg|Anatomy|false|false||lower Left legnull|Body Site Modifier - Lower|Anatomy|false|false|C2003888|lowernull|Lower (action)|Event|false|false|C1548802|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|numbness of left leg|Finding|false|false|C1140621;C0023216;C0230443;C0230416|Left leg numbnessnull|Structure of left lower leg|Anatomy|false|false|C2219779|Left leg
null|Left lower extremity|Anatomy|false|false|C2219779|Left legnull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Numbness in leg|Finding|false|false|C1140621;C0023216|leg numbnessnull|Lower Extremity|Anatomy|false|false|C2219779;C0857160|leg
null|Leg|Anatomy|false|false|C2219779;C0857160|legnull|Numbness|Finding|false|false||numbness
null|Hypesthesia|Finding|false|false||numbnessnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Evening|Time|false|false||eveningnull|Ultrasonic|Finding|false|false|C0023216;C1548802|ultrasoundnull|Urological ultrasound|Procedure|false|false|C0278454;C0015385;C1548802;C0023216|ultrasound
null|Ultrasonography|Procedure|false|false|C0278454;C0015385;C1548802;C0023216|ultrasoundnull|ultrasound device|Device|false|false||ultrasoundnull|Ultrasonic Shockwave|Phenomenon|false|false|C0023216|ultrasound
null|Ultrasonics (sound)|Phenomenon|false|false|C0023216|ultrasoundnull|Bilateral|Modifier|false|false||bilateralnull|Lower Extremity|Anatomy|false|false|C0220934;C2003888;C0041621;C1456803;C1315081;C0041618|lower extremitiesnull|Body Site Modifier - Lower|Anatomy|false|false|C2003888;C0220934;C1315081;C0041618|lowernull|Lower (action)|Event|false|false|C1548802;C0023216|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|All extremities|Anatomy|false|false|C1315081;C0041618|extremities
null|Limb structure|Anatomy|false|false|C1315081;C0041618|extremitiesnull|Bilateral|Modifier|false|false||bilateralnull|Structure of posterior tibial vein|Anatomy|false|false|C0398102;C0149871;C0151950;C0751438;C2926618|posterior tibial veinsnull|Posterior pituitary disease|Disorder|false|false|C0447138;C0226832|posteriornull|Dorsal|Modifier|false|false||posteriornull|Tibial vein structure|Anatomy|false|false|C0398102;C0149871;C0151950;C0751438;C2926618|tibial veinsnull|Bone structure of tibia|Anatomy|false|false|C0149871;C0151950;C0398102|tibialnull|Procedure on vein|Procedure|false|false|C0447138;C5239664;C0226832;C0040184;C0042449|veinsnull|Veins|Anatomy|false|false|C0149871;C0151950;C0398102|veinsnull|Deep thrombophlebitis|Disorder|false|false|C0042449;C0447138;C0226832;C0040184;C5239664|DVT
null|Deep Vein Thrombosis|Disorder|false|false|C0042449;C0447138;C0226832;C0040184;C5239664|DVTnull|area DVT|Anatomy|false|false|C0398102;C2926618;C0149871;C0151950|DVTnull|null|Attribute|false|false|C5239664;C0447138;C0226832|DVTnull|Bilateral|Modifier|false|false||Bilateralnull|Deep thrombophlebitis|Disorder|false|false||DVTsnull|Clinical NEC (not elsewhere classified in LNC)|Finding|false|false||clinicalnull|Clinical|Modifier|false|false||clinicalnull|Aspects of signs|Finding|true|false||signs
null|Physical findings|Finding|true|false||signsnull|Manufactured sign|Device|true|false||signsnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|BRAF Gene Rearrangement|Disorder|false|false||positivenull|Rh Positive Blood Group|Finding|false|false||positive
null|Positive Finding|Finding|false|false||positive
null|Positive|Finding|false|false||positivenull|Positive Charge|Modifier|false|false||positivenull|Positive Number|LabModifier|false|false||positivenull|Bilateral|Modifier|false|false||bilateralnull|Deep thrombophlebitis|Disorder|false|false||DVTsnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|ANTICOAGULATION (finding)|Finding|false|false||anticoagulation
null|Anticoagulation function|Finding|false|false||anticoagulation
null|Decreased Coagulation Activity [PE]|Finding|false|false||anticoagulationnull|Anticoagulation Therapy|Procedure|false|false||anticoagulationnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|Therapeutic brand of coal tar|Drug|false|false||therapeutic
null|Therapeutic brand of coal tar|Drug|false|false||therapeuticnull|Therapeutic - Location Service Code|Finding|false|false||therapeutic
null|Therapeutic|Finding|false|false||therapeuticnull|Therapeutic procedure|Procedure|false|false||therapeuticnull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|Coagulation tissue factor induced.INR goal|Attribute|false|false||INR goalnull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|objective (goal)|Finding|false|false||goal
null|Act Mood - Goal|Finding|false|false||goalnull|Due to|Finding|false|false||Due
null|Due|Finding|false|false||Duenull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|Diagnostic Service Section ID - Hematology|Finding|false|false||hematologynull|diagnostic service sources hematology (procedure)|Procedure|false|false||hematology
null|Hematology procedure|Procedure|false|false||hematology
null|Hematologic Tests|Procedure|false|false||hematologynull|hematology (field)|Title|false|false||hematologynull|Further|Modifier|false|false||furthernull|heparin, porcine|Drug|false|false||Heparin
null|heparin, porcine|Drug|false|false||Heparin
null|heparin, porcine|Drug|false|false||Heparin
null|heparin|Drug|false|false||Heparin
null|heparin|Drug|false|false||Heparin
null|heparin|Drug|false|false||Heparinnull|clopidogrel|Drug|false|false||Clopidogrel
null|clopidogrel|Drug|false|false||Clopidogrelnull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Cardiologists|Subject|false|false||cardiologistnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|Appropriate|Modifier|false|false||appropriatenull|Screening for cancer|Procedure|false|false||cancer screeningnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Screening - procedure intent|Finding|false|false||screening
null|Special screening finding|Finding|false|false||screening
null|Aspects of disease screening|Finding|false|false||screeningnull|Screening for cancer|Procedure|false|false||screening
null|Disease Screening|Procedure|false|false||screening
null|research subject screening|Procedure|false|false||screening
null|Screening|Procedure|false|false||screening
null|Screening procedure|Procedure|false|false||screeningnull|Consent Type - Colonoscopy|Procedure|false|false||colonoscopy
null|colonoscopy|Procedure|false|false||colonoscopynull|Encounter due to Screening for malignant neoplasm of breast|Finding|false|false||mammogramnull|Mammography|Procedure|false|false||mammogramnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Clinic|Device|false|false||clinic
null|Ambulatory Care Facilities|Device|false|false||clinicnull|Clinic|Entity|false|false||clinic
null|Ambulatory Care Facilities|Entity|false|false||clinicnull|Patient location type - Clinic|Modifier|false|false||clinic
null|Person location type - Clinic|Modifier|false|false||clinicnull|ANTICOAGULATION (finding)|Finding|false|false||anticoagulation
null|Anticoagulation function|Finding|false|false||anticoagulation
null|Decreased Coagulation Activity [PE]|Finding|false|false||anticoagulationnull|Anticoagulation Therapy|Procedure|false|false||anticoagulationnull|Disease Management|Procedure|false|false||managementnull|Management Occupations|Subject|false|false||managementnull|Management procedure|Event|false|false||management
null|Administration occupational activities|Event|false|false||managementnull|on warfarin|Procedure|false|false||on warfarinnull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|3 Months|Time|false|false||3 monthsnull|month|Time|false|false||monthsnull|Upper gastrointestinal hemorrhage|Finding|false|false||Upper GI bleednull|Upper gastrointestinal tract series|Procedure|false|false||Upper GInull|Upper Surface|Modifier|false|false||Upper
null|Upper|Modifier|false|false||Uppernull|Gastrointestinal Hemorrhage|Finding|false|false||GI bleednull|Hemorrhage|Finding|false|false||bleednull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Episode of|Time|false|false||episodenull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|Coffee|Drug|false|false||coffeenull|Coffea <Coffeeae>|Entity|false|false||coffeenull|Emesis [PE]|Finding|false|false||emesis
null|Vomiting|Finding|false|false||emesis
null|Vomitus|Finding|false|false||emesisnull|Emesis <Emesidini>|Entity|false|false||emesis
null|Emesis <subgenus>|Entity|false|false||emesisnull|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Packed red blood cells|Drug|false|false||pRBCs
null|Packed red blood cells|Drug|false|false||pRBCsnull|Esophagogastroduodenoscopy|Procedure|false|false||EGDnull|Gastritis|Disorder|false|false||gastritisnull|Superficial|Modifier|false|false||superficialnull|Superficial ulcer|Disorder|false|false||erosionsnull|Erosion lesion|Finding|false|false||erosionsnull|Hemorrhage|Finding|true|false||bleedingnull|Incidental Findings|Finding|false|false||Incidental findingnull|Incidental|Finding|false|false||Incidentalnull|Experimental Finding|Finding|false|false||finding
null|Signs and Symptoms|Finding|false|false||finding
null|Finding|Finding|false|false||findingnull|Medium (Substance)|Drug|false|false||medium
null|Culture Media|Drug|false|false||mediumnull|A Medium Amount of Time|Finding|false|false||medium
null|Communications Media|Finding|false|false||medium
null|A Medium Amount|Finding|false|false||mediumnull|Message Waiting Priority - Medium|Modifier|false|false||medium
null|medium exposure|Modifier|false|false||mediumnull|Medium|LabModifier|false|false||mediumnull|Hiatal Hernia|Disorder|false|false||hiatal hernianull|Hernia|Disorder|false|false||hernianull|Feces|Finding|false|false||Stoolnull|Stool seat|Device|false|false||Stoolnull|Antigens|Drug|false|false||antigennull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|week|Time|false|false||weeksnull|High dose|LabModifier|false|false||high dosenull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Proton Pump Inhibitors|Drug|false|false||PPInull|Prepulse Inhibition|Finding|false|false||PPInull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Antecubital|Anatomy|false|false||antecubitalnull|Hematoma|Finding|false|false||hematomanull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Antecubital|Anatomy|false|false|C2959585;C0542559;C2183248;C0018944;C5552692;C0030605;C0190979;C0684257;C0031555|antecubitalnull|Hematoma|Finding|false|false|C1549091|hematomanull|contextual factors|Finding|false|false|C1549091|settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|diagnostic service sources phlebotomy|Finding|false|false|C1549091|phlebotomynull|Phlebotomy, therapeutic (separate procedure)|Procedure|false|false|C1549091|phlebotomy
null|Venous blood sampling|Procedure|false|false|C1549091|phlebotomy
null|Venesection|Procedure|false|false|C1549091|phlebotomynull|Proliferating trichilemmal tumor|Disorder|false|false|C1549091|PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false|C1549091|PTT
null|Partial Thromboplastin Time|Procedure|false|false|C1549091|PTTnull|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|Drops - Drug Form|Drug|false|false||gttnull|Gestational Trophoblastic Neoplasms|Disorder|false|false||gttnull|Glucose tolerance test|Procedure|false|false||gttnull|Drop Dosing Unit|LabModifier|false|false||gtt
null|Medical Drop|LabModifier|false|false||gttnull|heparin, porcine|Drug|false|false||Heparin
null|heparin, porcine|Drug|false|false||Heparin
null|heparin, porcine|Drug|false|false||Heparin
null|heparin|Drug|false|false||Heparin
null|heparin|Drug|false|false||Heparin
null|heparin|Drug|false|false||Heparinnull|Hematoma|Finding|false|false||hematomanull|Repeat Object|Finding|false|false||Repeat
null|Repeat|Finding|false|false||Repeatnull|Repeat Pattern|Time|false|false||Repeatnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Admission Level of Care Code - Acute|Finding|false|false||Acute
null|Acute - Triage Code|Finding|false|false||Acutenull|acute|Time|false|false||Acutenull|Chronic Kidney Diseases|Disorder|false|false||CKDnull|Stage level 4|Finding|false|false||Stage IVnull|Tumor stage|Attribute|false|false||Stagenull|Stage|Time|false|false||Stage
null|Phase|Time|false|false||Stagenull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|creatinine|Drug|false|false||creatinine
null|creatinine|Drug|false|false||creatininenull|Creatinine metabolic function|Finding|false|false||creatininenull|Creatinine measurement|Procedure|false|false||creatininenull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Hydration status|Finding|false|false||hydration
null|Hydration|Finding|false|false||hydrationnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|Lasix|Drug|false|false||lasix
null|Lasix|Drug|false|false||lasixnull|lisinopril|Drug|false|false||lisinopril
null|lisinopril|Drug|false|false||lisinoprilnull|Initially|Time|false|false||initiallynull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|Lasix|Drug|false|false||lasix
null|Lasix|Drug|false|false||lasixnull|On discharge|Time|false|false||on dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Daily|Time|false|false||dailynull|Anemia|Disorder|false|false||Anemianull|Anemia <Anemiaceae>|Entity|false|false||Anemianull|Has patient|Finding|false|false||Patient hasnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Anemia|Disorder|false|false||anemianull|Anemia <Anemiaceae>|Entity|false|false||anemianull|Rectal examination|Procedure|false|false||Rectal examnull|Rectal Dosage Form|Drug|false|false||Rectalnull|Rectal Route of Administration|Finding|false|false||Rectal
null|Rectal (intended site)|Finding|false|false||Rectalnull|TUBE,RECTAL,24FR,PLASTIC B#6510|Device|false|false||Rectalnull|rectal|Modifier|false|false||Rectalnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|guaiac|Drug|false|false||guaiac
null|guaiac|Drug|false|false||guaiacnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|EPO protein, human|Drug|false|false||EPO
null|epoetin alfa|Drug|false|false||EPO
null|epoetin alfa|Drug|false|false||EPO
null|Erythropoietin|Drug|false|false||EPO
null|Erythropoietin|Drug|false|false||EPO
null|Erythropoietin|Drug|false|false||EPO
null|EPO protein, human|Drug|false|false||EPOnull|EPO gene|Finding|false|false||EPO
null|TIMP1 wt Allele|Finding|false|false||EPO
null|EPX gene|Finding|false|false||EPO
null|TIMP1 gene|Finding|false|false||EPO
null|Exclusive Provider Organization Plan|Finding|false|false||EPOnull|Esperanto Language|Entity|false|false||EPOnull|Science of Etiology|Finding|false|false||Etiology
null|Etiology aspects|Finding|false|false||Etiology
null|Etiology|Finding|false|false||Etiologynull|Adverse Event Probably Related to Intervention|Modifier|false|false||likely relatednull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Relate - vinyl resin|Drug|false|false||relatednull|Role Link Type - related|Finding|false|false||related
null|Related (finding)|Finding|false|false||relatednull|Definitely Related to Intervention|Modifier|false|false||related
null|Relationships|Modifier|false|false||relatednull|Chronic Kidney Diseases|Disorder|false|false||CKDnull|Slow|Modifier|false|false||slownull|Gastrointestinal Hemorrhage|Finding|false|false||GI bleednull|Hemorrhage|Finding|false|false||bleednull|Has patient|Finding|false|false||patient hasnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Gastritis|Disorder|false|false||gastritisnull|Duodenitis|Disorder|false|false||duodenitis
null|Acute Enteritis of the Mouse Intestinal Tract|Disorder|false|false||duodenitisnull|Esophagogastroduodenoscopy|Procedure|false|false||EGDnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Hemorrhage|Finding|true|false||bleedingnull|iron studies|Procedure|false|false||Iron studiesnull|Iron Drug Class|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||Ironnull|Iron measurement|Procedure|false|false||Ironnull|Scientific Study|Procedure|false|false||studiesnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|furosemide|Drug|false|false||furosemide
null|furosemide|Drug|false|false||furosemidenull|lisinopril|Drug|false|false||Lisinopril
null|lisinopril|Drug|false|false||Lisinoprilnull|On admission|Time|false|false||on admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Gastrointestinal Hemorrhage|Finding|false|false||GI bleednull|Hemorrhage|Finding|false|false||bleednull|carvedilol|Drug|false|false||Carvedilol
null|carvedilol|Drug|false|false||Carvedilolnull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Table Frame - above|Finding|false|false||abovenull|Upper|Modifier|false|false||abovenull|nifedipine|Drug|false|false||Nifedipine
null|nifedipine|Drug|false|false||Nifedipinenull|BID protein, human|Drug|false|false||bid
null|BID protein, human|Drug|false|false||bidnull|Body integrity dysphoria|Disorder|false|false||bidnull|BID gene|Finding|false|false||bidnull|Twice a day|Time|false|false||bidnull|Lasix|Drug|false|false||lasix
null|Lasix|Drug|false|false||lasixnull|Daily|Time|false|false||dailynull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Burning Mouth Syndrome|Disorder|false|false||BMSnull|Circumflex|Modifier|false|false||circumflexnull|PROGRESSIVE ENCEPHALOMYELITIS WITH RIGIDITY|Disorder|false|false|C0449201|Pernull|Per - dosing instruction fragment|Finding|false|false|C0449201|Per
null|PER1 gene|Finding|false|false|C0449201|Per
null|Follow|Finding|false|false|C0449201|Per
null|PER1 wt Allele|Finding|false|false|C0449201|Pernull|PER (body structure)|Anatomy|false|false|C3273590;C4281991;C1418464;C1704764;C1861457|Pernull|Per (qualifier)|Modifier|false|false||Pernull|Discussion (procedure)|Procedure|false|false||discussionsnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Cardiologists|Subject|false|false||cardiologistnull|clopidogrel|Drug|false|false||clopidogrel
null|clopidogrel|Drug|false|false||clopidogrelnull|Gastrointestinal Hemorrhage|Finding|false|false||GI bleednull|Hemorrhage|Finding|false|false||bleednull|Transcription Initiation|Finding|false|false||initiation
null|Initiation|Finding|false|false||initiation
null|null|Finding|false|false||initiationnull|AOD use initiation|Time|false|false||initiationnull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|Lasix|Drug|false|false||Lasix
null|Lasix|Drug|false|false||Lasixnull|Initially|Time|false|false||initiallynull|Table Frame - above|Finding|false|false||abovenull|Upper|Modifier|false|false||abovenull|On discharge|Time|false|false||on dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Daily|Time|false|false||dailynull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|Arylsulfatase A, human|Drug|false|false||ASA
null|Arylsulfatase A, human|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASAnull|ARSA gene|Finding|false|false||ASAnull|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Drug|false|false||statin
null|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Drug|false|false||statinnull|EEF1A2 gene|Finding|false|false||statinnull|3-hydroxy-3-methylglutaryl-coenzyme A reductase inhibitor (disposition)|Modifier|false|false||statinnull|carvedilol|Drug|false|false||carvedilol
null|carvedilol|Drug|false|false||carvedilolnull|Hypertensive disease|Disorder|false|false||HTNnull|nifedipine|Drug|false|false||Nifedipine
null|nifedipine|Drug|false|false||Nifedipinenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Numerous|LabModifier|false|false||multiplenull|Bleeding episodes|Finding|false|false||bleeding episodesnull|Hemorrhage|Finding|false|false||bleedingnull|Episode of|Time|false|false||episodesnull|Systemic arterial pressure|Finding|false|false||blood pressuresnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Pressure (finding)|Finding|false|false||pressuresnull|null|Phenomenon|false|false||pressuresnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|carvedilol|Drug|false|false||carvedilol
null|carvedilol|Drug|false|false||carvedilolnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|nifedipine|Drug|false|false||nifedipine
null|nifedipine|Drug|false|false||nifedipinenull|Daily|Time|false|false||dailynull|Acute hemorrhage|Finding|false|false||acute bleednull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Hemorrhage|Finding|false|false||bleednull|Structure of subparietal sulcus|Anatomy|false|false||SBPsnull|Lasix|Drug|false|false||Lasix
null|Lasix|Drug|false|false||Lasixnull|Daily|Time|false|false||dailynull|Daily|Time|false|false||dailynull|Diabetes Mellitus|Disorder|false|false||Diabetes Mellitusnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Diabetes
null|Diabetes|Disorder|false|false||Diabetes
null|Diabetes Mellitus|Disorder|false|false||Diabetesnull|Patient Condition Code - Stable|Finding|false|false||Stablenull|Stable status|Modifier|false|false||Stablenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Unit - NCI Thesaurus Property|LabModifier|false|false||units
null|Unit of Measure|LabModifier|false|false||units
null|Unit|LabModifier|false|false||unitsnull|insulin, regular, human|Drug|false|false||insulin
null|Insulin [EPC]|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulinnull|INS gene|Finding|false|false||insulinnull|Insulin measurement|Procedure|false|false||insulinnull|Bedtime (qualifier value)|Time|false|false||bedtime
null|Once a day, at bedtime|Time|false|false||bedtimenull|Marketing basis - Transitional|Finding|false|false||TRANSITIONALnull|Transitional cell morphology|Modifier|false|false||TRANSITIONALnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Work-up|Procedure|false|false||work upnull|Work|Event|false|false||worknull|Screening - procedure intent|Finding|false|false||screening
null|Special screening finding|Finding|false|false||screening
null|Aspects of disease screening|Finding|false|false||screeningnull|research subject screening|Procedure|false|false||screening
null|Disease Screening|Procedure|false|false||screening
null|Screening|Procedure|false|false||screening
null|Screening for cancer|Procedure|false|false||screening
null|Screening procedure|Procedure|false|false||screeningnull|Consent Type - Colonoscopy|Procedure|false|false||colonoscopy
null|colonoscopy|Procedure|false|false||colonoscopynull|Last|Modifier|false|false||lastnull|Encounter due to Screening for malignant neoplasm of breast|Finding|false|false||mammogramnull|Mammography|Procedure|false|false||mammogramnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Course|Time|false|false||coursenull|High dose|LabModifier|false|false||high dosenull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Proton Pump Inhibitors|Drug|false|false||PPInull|Prepulse Inhibition|Finding|false|false||PPInull|pantoprazole|Drug|false|false||pantoprazole
null|pantoprazole|Drug|false|false||pantoprazolenull|Twice a day|Time|false|false||twice dailynull|Daily|Time|false|false||dailynull|End date|Time|false|false||end datenull|Endoglin, human|Drug|false|false||end
null|Endoglin, human|Drug|false|false||endnull|end - ActRelationshipCheckpoint|Finding|false|false||end
null|ENG gene|Finding|false|false||end
null|ENG wt Allele|Finding|false|false||endnull|Stop (qualifier value)|Time|false|false||endnull|End|Modifier|false|false||endnull|Upper gastrointestinal hemorrhage|Finding|false|false||upper GI bleednull|Upper gastrointestinal tract series|Procedure|false|false||upper GInull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Gastrointestinal Hemorrhage|Finding|false|false||GI bleednull|Hemorrhage|Finding|false|false||bleednull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Gastritis|Disorder|false|false||gastritisnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|hypertensive agents|Drug|false|false||hypertension medicationsnull|Hypertensive disease|Disorder|false|false||hypertensionnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|lisinopril|Drug|false|false||Lisinopril
null|lisinopril|Drug|false|false||Lisinoprilnull|nifedipine|Drug|false|false||nifedipine
null|nifedipine|Drug|false|false||nifedipinenull|Upper gastrointestinal hemorrhage|Finding|false|false||upper GI bleednull|Upper gastrointestinal tract series|Procedure|false|false||upper GInull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Gastrointestinal Hemorrhage|Finding|false|false||GI bleednull|Hemorrhage|Finding|false|false||bleednull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|furosemide|Drug|false|false||furosemide
null|furosemide|Drug|false|false||furosemidenull|Daily|Time|false|false||dailynull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|nifedipine|Drug|false|false||nifedipine
null|nifedipine|Drug|false|false||nifedipinenull|Daily|Time|false|false||dailynull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Hemorrhage|Finding|false|false|C0228216|bleednull|Structure of subparietal sulcus|Anatomy|false|false|C0019080|SBPsnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Coumadin|Drug|false|false||Coumadin
null|Coumadin|Drug|false|false||Coumadinnull|clopidogrel|Drug|false|false||Clopidogrel
null|clopidogrel|Drug|false|false||Clopidogrelnull|Cardiovascular system|Anatomy|false|false||cardiologynull|cardiology (field)|Title|false|false||cardiologynull|Cardiology service|Entity|false|false||cardiologynull|Arylsulfatase A, human|Drug|false|false||ASA
null|Arylsulfatase A, human|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASAnull|ARSA gene|Finding|false|false||ASAnull|MDF Attribute Type - Address|Finding|false|false||address
null|Address (property)|Finding|false|false||address
null|Address|Finding|false|false||address
null|Value type - Address|Finding|false|false||address
null|Addresses (publication format)|Finding|false|false||address
null|Address Data Type|Finding|false|false||addressnull|null|Attribute|false|false||addressnull|Patient's home|Device|false|false||patient's homenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|home environment (history)|Finding|false|false||home environmentnull|Home environment|Modifier|false|false||home environmentnull|Address type - Home|Finding|false|false||home
null|Visit User Code - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Home environment|Modifier|false|false||home
null|Person location type - Home|Modifier|false|false||homenull|Environment|Modifier|false|false||environmentnull|At increased risk for falls|Finding|false|false||fall risknull|Falls|Finding|false|false||fallnull|Autumn|Time|false|false||fallnull|Risk|Finding|false|false||risknull|Recent|Time|false|false||recentnull|triptorelin|Drug|false|false||trip
null|triptorelin|Drug|false|false||trip
null|triptorelin|Drug|false|false||tripnull|TRAIP wt Allele|Finding|false|false||trip
null|TRAIP gene|Finding|false|false||trip
null|PIK3IP1 gene|Finding|false|false||trip
null|LRRFIP1 gene|Finding|false|false||tripnull|Tripping|Phenomenon|false|false||tripnull|At home|Finding|false|false||at homenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|ANTICOAGULATION (finding)|Finding|false|false||anticoagulation
null|Anticoagulation function|Finding|false|false||anticoagulation
null|Decreased Coagulation Activity [PE]|Finding|false|false||anticoagulationnull|Anticoagulation Therapy|Procedure|false|false||anticoagulationnull|Has patient|Finding|false|false||patient hasnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Patient Class - Outpatient|Finding|false|false||outpatient
null|Referral category - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|ANTICOAGULATION (finding)|Finding|false|false||anticoagulation
null|Anticoagulation function|Finding|false|false||anticoagulation
null|Decreased Coagulation Activity [PE]|Finding|false|false||anticoagulationnull|Anticoagulation Therapy|Procedure|false|false||anticoagulationnull|Disease Management|Procedure|false|false||managementnull|Management Occupations|Subject|false|false||managementnull|Management procedure|Event|false|false||management
null|Administration occupational activities|Event|false|false||managementnull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Rehabilitation therapy|Procedure|false|false||rehabnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Accurate (qualifier value)|Modifier|false|false||accuratenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|lisinopril|Drug|false|false||Lisinopril
null|lisinopril|Drug|false|false||Lisinoprilnull|Daily|Time|false|false||DAILYnull|allopurinol|Drug|false|false||Allopurinol
null|allopurinol|Drug|false|false||Allopurinolnull|Daily|Time|false|false||DAILYnull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|carvedilol|Drug|false|false||Carvedilol
null|carvedilol|Drug|false|false||Carvedilolnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|clopidogrel|Drug|false|false||Clopidogrel
null|clopidogrel|Drug|false|false||Clopidogrelnull|Daily|Time|false|false||DAILYnull|furosemide|Drug|false|false||Furosemide
null|furosemide|Drug|false|false||Furosemidenull|Daily|Time|false|false||DAILYnull|ranitidine|Drug|false|false||Ranitidine
null|ranitidine|Drug|false|false||Ranitidinenull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Reflux|Finding|false|false||refluxnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||DAILYnull|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitaminsnull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|Daily|Time|false|false||DAILYnull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|Storage Unit|Device|false|false||UNIT
null|Unit device|Device|false|false||UNITnull|Unit - NCI Thesaurus Property|LabModifier|false|false||UNIT
null|Unit of Measure|LabModifier|false|false||UNIT
null|Unit|LabModifier|false|false||UNIT
null|Enzyme Unit|LabModifier|false|false||UNITnull|Daily|Time|false|false||DAILYnull|nifedipine|Drug|false|false||NIFEdipine
null|nifedipine|Drug|false|false||NIFEdipinenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|nitroglycerin|Drug|false|false||Nitroglycerin
null|nitroglycerin|Drug|false|false||Nitroglycerinnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0008031;C1549543;C0030193;C2926613;C0741025|chest
null|Anterior thoracic region|Anatomy|false|false|C0008031;C1549543;C0030193;C2926613;C0741025|chestnull|Administration Method - Pain|Finding|false|false|C1527391;C0817096|pain
null|Pain|Finding|false|false|C1527391;C0817096|painnull|null|Attribute|false|false||painnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Units
null|Unit of Measure|LabModifier|false|false||Units
null|Unit|LabModifier|false|false||Unitsnull|Dinner|Finding|false|false||Dinnernull|With dinner|Time|false|false||Dinnernull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|allopurinol|Drug|false|false||Allopurinol
null|allopurinol|Drug|false|false||Allopurinolnull|Transaction counts and value totals - day|Finding|false|false||DAY
null|Precision - day|Finding|false|false||DAYnull|Land Dayak Languages|Entity|false|false||DAYnull|day|Time|false|false||DAY
null|Daily|Time|false|false||DAYnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||DAILYnull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|carvedilol|Drug|false|false||Carvedilol
null|carvedilol|Drug|false|false||Carvedilolnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Units
null|Unit of Measure|LabModifier|false|false||Units
null|Unit|LabModifier|false|false||Unitsnull|Dinner|Finding|false|false||Dinnernull|With dinner|Time|false|false||Dinnernull|lisinopril|Drug|false|false||Lisinopril
null|lisinopril|Drug|false|false||Lisinoprilnull|Daily|Time|false|false||DAILYnull|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitaminsnull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|Daily|Time|false|false||DAILYnull|nifedipine|Drug|false|false||NIFEdipine
null|nifedipine|Drug|false|false||NIFEdipinenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|Storage Unit|Device|false|false||UNIT
null|Unit device|Device|false|false||UNITnull|Unit - NCI Thesaurus Property|LabModifier|false|false||UNIT
null|Unit of Measure|LabModifier|false|false||UNIT
null|Unit|LabModifier|false|false||UNIT
null|Enzyme Unit|LabModifier|false|false||UNITnull|Daily|Time|false|false||DAILYnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|gabapentin|Drug|false|false||Gabapentin
null|gabapentin|Drug|false|false||Gabapentinnull|Once a day, at bedtime|Time|false|false||QHSnull|Neuropathic pain|Finding|false|false||neuropathic pain
null|Neuralgia|Finding|false|false||neuropathic painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|pantoprazole|Drug|false|false||Pantoprazole
null|pantoprazole|Drug|false|false||Pantoprazolenull|Every twelve hours|Time|false|false||Q12Hnull|sennosides, USP|Drug|false|false||Senna
null|sennosides, USP|Drug|false|false||Sennanull|Senna alexandrina|Entity|false|false||Senna
null|Senna Plant|Entity|false|false||Sennanull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Constipation|Finding|false|false||constipationnull|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarinnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|nitroglycerin|Drug|false|false||Nitroglycerin
null|nitroglycerin|Drug|false|false||Nitroglycerinnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0741025;C2926613;C0008031;C1549543;C0030193|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025;C2926613;C0008031;C1549543;C0030193|chestnull|Administration Method - Pain|Finding|false|false|C1527391;C0817096|pain
null|Pain|Finding|false|false|C1527391;C0817096|painnull|null|Attribute|false|false||painnull|furosemide|Drug|false|false||Furosemide
null|furosemide|Drug|false|false||Furosemidenull|Daily|Time|false|false||DAILYnull|polyethylene glycols|Drug|false|false||Polyethylene Glycol
null|polyethylene glycols|Drug|false|false||Polyethylene Glycolnull|high-density polyethylene|Drug|false|false||Polyethylene
null|high-density polyethylene|Drug|false|false||Polyethylene
null|polyethylenes|Drug|false|false||Polyethylene
null|polyethylenes|Drug|false|false||Polyethylene
null|Polyethylene|Drug|false|false||Polyethylene
null|Polyethylene|Drug|false|false||Polyethylenenull|ethylene glycol|Drug|false|false||Glycol
null|Glycol|Drug|false|false||Glycol
null|ethylene glycol|Drug|false|false||Glycol
null|Glycols|Drug|false|false||Glycolnull|Daily|Time|false|false||DAILYnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|long-term care|Procedure|false|false||Extended Carenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|True primary (qualifier value)|Time|false|false||Primarynull|Primary|Modifier|false|false||Primarynull|Deep Vein Thrombosis|Disorder|false|false|C5239664;C0226514;C0042449|Deep vein thrombosis (DVT)null|Deep vein thrombosis of lower limb|Disorder|false|false|C0042449;C0226514|Deep vein thrombosis
null|Deep Vein Thrombosis|Disorder|false|false|C0042449;C0226514|Deep vein thrombosisnull|Structure of deep vein|Anatomy|false|false|C0149871;C0151950;C0042487;C0040053;C0149871;C0340708;C0149871|Deep veinnull|Deep Resection Margin|Attribute|false|false||Deepnull|Deep (qualifier value)|Modifier|false|false||Deepnull|Venous Thrombosis|Finding|false|false|C0226514;C0042449|vein thrombosisnull|Veins|Anatomy|false|false|C0149871;C0340708;C0149871;C0040053;C0149871;C0151950;C0042487|veinnull|Thrombosis|Finding|false|false|C0226514;C0042449|thrombosisnull|Deep Vein Thrombosis|Disorder|false|false|C0226514;C5239664;C0042449|DVT
null|Deep thrombophlebitis|Disorder|false|false|C0226514;C5239664;C0042449|DVTnull|area DVT|Anatomy|false|false|C0149871;C2926618;C0149871;C0151950|DVTnull|null|Attribute|false|false|C5239664|DVTnull|Neoplasm Metastasis|Disorder|false|false||Secondarynull|metastatic qualifier|Finding|false|false||Secondarynull|Secondary to|Modifier|false|false||Secondarynull|second (number)|LabModifier|false|false||Secondarynull|Upper gastrointestinal hemorrhage|Finding|false|false||Upper GI bleednull|Upper gastrointestinal tract series|Procedure|false|false||Upper GInull|Upper Surface|Modifier|false|false||Upper
null|Upper|Modifier|false|false||Uppernull|Gastrointestinal Hemorrhage|Finding|false|false||GI bleednull|Hemorrhage|Finding|false|false||bleednull|Left arm|Anatomy|false|false|C3495676;C1824218;C3715044;C1522541;C5400986;C4761640;C0018944|L armnull|Anorectal Malformations|Disorder|false|false|C5779993;C0446516;C1140618;C1269078|armnull|AKR1A1 wt Allele|Finding|false|false|C0446516;C1140618;C1269078;C5779993|arm
null|ARMC9 gene|Finding|false|false|C0446516;C1140618;C1269078;C5779993|armnull|Protocol Treatment Arm|Procedure|false|false|C0446516;C1140618;C1269078;C5779993|arm
null|Axillary Reverse Mapping|Procedure|false|false|C0446516;C1140618;C1269078;C5779993|arm
null|Study Arm|Procedure|false|false|C0446516;C1140618;C1269078;C5779993|armnull|Upper arm|Anatomy|false|false|C0018944;C1824218;C3715044;C1522541;C5400986;C4761640;C3495676|arm
null|null|Anatomy|false|false|C0018944;C1824218;C3715044;C1522541;C5400986;C4761640;C3495676|arm
null|Upper Extremity|Anatomy|false|false|C0018944;C1824218;C3715044;C1522541;C5400986;C4761640;C3495676|armnull|Hematoma|Finding|false|false|C0446516;C1140618;C1269078;C5779993|hematomanull|Superficial Thrombophlebitis|Disorder|false|false||Superficial thrombophlebitisnull|Superficial|Modifier|false|false||Superficialnull|Thrombophlebitis|Finding|false|false||thrombophlebitisnull|Antecubital Fossa|Anatomy|false|false||antecubital fossanull|Antecubital|Anatomy|false|false||antecubitalnull|Fossa|Anatomy|false|false||fossanull|Fossa <Euplerinae>|Entity|false|false||fossa
null|Cryptoprocta ferox|Entity|false|false||fossanull|Chronic Kidney Diseases|Disorder|false|false|C0227665;C0022646|Chronic kidney diseasenull|Chronic - Admission Level of Care Code|Finding|false|false||Chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||Chronicnull|chronic|Time|false|false||Chronicnull|Kidney Diseases|Disorder|false|false|C0227665;C0022646|kidney diseasenull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false|C0227665;C0022646|kidney
null|Benign neoplasm of kidney|Disorder|false|false|C0227665;C0022646|kidneynull|Kidney problem|Finding|false|false|C0227665;C0022646|kidneynull|examination of kidney|Procedure|false|false|C0227665;C0022646|kidney
null|Procedures on Kidney|Procedure|false|false|C0227665;C0022646|kidneynull|Kidney|Anatomy|false|false|C0012634;C0496927;C0496892;C0812426;C0022658;C1561643;C4554465;C0869841|kidney
null|Both kidneys|Anatomy|false|false|C0012634;C0496927;C0496892;C0812426;C0022658;C1561643;C4554465;C0869841|kidneynull|Disease|Disorder|false|false|C0227665;C0022646|diseasenull|Tumor stage|Attribute|false|false||Stagenull|Stage|Time|false|false||Stage
null|Phase|Time|false|false||Stagenull|Peripheral Vascular Diseases|Disorder|false|false|C0005847|Peripheral vascular diseasenull|Peripheral|Modifier|false|false||Peripheralnull|Vascular Diseases|Disorder|false|false|C0005847|vascular diseasenull|Blood Vessel|Anatomy|false|false|C0085096;C0012634;C0042373|vascularnull|Vascular|Modifier|false|false||vascularnull|Disease|Disorder|false|false|C0005847|diseasenull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Diabetes mellitus type IInull|Diabetes Mellitus|Disorder|false|false||Diabetes mellitusnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Diabetes
null|Diabetes|Disorder|false|false||Diabetes
null|Diabetes Mellitus|Disorder|false|false||Diabetesnull|Type - ParameterizedDataType|Finding|false|false||type
null|SGCG gene|Finding|false|false||typenull|null|Modifier|false|false||typenull|Coronary Artery Disease|Disorder|false|false|C0018787;C0205042;C0226004;C0003842|Coronary artery disease
null|Coronary Arteriosclerosis|Disorder|false|false|C0018787;C0205042;C0226004;C0003842|Coronary artery diseasenull|Coronary artery|Anatomy|false|false|C0012634;C1956346;C0010054;C0852949|Coronary arterynull|Heart|Anatomy|false|false|C1956346;C0010054|Coronarynull|Coronary|Modifier|false|false||Coronarynull|Arteriopathic disease|Disorder|false|false|C0226004;C0003842;C0205042|artery diseasenull|Arterial system|Anatomy|false|false|C0852949;C1956346;C0010054;C0012634|artery
null|Arteries|Anatomy|false|false|C0852949;C1956346;C0010054;C0012634|arterynull|Disease|Disorder|false|false|C0205042;C0226004;C0003842|diseasenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Disease|Disorder|false|false||Conditionnull|Logical Condition|Finding|false|false||Conditionnull|null|Attribute|false|false||Conditionnull|Condition|Modifier|false|false||Conditionnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Discharge instructions|Finding|false|false||Discharge Instructionsnull|hospital discharge instructions (treatment)|Procedure|false|false||Discharge Instructionsnull|null|Attribute|false|false||Discharge Instructionsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|FBXW7-AS1 gene|Finding|false|false||Dearnull|Production Class Code - Pleasure|Finding|false|false||pleasure
null|pleasurable emotion|Finding|false|false||pleasurenull|Pleasure - Animals raised for recreation|Entity|false|false||pleasurenull|Swelling of lower limb|Finding|false|false|C1140621;C0023216|leg swellingnull|Leg|Anatomy|false|false|C0581394;C1549543;C0030193;C0013604;C0038999|leg
null|Lower Extremity|Anatomy|false|false|C0581394;C1549543;C0030193;C0013604;C0038999|legnull|Swelling|Finding|false|false|C1140621;C0023216|swelling
null|Edema|Finding|false|false|C1140621;C0023216|swellingnull|Administration Method - Pain|Finding|false|false|C1140621;C0023216|pain
null|Pain|Finding|false|false|C1140621;C0023216|painnull|null|Attribute|false|false||painnull|Diagnostic tests|Procedure|false|false||Diagnostic testsnull|diagnostic tests device|Device|false|false||Diagnostic testsnull|Diagnostic agents|Drug|false|false||Diagnosticnull|Location Service Code - Diagnostic|Finding|false|false||Diagnostic
null|Diagnostic|Finding|false|false||Diagnosticnull|Diagnostic dental procedure|Procedure|false|false||Diagnostic
null|Diagnosis|Procedure|false|false||Diagnosticnull|Tests (qualifier value)|Finding|false|false||testsnull|Laboratory Procedures|Procedure|false|false||testsnull|Deep vein thrombosis of lower limb|Disorder|false|false|C0042449;C0226514|deep vein thrombosis
null|Deep Vein Thrombosis|Disorder|false|false|C0042449;C0226514|deep vein thrombosisnull|Structure of deep vein|Anatomy|false|false|C0149871;C0340708|deep veinnull|Deep Resection Margin|Attribute|false|false||deepnull|Deep (qualifier value)|Modifier|false|false||deepnull|Venous Thrombosis|Finding|false|false|C0042449|vein thrombosisnull|Veins|Anatomy|false|false|C0149871;C0340708;C0042487|veinnull|Thrombosis|Finding|false|false||thrombosisnull|Blood Clot|Finding|false|false||blood clots
null|Thrombus|Finding|false|false||blood clotsnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|In Blood|Finding|false|false||blood
null|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||bloodnull|Blood Clot|Finding|false|false||clotsnull|Leg|Anatomy|false|false|C5781420|legsnull|null|Attribute|false|false|C1140621|legsnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Thinning Weight Loss|Finding|false|false||thinningnull|Decreased thickness|Modifier|false|false||thinningnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|At home|Finding|false|false||at homenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Episode of|Time|false|false||episode ofnull|Episode of|Time|false|false||episodenull|Upper gastrointestinal hemorrhage|Finding|false|false||upper GI bleedingnull|Upper gastrointestinal tract series|Procedure|false|false||upper GInull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Gastrointestinal Hemorrhage|Finding|false|false||GI bleedingnull|Hemorrhage|Finding|false|false||bleedingnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Esophagogastroduodenoscopy|Procedure|false|false||EGDnull|Left upper arm structure|Anatomy|false|false|C1522541;C5400986;C4761640;C1824218;C3715044;C3495676|left arm
null|Left arm|Anatomy|false|false|C1522541;C5400986;C4761640;C1824218;C3715044;C3495676|left armnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Anorectal Malformations|Disorder|false|false|C0230347;C5779993;C0446516;C1140618;C1269078|armnull|AKR1A1 wt Allele|Finding|false|false|C0230347;C5779993;C0446516;C1140618;C1269078|arm
null|ARMC9 gene|Finding|false|false|C0230347;C5779993;C0446516;C1140618;C1269078|armnull|Protocol Treatment Arm|Procedure|false|false|C0446516;C1140618;C1269078;C0230347;C5779993|arm
null|Axillary Reverse Mapping|Procedure|false|false|C0446516;C1140618;C1269078;C0230347;C5779993|arm
null|Study Arm|Procedure|false|false|C0446516;C1140618;C1269078;C0230347;C5779993|armnull|Upper arm|Anatomy|false|false|C1522541;C5400986;C4761640;C1824218;C3715044;C3495676|arm
null|null|Anatomy|false|false|C1522541;C5400986;C4761640;C1824218;C3715044;C3495676|arm
null|Upper Extremity|Anatomy|false|false|C1522541;C5400986;C4761640;C1824218;C3715044;C3495676|armnull|Hematoma|Finding|false|false||hematomanull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Own|Finding|false|false||ownnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Blood Clot|Finding|false|false||blood clots
null|Thrombus|Finding|false|false||blood clotsnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Blood Clot|Finding|false|false||clotsnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Pharmaceutical Preparations|Drug|false|false||drug
null|Pharmacologic Substance|Drug|false|false||drugnull|Drug problem|Finding|false|false||drugnull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Upper gastrointestinal hemorrhage|Finding|false|false||upper GI bleednull|Upper gastrointestinal tract series|Procedure|false|false||upper GInull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Gastrointestinal Hemorrhage|Finding|false|false||GI bleednull|Hemorrhage|Finding|false|false||bleednull|pantoprazole|Drug|false|false||Pantoprazole
null|pantoprazole|Drug|false|false||Pantoprazolenull|Twice a day|Time|false|false||twice dailynull|Daily|Time|false|false||dailynull|Pharmaceutical Preparations|Drug|false|false||drug
null|Pharmacologic Substance|Drug|false|false||drugnull|Drug problem|Finding|false|false||drugnull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|week|Time|false|false||weeksnull|clopidogrel|Drug|false|false||Clopidogrel
null|clopidogrel|Drug|false|false||Clopidogrelnull|Plavix|Drug|false|false||Plavix
null|Plavix|Drug|false|false||Plavixnull|Cardiologists|Subject|false|false||cardiologistnull|Production Class Code - Pleasure|Finding|false|false||pleasure
null|pleasurable emotion|Finding|false|false||pleasurenull|Pleasure - Animals raised for recreation|Entity|false|false||pleasurenull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Hospital Stay|Time|false|false||hospital staynull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Care team|Finding|false|false||Care Teamnull|null|Attribute|false|false||Care Teamnull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|Team|Subject|false|false||Teamnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions