 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|42,51|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|42,51|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|42,56|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|76,85|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|76,85|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|76,90|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|132,135|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|143,150|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|143,150|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|152,160|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Drug|Indicator, Reagent, or Diagnostic Aid|Allergies|178,181|false|false|false|C0013343|Dyes|Dye
Event|Event|Allergies|178,181|false|false|false|||Dye
Drug|Biologically Active Substance|Allergies|183,189|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Drug|Element, Ion, or Isotope|Allergies|183,189|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Drug|Pharmacologic Substance|Allergies|183,189|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Event|Activity|Allergies|190,200|false|false|false|C2700400|Contain (action)|Containing
Finding|Functional Concept|Allergies|190,200|false|false|false|C0332256|Containing (qualifier value)|Containing
Drug|Indicator, Reagent, or Diagnostic Aid|Allergies|201,209|false|false|false|C0009924|Contrast Media|Contrast
Drug|Indicator, Reagent, or Diagnostic Aid|Allergies|201,215|false|false|false|C0009924|Contrast Media|Contrast Media
Anatomy|Tissue|Allergies|210,215|false|false|false|C0162867;C1254021|Media layer;Tunica Media|Media
Finding|Intellectual Product|Allergies|210,215|false|false|false|C0009458;C0677540|Communications Media;PAMS Media|Media
Drug|Organic Chemical|Allergies|218,227|false|false|false|C0030049|oxycodone|Oxycodone
Drug|Pharmacologic Substance|Allergies|218,227|false|false|false|C0030049|oxycodone|Oxycodone
Event|Event|Allergies|218,227|false|false|false|||Oxycodone
Procedure|Laboratory Procedure|Allergies|218,227|false|false|false|C0524222|Oxycodone measurement|Oxycodone
Drug|Organic Chemical|Allergies|231,241|false|false|false|C0055729|cilostazol|cilostazol
Drug|Pharmacologic Substance|Allergies|231,241|false|false|false|C0055729|cilostazol|cilostazol
Event|Event|Allergies|231,241|false|false|false|||cilostazol
Drug|Organic Chemical|Allergies|244,255|false|false|false|C1569608|varenicline|Varenicline
Drug|Pharmacologic Substance|Allergies|244,255|false|false|false|C1569608|varenicline|Varenicline
Event|Event|Allergies|244,255|false|false|false|||Varenicline
Event|Event|Allergies|258,267|false|false|false|||Attending
Finding|Functional Concept|Allergies|258,267|false|false|false|C1999232|Attending (action)|Attending
Event|Event|Chief Complaint|293,302|false|false|false|||Shortness
Attribute|Clinical Attribute|Chief Complaint|293,312|false|false|false|C2707305||Shortness of breath
Finding|Sign or Symptom|Chief Complaint|293,312|false|false|false|C0013404|Dyspnea|Shortness of breath
Finding|Body Substance|Chief Complaint|306,312|false|false|false|C0225386|Breath|breath
Finding|Classification|Chief Complaint|315,320|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|321,329|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|321,329|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|333,351|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|342,351|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|342,351|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|342,351|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|342,351|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|342,351|false|false|false|C0184661|Interventional procedure|Procedure
Disorder|Disease or Syndrome|History of Present Illness|414,418|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|History of Present Illness|414,418|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|History of Present Illness|414,418|false|false|false|||COPD
Finding|Gene or Genome|History of Present Illness|414,418|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|History of Present Illness|422,426|false|false|false|||home
Finding|Idea or Concept|History of Present Illness|422,426|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|History of Present Illness|422,426|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|History of Present Illness|422,426|false|false|false|C1553498|home health encounter|home
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|431,437|false|false|false|C0018792|Heart Atrium|atrial
Disorder|Disease or Syndrome|History of Present Illness|439,451|false|false|false|C0232197|Fibrillation|fibrillation
Event|Event|History of Present Illness|439,451|false|false|false|||fibrillation
Drug|Organic Chemical|History of Present Illness|455,463|false|false|false|C1831808|apixaban|apixaban
Drug|Pharmacologic Substance|History of Present Illness|455,463|false|false|false|C1831808|apixaban|apixaban
Event|Event|History of Present Illness|455,463|false|false|false|||apixaban
Disorder|Disease or Syndrome|History of Present Illness|465,477|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|History of Present Illness|465,477|false|false|false|||hypertension
Disorder|Disease or Syndrome|History of Present Illness|479,482|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|479,482|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|History of Present Illness|479,482|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|History of Present Illness|479,482|false|false|false|||CAD
Finding|Gene or Genome|History of Present Illness|479,482|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|History of Present Illness|479,482|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|History of Present Illness|479,482|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|479,482|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|History of Present Illness|488,502|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|hyperlipidemia
Event|Event|History of Present Illness|488,502|false|false|false|||hyperlipidemia
Finding|Finding|History of Present Illness|488,502|false|false|false|C0428465|Serum lipids high (finding)|hyperlipidemia
Event|Event|History of Present Illness|520,536|false|false|false|||hospitalizations
Procedure|Health Care Activity|History of Present Illness|520,536|false|false|false|C0019993|Hospitalization|hospitalizations
Disorder|Disease or Syndrome|History of Present Illness|541,545|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|History of Present Illness|541,545|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|History of Present Illness|541,545|false|false|false|||COPD
Finding|Gene or Genome|History of Present Illness|541,545|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|History of Present Illness|546,559|false|false|false|||exacerbations
Event|Event|History of Present Illness|566,575|false|false|false|||presented
Event|Event|History of Present Illness|581,588|false|false|false|||dyspnea
Finding|Finding|History of Present Illness|581,588|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|History of Present Illness|581,588|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Event|Event|History of Present Illness|620,630|false|false|false|||admissions
Procedure|Health Care Activity|History of Present Illness|620,630|false|false|false|C0184666|Hospital admission|admissions
Event|Event|History of Present Illness|635,642|false|false|false|||dyspnea
Finding|Finding|History of Present Illness|635,642|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|History of Present Illness|635,642|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Event|Event|History of Present Illness|662,672|false|false|false|||discharged
Finding|Idea or Concept|History of Present Illness|688,691|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|History of Present Illness|688,691|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|History of Present Illness|692,701|false|false|false|||inpatient
Finding|Idea or Concept|History of Present Illness|692,701|false|false|false|C1548438;C1549404|Patient Class - Inpatient;Referral category - Inpatient|inpatient
Procedure|Health Care Activity|History of Present Illness|692,701|false|false|false|C1555324|inpatient encounter|inpatient
Event|Event|History of Present Illness|702,711|false|false|false|||admission
Procedure|Health Care Activity|History of Present Illness|702,711|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Disorder|Disease or Syndrome|History of Present Illness|717,721|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|History of Present Illness|717,721|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|History of Present Illness|717,721|false|false|false|||COPD
Finding|Gene or Genome|History of Present Illness|717,721|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|History of Present Illness|717,734|false|false|false|C0740304|COPD exacerbation|COPD exacerbation
Event|Event|History of Present Illness|722,734|false|false|false|||exacerbation
Finding|Finding|History of Present Illness|722,734|false|false|false|C4086268|Exacerbation|exacerbation
Event|Event|History of Present Illness|744,754|false|false|false|||discharged
Finding|Finding|History of Present Illness|758,766|false|false|false|C0231448;C5781021|Extended (finding);Extension|extended
Finding|Functional Concept|History of Present Illness|758,766|false|false|false|C0231448;C5781021|Extended (finding);Extension|extended
Drug|Hormone|History of Present Illness|767,777|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|History of Present Illness|767,777|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|History of Present Illness|767,777|false|false|false|C0032952|prednisone|prednisone
Event|Event|History of Present Illness|767,777|false|false|false|||prednisone
Event|Event|History of Present Illness|779,784|false|false|false|||taper
Procedure|Health Care Activity|History of Present Illness|779,784|false|false|false|C0441640||taper
Disorder|Disease or Syndrome|History of Present Illness|790,794|false|false|false|C0270724|Infantile Neuroaxonal Dystrophy|plan
Event|Event|History of Present Illness|790,794|false|false|false|||plan
Finding|Functional Concept|History of Present Illness|790,794|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Intellectual Product|History of Present Illness|790,794|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Mental Process|History of Present Illness|790,794|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Drug|Hormone|History of Present Illness|807,817|false|false|false|C0032952|prednisone|Prednisone
Drug|Organic Chemical|History of Present Illness|807,817|false|false|false|C0032952|prednisone|Prednisone
Drug|Pharmacologic Substance|History of Present Illness|807,817|false|false|false|C0032952|prednisone|Prednisone
Finding|Functional Concept|History of Present Illness|822,828|false|false|false|C1706059|Finish - dosing instruction imperative|finish
Event|Event|History of Present Illness|851,856|false|false|false|||taper
Procedure|Health Care Activity|History of Present Illness|851,856|false|false|false|C0441640||taper
Finding|Idea or Concept|History of Present Illness|897,900|false|false|false|C1548556|Etc.|etc
Event|Event|History of Present Illness|932,944|false|false|false|||presentation
Finding|Idea or Concept|History of Present Illness|932,944|false|false|false|C0449450|Presentation|presentation
Finding|Body Substance|History of Present Illness|946,953|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|946,953|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|946,953|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|977,986|false|false|false|||shortness
Attribute|Clinical Attribute|History of Present Illness|977,996|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|History of Present Illness|977,996|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|History of Present Illness|990,996|false|false|false|C0225386|Breath|breath
Drug|Organic Chemical|History of Present Illness|1012,1017|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|1012,1017|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|History of Present Illness|1012,1017|false|false|false|||cough
Finding|Sign or Symptom|History of Present Illness|1012,1017|false|false|false|C0010200|Coughing|cough
Event|Event|History of Present Illness|1022,1030|false|false|false|||wheezing
Finding|Sign or Symptom|History of Present Illness|1022,1030|false|false|false|C0043144|Wheezing|wheezing
Disorder|Disease or Syndrome|History of Present Illness|1042,1046|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|History of Present Illness|1042,1046|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|History of Present Illness|1042,1046|false|false|false|||COPD
Finding|Gene or Genome|History of Present Illness|1042,1046|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|History of Present Illness|1047,1060|false|false|false|||exacerbations
Event|Event|History of Present Illness|1066,1074|true|false|false|||reported
Event|Event|History of Present Illness|1082,1090|true|false|false|||inhalers
Event|Event|History of Present Illness|1095,1103|true|false|false|||directed
Drug|Organic Chemical|History of Present Illness|1113,1119|true|false|false|C0723011|Relief brand of phenylephrine|relief
Drug|Pharmacologic Substance|History of Present Illness|1113,1119|true|false|false|C0723011|Relief brand of phenylephrine|relief
Event|Event|History of Present Illness|1113,1119|true|false|false|||relief
Finding|Finding|History of Present Illness|1113,1119|true|false|false|C0564405|Feeling relief|relief
Finding|Body Substance|History of Present Illness|1125,1132|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1125,1132|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1125,1132|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|1133,1141|false|false|false|||reported
Event|Event|History of Present Illness|1163,1172|false|false|false|||identical
Event|Event|History of Present Illness|1185,1197|false|false|false|||presentation
Finding|Idea or Concept|History of Present Illness|1185,1197|false|false|false|C0449450|Presentation|presentation
Event|Event|History of Present Illness|1208,1212|false|false|false|||felt
Event|Event|History of Present Illness|1227,1233|true|false|false|||taking
Attribute|Clinical Attribute|History of Present Illness|1243,1254|true|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|History of Present Illness|1243,1254|true|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|History of Present Illness|1243,1254|true|false|false|||medications
Finding|Intellectual Product|History of Present Illness|1243,1254|true|false|false|C4284232|Medications|medications
Event|Event|History of Present Illness|1268,1272|true|false|false|||wish
Event|Event|History of Present Illness|1277,1285|true|false|false|||continue
Event|Event|History of Present Illness|1289,1293|true|false|false|||take
Drug|Hormone|History of Present Illness|1294,1304|true|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|History of Present Illness|1294,1304|true|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|History of Present Illness|1294,1304|true|false|false|C0032952|prednisone|prednisone
Event|Event|History of Present Illness|1294,1304|true|false|false|||prednisone
Finding|Body Substance|History of Present Illness|1310,1317|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1310,1317|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1310,1317|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|1327,1332|false|false|false|||noted
Event|Event|History of Present Illness|1342,1351|false|false|false|||increased
Event|Event|History of Present Illness|1355,1366|false|false|false|||requirement
Finding|Functional Concept|History of Present Illness|1355,1366|false|false|false|C1514873|Requirement|requirement
Event|Event|History of Present Illness|1379,1387|false|false|false|||referred
Event|Event|History of Present Illness|1415,1425|false|false|false|||management
Event|Occupational Activity|History of Present Illness|1415,1425|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|History of Present Illness|1415,1425|false|false|false|C0376636|Disease Management|management
Event|Event|History of Present Illness|1443,1446|false|false|false|||see
Procedure|Health Care Activity|History of Present Illness|1453,1462|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|History of Present Illness|1463,1467|false|false|false|||note
Event|Event|History of Present Illness|1473,1480|false|false|false|||details
Event|Event|History of Present Illness|1497,1506|false|false|false|||admission
Procedure|Health Care Activity|History of Present Illness|1497,1506|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Idea or Concept|History of Present Illness|1523,1530|false|false|false|C1555582|Initial (abbreviation)|initial
Drug|Food|History of Present Illness|1531,1536|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|vital
Attribute|Clinical Attribute|History of Present Illness|1531,1542|false|false|false|C0488614;C0518766|Vital signs|vital signs
Procedure|Health Care Activity|History of Present Illness|1531,1542|false|false|false|C0150404|Taking vital signs|vital signs
Event|Event|History of Present Illness|1537,1542|false|false|false|||signs
Finding|Finding|History of Present Illness|1537,1542|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|History of Present Illness|1537,1542|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Lab|Laboratory or Test Result|History of Present Illness|1571,1575|false|false|false|C0587081|Laboratory test finding|Labs
Event|Event|History of Present Illness|1582,1589|false|false|false|||notable
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1601,1604|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Hormone|History of Present Illness|1601,1604|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Pharmacologic Substance|History of Present Illness|1601,1604|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Event|Event|History of Present Illness|1601,1604|false|false|false|||BNP
Finding|Gene or Genome|History of Present Illness|1601,1604|false|false|false|C1417808;C2982014|NPPB gene;NPPB wt Allele|BNP
Procedure|Laboratory Procedure|History of Present Illness|1601,1604|false|false|false|C1095989|Brain natriuretic peptide measurement|BNP
Drug|Biologically Active Substance|History of Present Illness|1611,1621|false|false|false|C0010294|creatinine|creatinine
Drug|Organic Chemical|History of Present Illness|1611,1621|false|false|false|C0010294|creatinine|creatinine
Event|Event|History of Present Illness|1611,1621|false|false|false|||creatinine
Finding|Physiologic Function|History of Present Illness|1611,1621|false|false|false|C4551889|Creatinine metabolic function|creatinine
Procedure|Laboratory Procedure|History of Present Illness|1611,1621|false|false|false|C0201975|Creatinine measurement|creatinine
Finding|Body Substance|History of Present Illness|1630,1637|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|1630,1637|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|1630,1637|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Antibiotic|History of Present Illness|1649,1661|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|History of Present Illness|1649,1661|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|History of Present Illness|1649,1661|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Event|Event|History of Present Illness|1649,1661|false|false|false|||azithromycin
Drug|Organic Chemical|History of Present Illness|1666,1672|false|false|false|C0939692|DuoNeb|duoneb
Drug|Pharmacologic Substance|History of Present Illness|1666,1672|false|false|false|C0939692|DuoNeb|duoneb
Event|Event|History of Present Illness|1666,1672|false|false|false|||duoneb
Finding|Body Substance|History of Present Illness|1674,1681|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|1674,1681|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|1674,1681|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|History of Present Illness|1686,1695|false|false|false|||scheduled
Event|Event|History of Present Illness|1736,1748|true|false|false|||administered
Event|Activity|History of Present Illness|1755,1762|true|false|false|C1706079||arrival
Event|Event|History of Present Illness|1755,1762|true|false|false|||arrival
Finding|Functional Concept|History of Present Illness|1755,1762|true|false|false|C1555577|arrival - ActRelationshipType|arrival
Anatomy|Anatomical Structure|History of Present Illness|1771,1776|false|false|false|C3714591|Floor (anatomic)|floor
Event|Activity|History of Present Illness|1786,1793|false|false|false|C1706079||arrival
Event|Event|History of Present Illness|1786,1793|false|false|false|||arrival
Finding|Functional Concept|History of Present Illness|1786,1793|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Anatomy|Anatomical Structure|History of Present Illness|1801,1806|false|false|false|C3714591|Floor (anatomic)|floor
Event|Event|History of Present Illness|1812,1822|false|false|false|||complained
Event|Event|History of Present Illness|1826,1834|false|false|false|||wheezing
Finding|Sign or Symptom|History of Present Illness|1826,1834|false|false|false|C0043144|Wheezing|wheezing
Event|Event|History of Present Illness|1839,1842|false|false|false|||SOB
Finding|Sign or Symptom|History of Present Illness|1839,1842|false|false|false|C0013404|Dyspnea|SOB
Event|Event|History of Present Illness|1859,1863|false|false|false|||felt
Finding|Finding|History of Present Illness|1864,1868|false|false|false|C5575035|Well (answer to question)|well
Event|Event|History of Present Illness|1874,1880|false|false|false|||agreed
Event|Event|History of Present Illness|1893,1908|false|false|false|||methyprednisone
Event|Event|History of Present Illness|1923,1927|true|false|false|||wish
Drug|Hormone|History of Present Illness|1936,1946|true|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|History of Present Illness|1936,1946|true|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|History of Present Illness|1936,1946|true|false|false|C0032952|prednisone|prednisone
Event|Event|History of Present Illness|1936,1946|true|false|false|||prednisone
Event|Event|History of Present Illness|1961,1967|false|false|false|||REVIEW
Finding|Idea or Concept|History of Present Illness|1961,1967|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|REVIEW
Finding|Intellectual Product|History of Present Illness|1961,1967|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|REVIEW
Finding|Functional Concept|History of Present Illness|1961,1970|false|false|false|C0699752|Review of|REVIEW OF
Attribute|Clinical Attribute|History of Present Illness|1961,1978|false|false|false|C0488564;C0488565||REVIEW OF SYSTEMS
Procedure|Health Care Activity|History of Present Illness|1961,1978|false|false|false|C0489633|Review of systems (procedure)|REVIEW OF SYSTEMS
Event|Event|History of Present Illness|1971,1978|false|false|false|||SYSTEMS
Finding|Functional Concept|History of Present Illness|1971,1978|false|false|false|C0449913|System|SYSTEMS
Disorder|Disease or Syndrome|History of Present Illness|1984,1987|false|false|false|C0268529|Proline dehydrogenase deficiency|HPI
Event|Event|History of Present Illness|1984,1987|false|false|false|||HPI
Finding|Finding|History of Present Illness|1984,1987|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Finding|Molecular Function|History of Present Illness|1984,1987|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Event|Event|History of Present Illness|1989,1995|false|false|false|||Denies
Event|Event|History of Present Illness|1996,2004|true|false|false|||headache
Finding|Sign or Symptom|History of Present Illness|1996,2004|true|false|false|C0018681|Headache|headache
Finding|Functional Concept|History of Present Illness|2006,2012|true|false|false|C0234621|Visual|visual
Finding|Finding|History of Present Illness|2006,2020|true|false|false|C0750280|Visual changes|visual changes
Event|Event|History of Present Illness|2013,2020|true|false|false|||changes
Finding|Functional Concept|History of Present Illness|2013,2020|true|false|false|C0392747|Changing|changes
Disorder|Disease or Syndrome|History of Present Illness|2023,2034|true|false|false|C0031350|Pharyngitis|pharyngitis
Event|Event|History of Present Illness|2023,2034|true|false|false|||pharyngitis
Event|Event|History of Present Illness|2036,2042|false|false|false|||fevers
Finding|Sign or Symptom|History of Present Illness|2036,2042|false|false|false|C0015967|Fever|fevers
Event|Event|History of Present Illness|2044,2050|false|false|false|||chills
Finding|Sign or Symptom|History of Present Illness|2044,2050|false|false|false|C0085593|Chills|chills
Event|Event|History of Present Illness|2052,2058|false|false|false|||sweats
Finding|Body Substance|History of Present Illness|2052,2058|false|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Finding|Finding|History of Present Illness|2052,2058|false|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Attribute|Clinical Attribute|History of Present Illness|2060,2066|false|false|false|C0944911||weight
Event|Event|History of Present Illness|2060,2066|false|false|false|||weight
Finding|Finding|History of Present Illness|2060,2066|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|History of Present Illness|2060,2066|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|History of Present Illness|2060,2066|false|false|false|C1305866|Weighing patient|weight
Finding|Finding|History of Present Illness|2060,2071|false|false|false|C1262477;C3540682|Losing Weight (question);Weight Loss|weight loss
Finding|Intellectual Product|History of Present Illness|2060,2071|false|false|false|C1262477;C3540682|Losing Weight (question);Weight Loss|weight loss
Event|Event|History of Present Illness|2067,2071|false|false|false|||loss
Finding|Finding|History of Present Illness|2067,2071|false|false|false|C5890125|Loss (adaptation)|loss
Anatomy|Body Location or Region|History of Present Illness|2073,2078|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|2073,2078|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|2073,2083|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|2073,2083|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|2079,2083|false|true|false|C2598155||pain
Event|Event|History of Present Illness|2079,2083|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|2079,2083|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|2079,2083|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Location or Region|History of Present Illness|2086,2095|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|History of Present Illness|2086,2100|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|History of Present Illness|2096,2100|false|false|false|C2598155||pain
Event|Event|History of Present Illness|2096,2100|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|2096,2100|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|2096,2100|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|History of Present Illness|2102,2108|false|false|false|C4255480||nausea
Event|Event|History of Present Illness|2102,2108|false|false|false|||nausea
Finding|Sign or Symptom|History of Present Illness|2102,2108|false|false|false|C0027497|Nausea|nausea
Event|Event|History of Present Illness|2110,2118|false|false|false|||vomiting
Finding|Sign or Symptom|History of Present Illness|2110,2118|false|false|false|C0042963|Vomiting|vomiting
Event|Event|History of Present Illness|2120,2128|false|false|false|||diarrhea
Finding|Finding|History of Present Illness|2120,2128|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|History of Present Illness|2120,2128|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Event|Event|History of Present Illness|2130,2142|false|false|false|||constipation
Finding|Sign or Symptom|History of Present Illness|2130,2142|false|false|false|C0009806|Constipation|constipation
Disorder|Disease or Syndrome|History of Present Illness|2145,2157|false|false|false|C0018932|Hematochezia|hematochezia
Event|Event|History of Present Illness|2145,2157|false|false|false|||hematochezia
Finding|Sign or Symptom|History of Present Illness|2145,2157|false|false|false|C1321898|Blood in stool|hematochezia
Event|Event|History of Present Illness|2159,2166|false|false|false|||dysuria
Finding|Sign or Symptom|History of Present Illness|2159,2166|false|false|false|C0013428|Dysuria|dysuria
Disorder|Disease or Syndrome|History of Present Illness|2168,2172|false|false|false|C5779629|Eruption of skin (disorder)|rash
Event|Event|History of Present Illness|2168,2172|false|false|false|||rash
Finding|Pathologic Function|History of Present Illness|2168,2172|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|History of Present Illness|2168,2172|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Disorder|Disease or Syndrome|History of Present Illness|2174,2186|false|false|false|C0030554|Paresthesia|paresthesias
Event|Event|History of Present Illness|2174,2186|false|false|false|||paresthesias
Event|Event|History of Present Illness|2192,2200|false|false|false|||weakness
Finding|Sign or Symptom|History of Present Illness|2192,2200|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Disorder|Disease or Syndrome|Past Medical History|2228,2232|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Past Medical History|2228,2232|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Past Medical History|2228,2232|false|false|false|||COPD
Finding|Gene or Genome|Past Medical History|2228,2232|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|Past Medical History|2233,2239|false|false|false|C0004096|Asthma|Asthma
Event|Event|Past Medical History|2233,2239|false|false|false|||Asthma
Event|Event|Past Medical History|2243,2247|false|false|false|||home
Finding|Idea or Concept|Past Medical History|2243,2247|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Past Medical History|2243,2247|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Past Medical History|2243,2247|false|false|false|C1553498|home health encounter|home
Finding|Finding|Past Medical History|2256,2264|false|false|false|C0741302|atypia morphology|Atypical
Finding|Sign or Symptom|Past Medical History|2256,2275|false|false|false|C0262384|Atypical chest pain|Atypical Chest Pain
Anatomy|Body Location or Region|Past Medical History|2265,2270|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|Past Medical History|2265,2270|false|false|false|C0741025|Chest problem|Chest
Attribute|Clinical Attribute|Past Medical History|2265,2275|false|false|false|C2926613||Chest Pain
Finding|Sign or Symptom|Past Medical History|2265,2275|false|false|false|C0008031|Chest Pain|Chest Pain
Attribute|Clinical Attribute|Past Medical History|2271,2275|false|true|false|C2598155||Pain
Event|Event|Past Medical History|2271,2275|false|false|false|||Pain
Finding|Functional Concept|Past Medical History|2271,2275|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Past Medical History|2271,2275|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Disorder|Disease or Syndrome|Past Medical History|2278,2290|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|Past Medical History|2278,2290|false|false|false|||Hypertension
Disorder|Disease or Syndrome|Past Medical History|2293,2307|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|Hyperlipidemia
Event|Event|Past Medical History|2293,2307|false|false|false|||Hyperlipidemia
Finding|Finding|Past Medical History|2293,2307|false|false|false|C0428465|Serum lipids high (finding)|Hyperlipidemia
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2328,2334|false|false|false|C0018792|Heart Atrium|Atrial
Attribute|Clinical Attribute|Past Medical History|2328,2347|false|false|false|C2926591||Atrial Fibrillation
Disorder|Disease or Syndrome|Past Medical History|2328,2347|false|false|false|C0004238|Atrial Fibrillation|Atrial Fibrillation
Lab|Laboratory or Test Result|Past Medical History|2328,2347|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Atrial Fibrillation
Disorder|Disease or Syndrome|Past Medical History|2335,2347|false|false|false|C0232197|Fibrillation|Fibrillation
Event|Event|Past Medical History|2335,2347|false|false|false|||Fibrillation
Drug|Organic Chemical|Past Medical History|2351,2359|false|false|false|C1831808|apixaban|Apixaban
Drug|Pharmacologic Substance|Past Medical History|2351,2359|false|false|false|C1831808|apixaban|Apixaban
Disorder|Mental or Behavioral Dysfunction|Past Medical History|2362,2369|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|Anxiety
Event|Event|Past Medical History|2362,2369|false|false|false|||Anxiety
Finding|Sign or Symptom|Past Medical History|2362,2369|false|false|false|C0860603|Anxiety symptoms|Anxiety
Anatomy|Body Location or Region|Past Medical History|2372,2380|false|false|false|C0027530|Neck|Cervical
Disorder|Disease or Syndrome|Past Medical History|2372,2392|false|false|false|C0263884|Cervical radiculitis|Cervical Radiculitis
Disorder|Disease or Syndrome|Past Medical History|2381,2392|false|false|false|C0034544|Radiculitis|Radiculitis
Event|Event|Past Medical History|2381,2392|false|false|false|||Radiculitis
Anatomy|Body Location or Region|Past Medical History|2395,2403|false|false|false|C0027530|Neck|Cervical
Disorder|Disease or Syndrome|Past Medical History|2395,2415|false|false|false|C0158241;C1384641|Cervical spondylosis;Cervical spondylosis without myelopathy|Cervical Spondylosis
Disorder|Disease or Syndrome|Past Medical History|2404,2415|false|false|false|C0038019|Spondylosis|Spondylosis
Event|Event|Past Medical History|2404,2415|false|false|false|||Spondylosis
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2418,2426|false|false|false|C0018787|Heart|Coronary
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2418,2433|false|false|false|C0205042|Coronary artery|Coronary Artery
Disorder|Disease or Syndrome|Past Medical History|2418,2441|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|Coronary Artery Disease
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2427,2433|false|false|false|C0003842;C0226004|Arterial system;Arteries|Artery
Anatomy|Body System|Past Medical History|2427,2433|false|false|false|C0003842;C0226004|Arterial system;Arteries|Artery
Disorder|Disease or Syndrome|Past Medical History|2427,2441|false|false|false|C0852949|Arteriopathic disease|Artery Disease
Disorder|Disease or Syndrome|Past Medical History|2434,2441|false|false|false|C0012634|Disease|Disease
Event|Event|Past Medical History|2434,2441|false|false|false|||Disease
Finding|Sign or Symptom|Past Medical History|2444,2452|false|false|false|C0018681|Headache|Headache
Disorder|Disease or Syndrome|Past Medical History|2455,2461|false|false|false|C0019340;C0854331|Herpes simplex dermatitis|Herpes
Disorder|Disease or Syndrome|Past Medical History|2455,2468|false|false|false|C0019360;C0042338|Herpes zoster (disorder);herpesvirus 3, human|Herpes Zoster
Disorder|Virus|Past Medical History|2455,2468|false|false|false|C0019360;C0042338|Herpes zoster (disorder);herpesvirus 3, human|Herpes Zoster
Disorder|Disease or Syndrome|Past Medical History|2462,2468|false|false|false|C0019360|Herpes zoster (disorder)|Zoster
Event|Event|Past Medical History|2462,2468|false|false|false|||Zoster
Finding|Pathologic Function|Past Medical History|2471,2482|false|false|false|C0017181|Gastrointestinal Hemorrhage|GI Bleeding
Event|Event|Past Medical History|2474,2482|false|false|false|||Bleeding
Finding|Pathologic Function|Past Medical History|2474,2482|false|false|false|C0019080|Hemorrhage|Bleeding
Disorder|Disease or Syndrome|Past Medical History|2485,2512|false|false|false|C0085096|Peripheral Vascular Diseases|Peripheral Vascular Disease
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2496,2504|false|false|false|C0005847|Blood Vessel|Vascular
Disorder|Disease or Syndrome|Past Medical History|2496,2512|false|false|false|C0042373|Vascular Diseases|Vascular Disease
Disorder|Disease or Syndrome|Past Medical History|2505,2512|false|false|false|C0012634|Disease|Disease
Event|Event|Past Medical History|2505,2512|false|false|false|||Disease
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2527,2532|false|false|false|C0020889|Bone structure of ilium|iliac
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2527,2539|false|false|false|C0850459|iliac stents|iliac stents
Event|Event|Past Medical History|2533,2539|false|false|false|||stents
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2546,2549|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|Past Medical History|2546,2549|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|Past Medical History|2546,2549|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|Past Medical History|2546,2549|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|Past Medical History|2546,2549|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2546,2549|false|false|false|C1292890|Procedure on hip|hip
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2546,2561|false|false|false|C0392806|Prosthetic arthroplasty of hip (procedure)|hip replacement
Event|Event|Past Medical History|2550,2561|false|false|false|||replacement
Finding|Functional Concept|Past Medical History|2550,2561|false|false|false|C0559956|Replacement|replacement
Procedure|Health Care Activity|Past Medical History|2550,2561|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2550,2561|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Event|Event|Family Medical History|2600,2606|false|false|false|||Mother
Finding|Idea or Concept|Family Medical History|2600,2606|false|false|false|C1546508|Relationship - Mother|Mother
Disorder|Disease or Syndrome|Family Medical History|2612,2618|false|false|false|C0004096|Asthma|asthma
Event|Event|Family Medical History|2612,2618|false|false|false|||asthma
Disorder|Disease or Syndrome|Family Medical History|2623,2635|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|Family Medical History|2623,2635|false|false|false|||hypertension
Finding|Conceptual Entity|Family Medical History|2637,2643|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|Family Medical History|2637,2643|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2649,2654|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|Family Medical History|2649,2654|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|Family Medical History|2649,2654|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Finding|Finding|Family Medical History|2649,2654|false|false|false|C0750873|COLON PROBLEM|colon
Disorder|Neoplastic Process|Family Medical History|2649,2661|false|false|false|C0007102;C0346629;C0699790|Colon Carcinoma;Malignant neoplasm of large intestine;Malignant tumor of colon|colon cancer
Disorder|Neoplastic Process|Family Medical History|2655,2661|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Family Medical History|2655,2661|false|false|false|||cancer
Event|Event|Family Medical History|2664,2671|false|false|false|||Brother
Finding|Conceptual Entity|Family Medical History|2664,2671|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Idea or Concept|Family Medical History|2664,2671|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Disorder|Neoplastic Process|Family Medical History|2677,2685|false|false|false|C0023418|leukemia|leukemia
Event|Event|Family Medical History|2677,2685|false|false|false|||leukemia
Finding|Finding|General Exam|2705,2713|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|General Exam|2705,2713|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|General Exam|2705,2713|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|General Exam|2705,2725|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAMINATION
Procedure|Health Care Activity|General Exam|2705,2725|false|false|false|C0031809|Physical Examination|PHYSICAL EXAMINATION
Event|Activity|General Exam|2714,2725|false|false|false|C4321457|Examination|EXAMINATION
Event|Event|General Exam|2714,2725|false|false|false|||EXAMINATION
Procedure|Health Care Activity|General Exam|2714,2725|false|false|false|C0031809;C0582103|Medical Examination;Physical Examination|EXAMINATION
Procedure|Health Care Activity|General Exam|2729,2738|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|General Exam|2776,2782|false|false|false|||VITALS
Event|Event|General Exam|2817,2824|false|false|false|||GENERAL
Finding|Classification|General Exam|2817,2824|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|General Exam|2817,2824|false|false|false|C3812897|General medical service|GENERAL
Event|Event|General Exam|2826,2834|true|false|false|||Pleasant
Finding|Mental Process|General Exam|2826,2834|true|false|false|C2987187|Pleasant|Pleasant
Finding|Finding|General Exam|2836,2840|true|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|2841,2850|true|false|false|||appearing
Finding|Idea or Concept|General Exam|2858,2866|true|false|false|C0750489|apparent|apparent
Event|Event|General Exam|2867,2875|true|false|false|||distress
Finding|Finding|General Exam|2867,2875|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|General Exam|2867,2875|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|General Exam|2880,2885|false|false|false|C1512338|HEENT|HEENT
Event|Event|General Exam|2887,2900|true|false|false|||Normocephalic
Event|Event|General Exam|2902,2912|true|false|false|||atraumatic
Anatomy|Body Part, Organ, or Organ Component|General Exam|2917,2929|true|false|false|C0009758|conjunctiva|conjunctival
Finding|Functional Concept|General Exam|2917,2929|true|false|false|C1522483|Conjunctival Route of Administration|conjunctival
Finding|Finding|General Exam|2917,2936|true|false|false|C2071267|Conjunctival pallor|conjunctival pallor
Event|Event|General Exam|2930,2936|true|false|false|||pallor
Finding|Finding|General Exam|2930,2936|true|false|false|C0241137|Pallor of skin|pallor
Anatomy|Body Part, Organ, or Organ Component|General Exam|2941,2948|true|false|false|C0036410|Sclera|scleral
Finding|Finding|General Exam|2941,2956|true|false|false|C0240962|Scleral icterus|scleral icterus
Finding|Sign or Symptom|General Exam|2949,2956|true|false|false|C0022346|Icterus|icterus
Event|Event|General Exam|2958,2964|false|false|false|||PERRLA
Finding|Finding|General Exam|2958,2964|false|false|false|C2143306|PERRLA|PERRLA
Event|Event|General Exam|2966,2970|false|false|false|||EOMI
Event|Event|General Exam|2975,2980|false|false|false|||clear
Finding|Idea or Concept|General Exam|2975,2980|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Location or Region|General Exam|2985,2989|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|General Exam|2985,2989|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|General Exam|2985,2989|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|General Exam|2991,2997|true|false|false|||Supple
Finding|Functional Concept|General Exam|2991,2997|true|false|false|C0332254|Supple|Supple
Anatomy|Body Part, Organ, or Organ Component|General Exam|3002,3005|true|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|General Exam|3002,3005|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|General Exam|3002,3005|true|false|false|||LAD
Finding|Gene or Genome|General Exam|3002,3005|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Disorder|Disease or Syndrome|General Exam|3010,3021|true|false|false|C0018021|Goiter|thyromegaly
Event|Event|General Exam|3010,3021|true|false|false|||thyromegaly
Event|Event|General Exam|3023,3026|true|false|false|||JVP
Finding|Finding|General Exam|3023,3026|true|false|false|C0428897|Jugular venous pressure|JVP
Anatomy|Body Part, Organ, or Organ Component|General Exam|3036,3043|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|General Exam|3036,3043|false|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Event|General Exam|3062,3069|true|false|false|||murmurs
Finding|Finding|General Exam|3062,3069|true|false|false|C0018808|Heart murmur|murmurs
Event|Event|General Exam|3070,3074|true|false|false|||rubs
Finding|Finding|General Exam|3070,3074|true|false|false|C0232267|Pericardial friction rub|rubs
Event|Event|General Exam|3078,3085|true|false|false|||gallops
Anatomy|Body Part, Organ, or Organ Component|General Exam|3090,3099|false|false|false|C0024109|Lung|PULMONARY
Attribute|Clinical Attribute|General Exam|3090,3099|false|false|false|C2707265||PULMONARY
Finding|Finding|General Exam|3090,3099|false|false|false|C4522268|Pulmonary (intended site)|PULMONARY
Finding|Intellectual Product|General Exam|3101,3105|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Finding|Organism Function|General Exam|3106,3116|false|false|false|C0231800|Expiration, Respiratory|expiratory
Finding|Sign or Symptom|General Exam|3106,3124|false|false|false|C0231875|Expiratory wheezing|expiratory wheezes
Event|Event|General Exam|3117,3124|false|false|false|||wheezes
Finding|Sign or Symptom|General Exam|3117,3124|false|false|false|C0043144|Wheezing|wheezes
Anatomy|Body Location or Region|General Exam|3132,3136|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|General Exam|3132,3136|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|General Exam|3132,3136|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|General Exam|3132,3136|false|false|false|C0740941|Lung Problem|lung
Event|Event|General Exam|3137,3143|false|false|false|||fields
Anatomy|Body Location or Region|General Exam|3147,3154|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|General Exam|3147,3154|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|General Exam|3147,3154|false|false|false|||ABDOMEN
Finding|Finding|General Exam|3147,3154|false|false|false|C0941288|Abdomen problem|ABDOMEN
Anatomy|Body Part, Organ, or Organ Component|General Exam|3163,3168|false|false|false|C0021853|Intestines|bowel
Finding|Finding|General Exam|3163,3175|false|false|false|C0232693|Bowel sounds|bowel sounds
Event|Event|General Exam|3169,3175|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|General Exam|3169,3175|false|false|false|C0037709||sounds
Disorder|Disease or Syndrome|General Exam|3177,3181|true|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|General Exam|3177,3181|true|false|false|||soft
Event|Event|General Exam|3214,3226|true|false|false|||organomegaly
Finding|Finding|General Exam|3214,3226|true|false|false|C4054315|Organomegaly|organomegaly
Anatomy|Body Part, Organ, or Organ Component|General Exam|3231,3242|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Event|Event|General Exam|3244,3248|true|false|false|||Warm
Finding|Finding|General Exam|3244,3248|true|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|3244,3248|true|false|false|C0687712|warming process|Warm
Finding|Finding|General Exam|3250,3254|true|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|3255,3263|true|false|false|||perfused
Event|Event|General Exam|3268,3276|true|false|false|||cyanosis
Finding|Sign or Symptom|General Exam|3268,3276|true|false|false|C0010520|Cyanosis|cyanosis
Disorder|Anatomical Abnormality|General Exam|3278,3286|true|false|false|C0149651|Clubbing|clubbing
Event|Event|General Exam|3278,3286|true|false|false|||clubbing
Attribute|Clinical Attribute|General Exam|3291,3296|true|false|false|C1717255||edema
Event|Event|General Exam|3291,3296|true|false|false|||edema
Finding|Pathologic Function|General Exam|3291,3296|true|false|false|C0013604|Edema|edema
Anatomy|Body System|General Exam|3301,3305|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|General Exam|3301,3305|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|General Exam|3301,3305|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|General Exam|3301,3305|false|false|false|||SKIN
Finding|Body Substance|General Exam|3301,3305|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|General Exam|3301,3305|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Disorder|Disease or Syndrome|General Exam|3315,3319|true|false|false|C5779629|Eruption of skin (disorder)|rash
Event|Event|General Exam|3315,3319|true|false|false|||rash
Finding|Pathologic Function|General Exam|3315,3319|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|General Exam|3315,3319|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Event|Event|General Exam|3324,3334|false|false|false|||NEUROLOGIC
Event|Event|General Exam|3376,3385|false|false|false|||sensation
Finding|Finding|General Exam|3376,3385|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|General Exam|3376,3385|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|General Exam|3376,3385|false|false|false|C2229507|sensory exam|sensation
Event|Event|General Exam|3393,3401|false|false|false|||strength
Finding|Idea or Concept|General Exam|3393,3401|false|false|false|C0808080|Strength (attribute)|strength
Finding|Finding|General Exam|3422,3430|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|General Exam|3422,3430|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|General Exam|3422,3430|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|General Exam|3422,3442|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAMINATION
Procedure|Health Care Activity|General Exam|3422,3442|false|false|false|C0031809|Physical Examination|PHYSICAL EXAMINATION
Event|Activity|General Exam|3431,3442|false|false|false|C4321457|Examination|EXAMINATION
Event|Event|General Exam|3431,3442|false|false|false|||EXAMINATION
Procedure|Health Care Activity|General Exam|3431,3442|false|false|false|C0031809;C0582103|Medical Examination;Physical Examination|EXAMINATION
Finding|Body Substance|General Exam|3446,3455|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|3446,3455|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|3446,3455|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|3446,3455|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|General Exam|3493,3499|false|false|false|||VITALS
Event|Event|General Exam|3546,3553|false|false|false|||GENERAL
Finding|Classification|General Exam|3546,3553|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|General Exam|3546,3553|false|false|false|C3812897|General medical service|GENERAL
Event|Event|General Exam|3555,3563|true|false|false|||Pleasant
Finding|Mental Process|General Exam|3555,3563|true|false|false|C2987187|Pleasant|Pleasant
Finding|Finding|General Exam|3565,3569|true|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|3570,3579|true|false|false|||appearing
Finding|Idea or Concept|General Exam|3587,3595|true|false|false|C0750489|apparent|apparent
Event|Event|General Exam|3596,3604|true|false|false|||distress
Finding|Finding|General Exam|3596,3604|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|General Exam|3596,3604|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|General Exam|3609,3614|false|false|false|C1512338|HEENT|HEENT
Event|Event|General Exam|3616,3629|true|false|false|||Normocephalic
Event|Event|General Exam|3631,3641|true|false|false|||atraumatic
Anatomy|Body Part, Organ, or Organ Component|General Exam|3646,3658|true|false|false|C0009758|conjunctiva|conjunctival
Finding|Functional Concept|General Exam|3646,3658|true|false|false|C1522483|Conjunctival Route of Administration|conjunctival
Finding|Finding|General Exam|3646,3665|true|false|false|C2071267|Conjunctival pallor|conjunctival pallor
Event|Event|General Exam|3659,3665|true|false|false|||pallor
Finding|Finding|General Exam|3659,3665|true|false|false|C0241137|Pallor of skin|pallor
Anatomy|Body Part, Organ, or Organ Component|General Exam|3670,3677|true|false|false|C0036410|Sclera|scleral
Finding|Finding|General Exam|3670,3685|true|false|false|C0240962|Scleral icterus|scleral icterus
Finding|Sign or Symptom|General Exam|3678,3685|true|false|false|C0022346|Icterus|icterus
Event|Event|General Exam|3687,3693|false|false|false|||PERRLA
Finding|Finding|General Exam|3687,3693|false|false|false|C2143306|PERRLA|PERRLA
Event|Event|General Exam|3695,3699|false|false|false|||EOMI
Event|Event|General Exam|3704,3709|false|false|false|||clear
Finding|Idea or Concept|General Exam|3704,3709|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Location or Region|General Exam|3714,3718|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|General Exam|3714,3718|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|General Exam|3714,3718|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|General Exam|3720,3726|true|false|false|||Supple
Finding|Functional Concept|General Exam|3720,3726|true|false|false|C0332254|Supple|Supple
Anatomy|Body Part, Organ, or Organ Component|General Exam|3731,3734|true|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|General Exam|3731,3734|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|General Exam|3731,3734|true|false|false|||LAD
Finding|Gene or Genome|General Exam|3731,3734|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Disorder|Disease or Syndrome|General Exam|3739,3750|true|false|false|C0018021|Goiter|thyromegaly
Event|Event|General Exam|3739,3750|true|false|false|||thyromegaly
Event|Event|General Exam|3752,3755|true|false|false|||JVP
Finding|Finding|General Exam|3752,3755|true|false|false|C0428897|Jugular venous pressure|JVP
Anatomy|Body Part, Organ, or Organ Component|General Exam|3765,3772|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|General Exam|3765,3772|false|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Event|General Exam|3791,3798|true|false|false|||murmurs
Finding|Finding|General Exam|3791,3798|true|false|false|C0018808|Heart murmur|murmurs
Event|Event|General Exam|3799,3803|true|false|false|||rubs
Finding|Finding|General Exam|3799,3803|true|false|false|C0232267|Pericardial friction rub|rubs
Event|Event|General Exam|3807,3814|true|false|false|||gallops
Anatomy|Body Part, Organ, or Organ Component|General Exam|3819,3828|false|false|false|C0024109|Lung|PULMONARY
Attribute|Clinical Attribute|General Exam|3819,3828|false|false|false|C2707265||PULMONARY
Finding|Finding|General Exam|3819,3828|false|false|false|C4522268|Pulmonary (intended site)|PULMONARY
Drug|Inorganic Chemical|General Exam|3860,3863|true|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|General Exam|3860,3863|true|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|General Exam|3860,3863|true|false|false|C0001861;C3536832|Air (substance);air|air
Finding|Finding|General Exam|3860,3863|true|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|General Exam|3860,3863|true|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|General Exam|3860,3863|true|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Event|Event|General Exam|3864,3869|true|false|false|||entry
Finding|Functional Concept|General Exam|3864,3869|true|false|false|C1550548;C1705654|Entry (data);entry - ActRelationshipCheckpoint|entry
Finding|Intellectual Product|General Exam|3864,3869|true|false|false|C1550548;C1705654|Entry (data);entry - ActRelationshipCheckpoint|entry
Event|Event|General Exam|3874,3881|true|false|false|||wheezes
Finding|Sign or Symptom|General Exam|3874,3881|true|false|false|C0043144|Wheezing|wheezes
Anatomy|Body Location or Region|General Exam|3890,3894|true|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|General Exam|3890,3894|true|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|General Exam|3890,3894|true|false|false|C0024115|Lung diseases|lung
Finding|Finding|General Exam|3890,3894|true|false|false|C0740941|Lung Problem|lung
Event|Event|General Exam|3895,3901|true|false|false|||fields
Anatomy|Body Location or Region|General Exam|3905,3912|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|General Exam|3905,3912|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|General Exam|3905,3912|false|false|false|||ABDOMEN
Finding|Finding|General Exam|3905,3912|false|false|false|C0941288|Abdomen problem|ABDOMEN
Anatomy|Body Part, Organ, or Organ Component|General Exam|3921,3926|false|false|false|C0021853|Intestines|bowel
Finding|Finding|General Exam|3921,3933|false|false|false|C0232693|Bowel sounds|bowel sounds
Event|Event|General Exam|3927,3933|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|General Exam|3927,3933|false|false|false|C0037709||sounds
Disorder|Disease or Syndrome|General Exam|3935,3939|true|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|General Exam|3935,3939|true|false|false|||soft
Event|Event|General Exam|3972,3984|true|false|false|||organomegaly
Finding|Finding|General Exam|3972,3984|true|false|false|C4054315|Organomegaly|organomegaly
Anatomy|Body Part, Organ, or Organ Component|General Exam|3989,4000|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Event|Event|General Exam|4002,4006|true|false|false|||Warm
Finding|Finding|General Exam|4002,4006|true|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|4002,4006|true|false|false|C0687712|warming process|Warm
Finding|Finding|General Exam|4008,4012|true|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|4013,4021|true|false|false|||perfused
Event|Event|General Exam|4026,4034|true|false|false|||cyanosis
Finding|Sign or Symptom|General Exam|4026,4034|true|false|false|C0010520|Cyanosis|cyanosis
Disorder|Anatomical Abnormality|General Exam|4036,4044|true|false|false|C0149651|Clubbing|clubbing
Event|Event|General Exam|4036,4044|true|false|false|||clubbing
Attribute|Clinical Attribute|General Exam|4049,4054|true|false|false|C1717255||edema
Event|Event|General Exam|4049,4054|true|false|false|||edema
Finding|Pathologic Function|General Exam|4049,4054|true|false|false|C0013604|Edema|edema
Anatomy|Body System|General Exam|4059,4063|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|General Exam|4059,4063|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|General Exam|4059,4063|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|General Exam|4059,4063|false|false|false|||SKIN
Finding|Body Substance|General Exam|4059,4063|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|General Exam|4059,4063|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Disorder|Disease or Syndrome|General Exam|4073,4077|true|false|false|C5779629|Eruption of skin (disorder)|rash
Event|Event|General Exam|4073,4077|true|false|false|||rash
Finding|Pathologic Function|General Exam|4073,4077|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|General Exam|4073,4077|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Event|Event|General Exam|4082,4092|false|false|false|||NEUROLOGIC
Event|Event|General Exam|4134,4143|false|false|false|||sensation
Finding|Finding|General Exam|4134,4143|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|General Exam|4134,4143|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|General Exam|4134,4143|false|false|false|C2229507|sensory exam|sensation
Event|Event|General Exam|4151,4159|false|false|false|||strength
Finding|Idea or Concept|General Exam|4151,4159|false|false|false|C0808080|Strength (attribute)|strength
Event|Event|General Exam|4199,4203|false|false|false|||LABS
Lab|Laboratory or Test Result|General Exam|4199,4203|false|false|false|C0587081|Laboratory test finding|LABS
Procedure|Health Care Activity|General Exam|4207,4216|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Disorder|Disease or Syndrome|General Exam|4249,4254|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4249,4254|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4249,4254|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|4255,4258|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|4263,4266|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|4263,4266|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|4263,4266|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|4272,4275|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|4272,4275|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|4272,4275|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|4272,4275|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|4281,4284|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|4281,4284|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|4290,4293|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|4290,4293|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|4290,4293|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|4290,4293|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|4290,4293|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|4298,4301|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|4298,4301|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|4298,4301|false|false|false|||MCH
Finding|Gene or Genome|General Exam|4298,4301|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|4298,4301|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|4298,4301|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|4307,4311|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|4307,4311|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|4340,4343|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|4360,4365|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4360,4365|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4360,4365|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Body Substance|General Exam|4378,4384|false|false|false|C0024202|Lymph|Lymphs
Drug|Antibiotic|General Exam|4390,4395|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|General Exam|4390,4395|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|General Exam|4390,4395|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|General Exam|4401,4404|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Event|Event|General Exam|4401,4404|false|false|false|||Eos
Finding|Gene or Genome|General Exam|4401,4404|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|General Exam|4506,4511|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4506,4511|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4506,4511|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|4516,4519|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|General Exam|4516,4519|false|false|false|||PTT
Procedure|Laboratory Procedure|General Exam|4516,4519|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|General Exam|4541,4546|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4541,4546|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|4547,4550|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|4567,4572|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4567,4572|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4567,4572|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|4567,4580|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|4567,4580|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|4567,4580|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|4573,4580|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|4573,4580|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|4573,4580|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|4573,4580|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|4573,4580|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|4573,4580|false|false|false|C0337438|Glucose measurement|Glucose
Disorder|Disease or Syndrome|General Exam|4657,4662|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4657,4662|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4657,4662|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|4663,4666|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|4663,4666|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|General Exam|4663,4666|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|General Exam|4663,4666|false|false|false|||ALT
Finding|Gene or Genome|General Exam|4663,4666|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|General Exam|4663,4666|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|General Exam|4663,4666|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|General Exam|4663,4666|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|General Exam|4671,4674|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|General Exam|4671,4674|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|4671,4674|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|General Exam|4671,4674|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|General Exam|4671,4674|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|General Exam|4671,4674|false|false|false|||AST
Finding|Gene or Genome|General Exam|4671,4674|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|4678,4685|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|General Exam|4678,4685|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|General Exam|4713,4718|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4713,4718|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4713,4718|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|4719,4725|false|false|false|C0023764|lipase|Lipase
Drug|Enzyme|General Exam|4719,4725|false|false|false|C0023764|lipase|Lipase
Drug|Pharmacologic Substance|General Exam|4719,4725|false|false|false|C0023764|lipase|Lipase
Procedure|Laboratory Procedure|General Exam|4719,4725|false|false|false|C0373670|Lipase measurement|Lipase
Disorder|Disease or Syndrome|General Exam|4741,4746|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4741,4746|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4741,4746|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|4761,4767|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Drug|Hormone|General Exam|4761,4767|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Disorder|Disease or Syndrome|General Exam|4784,4789|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4784,4789|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4784,4789|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|4784,4797|false|false|false|C0853248|Blood albumin|BLOOD Albumin
Drug|Amino Acid, Peptide, or Protein|General Exam|4790,4797|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Biologically Active Substance|General Exam|4790,4797|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Pharmacologic Substance|General Exam|4790,4797|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Event|Event|General Exam|4790,4797|false|false|false|||Albumin
Finding|Gene or Genome|General Exam|4790,4797|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Finding|Physiologic Function|General Exam|4790,4797|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Procedure|Laboratory Procedure|General Exam|4790,4797|false|false|false|C0201838|Albumin measurement|Albumin
Event|Event|General Exam|4803,4807|false|false|false|||LABS
Lab|Laboratory or Test Result|General Exam|4803,4807|false|false|false|C0587081|Laboratory test finding|LABS
Event|Event|General Exam|4811,4821|false|false|false|||DISHCHARGE
Disorder|Disease or Syndrome|General Exam|4855,4860|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4855,4860|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4855,4860|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|4861,4864|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|4871,4874|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|4871,4874|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|4871,4874|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|4880,4883|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|4880,4883|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|4880,4883|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|4880,4883|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|4889,4892|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|4889,4892|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|4899,4902|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|4899,4902|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|4899,4902|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|4899,4902|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|4899,4902|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|4906,4909|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|4906,4909|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|4906,4909|false|false|false|||MCH
Finding|Gene or Genome|General Exam|4906,4909|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|4906,4909|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|4906,4909|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|4915,4919|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|4915,4919|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|4948,4951|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|4968,4973|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4968,4973|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|4974,4977|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|4994,4999|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4994,4999|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4994,4999|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|4994,5007|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|4994,5007|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|4994,5007|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|5000,5007|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|5000,5007|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|5000,5007|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|5000,5007|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|5000,5007|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|5000,5007|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|5052,5056|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|5052,5056|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|5052,5056|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|5081,5086|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|5081,5086|false|false|false|||BLOOD
Finding|Body Substance|General Exam|5081,5086|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|5081,5094|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|General Exam|5087,5094|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|5087,5094|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|5087,5094|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|5087,5094|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|5087,5094|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|General Exam|5087,5094|false|false|false|||Calcium
Finding|Physiologic Function|General Exam|5087,5094|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|5087,5094|false|false|false|C0201925|Calcium measurement|Calcium
Event|Event|General Exam|5117,5124|false|false|false|||IMAGING
Finding|Finding|General Exam|5117,5124|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|General Exam|5117,5124|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Event|Event|General Exam|5139,5142|false|false|false|||CXR
Procedure|Diagnostic Procedure|General Exam|5139,5142|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Intellectual Product|General Exam|5147,5152|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Location or Region|General Exam|5153,5168|true|false|false|C0553534|Cardiopulmonary|cardiopulmonary
Disorder|Disease or Syndrome|General Exam|5153,5168|true|false|false|C4072686|Cardiovascular disease+Pulmonary disease|cardiopulmonary
Anatomy|Body Part, Organ, or Organ Component|General Exam|5169,5176|true|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|General Exam|5169,5176|true|false|false|C1951340|Process Pharmacologic Substance|process
Event|Event|General Exam|5169,5176|true|false|false|||process
Finding|Functional Concept|General Exam|5169,5176|true|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|General Exam|5169,5176|true|false|false|C1522240|Process|process
Event|Event|Hospital Course|5218,5225|false|false|false|||history
Finding|Conceptual Entity|Hospital Course|5218,5225|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|5218,5225|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|5218,5225|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|5218,5228|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|Hospital Course|5229,5233|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|5229,5233|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|5229,5233|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|5229,5233|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|Hospital Course|5237,5241|false|false|false|||home
Finding|Idea or Concept|Hospital Course|5237,5241|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|5237,5241|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|5237,5241|false|false|false|C1553498|home health encounter|home
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5246,5252|false|false|false|C0018792|Heart Atrium|atrial
Attribute|Clinical Attribute|Hospital Course|5246,5265|false|false|false|C2926591||atrial fibrillation
Disorder|Disease or Syndrome|Hospital Course|5246,5265|false|false|false|C0004238|Atrial Fibrillation|atrial fibrillation
Lab|Laboratory or Test Result|Hospital Course|5246,5265|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|atrial fibrillation
Disorder|Disease or Syndrome|Hospital Course|5253,5265|false|false|false|C0232197|Fibrillation|fibrillation
Event|Event|Hospital Course|5253,5265|false|false|false|||fibrillation
Drug|Organic Chemical|Hospital Course|5270,5278|false|false|false|C1831808|apixaban|apixaban
Drug|Pharmacologic Substance|Hospital Course|5270,5278|false|false|false|C1831808|apixaban|apixaban
Event|Event|Hospital Course|5270,5278|false|false|false|||apixaban
Disorder|Disease or Syndrome|Hospital Course|5280,5292|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|Hospital Course|5280,5292|false|false|false|||hypertension
Disorder|Disease or Syndrome|Hospital Course|5294,5297|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5294,5297|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|5294,5297|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Hospital Course|5294,5297|false|false|false|||CAD
Finding|Gene or Genome|Hospital Course|5294,5297|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|5294,5297|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|5294,5297|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5294,5297|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|Hospital Course|5299,5313|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|hyperlipidemia
Event|Event|Hospital Course|5299,5313|false|false|false|||hyperlipidemia
Finding|Finding|Hospital Course|5299,5313|false|false|false|C0428465|Serum lipids high (finding)|hyperlipidemia
Event|Event|Hospital Course|5319,5328|false|false|false|||recurrent
Event|Event|Hospital Course|5330,5345|false|false|false|||hospitalization
Procedure|Health Care Activity|Hospital Course|5330,5345|false|false|false|C0019993|Hospitalization|hospitalization
Disorder|Disease or Syndrome|Hospital Course|5350,5354|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|5350,5354|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|5350,5354|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|5350,5354|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|Hospital Course|5350,5367|false|false|false|C0740304|COPD exacerbation|COPD exacerbation
Event|Event|Hospital Course|5355,5367|false|false|false|||exacerbation
Finding|Finding|Hospital Course|5355,5367|false|false|false|C4086268|Exacerbation|exacerbation
Event|Event|Hospital Course|5397,5406|false|false|false|||presented
Event|Event|Hospital Course|5412,5419|false|false|false|||dyspnea
Finding|Finding|Hospital Course|5412,5419|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|Hospital Course|5412,5419|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Event|Event|Hospital Course|5434,5442|false|false|false|||wheezing
Finding|Sign or Symptom|Hospital Course|5434,5442|false|false|false|C0043144|Wheezing|wheezing
Disorder|Neoplastic Process|Hospital Course|5443,5452|false|false|false|C0027627|Neoplasm Metastasis|secondary
Event|Event|Hospital Course|5443,5452|false|false|false|||secondary
Finding|Functional Concept|Hospital Course|5443,5452|false|false|false|C1522484|metastatic qualifier|secondary
Event|Event|Hospital Course|5457,5463|false|false|false|||severe
Finding|Finding|Hospital Course|5457,5463|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Hospital Course|5457,5463|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|Hospital Course|5464,5468|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|5464,5468|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|5464,5468|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|5464,5468|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|Hospital Course|5483,5487|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|5483,5487|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|5483,5487|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|5483,5487|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|Hospital Course|5483,5500|false|false|false|C0740304|COPD exacerbation|COPD exacerbation
Event|Event|Hospital Course|5488,5500|false|false|false|||exacerbation
Finding|Finding|Hospital Course|5488,5500|false|false|false|C4086268|Exacerbation|exacerbation
Finding|Body Substance|Hospital Course|5502,5509|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|5502,5509|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|5502,5509|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|5510,5519|false|false|false|||presented
Event|Event|Hospital Course|5525,5534|false|false|false|||increased
Finding|Finding|Hospital Course|5525,5534|false|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Functional Concept|Hospital Course|5525,5534|false|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Event|Event|Hospital Course|5536,5543|false|false|false|||dyspnea
Finding|Finding|Hospital Course|5536,5543|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|Hospital Course|5536,5543|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Finding|Hospital Course|5548,5564|false|false|false|C2089439|diffuse wheezing|diffuse wheezing
Event|Event|Hospital Course|5556,5564|false|false|false|||wheezing
Finding|Sign or Symptom|Hospital Course|5556,5564|false|false|false|C0043144|Wheezing|wheezing
Finding|Finding|Hospital Course|5566,5572|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|5566,5572|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Disorder|Neoplastic Process|Hospital Course|5573,5582|false|true|false|C0027627|Neoplasm Metastasis|secondary
Event|Event|Hospital Course|5573,5582|false|false|false|||secondary
Finding|Functional Concept|Hospital Course|5573,5582|false|true|false|C1522484|metastatic qualifier|secondary
Disorder|Disease or Syndrome|Hospital Course|5586,5590|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|5586,5590|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|5586,5590|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|5586,5590|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|Hospital Course|5592,5604|false|false|false|||exacerbation
Finding|Finding|Hospital Course|5592,5604|false|false|false|C4086268|Exacerbation|exacerbation
Event|Event|Hospital Course|5616,5623|false|false|false|||history
Finding|Conceptual Entity|Hospital Course|5616,5623|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|5616,5623|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|5616,5623|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|5616,5626|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|Hospital Course|5646,5650|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|5646,5650|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|5646,5650|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|5646,5650|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|Hospital Course|5652,5668|false|false|false|||hospitalizations
Procedure|Health Care Activity|Hospital Course|5652,5668|false|false|false|C0019993|Hospitalization|hospitalizations
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5683,5692|false|false|false|C0024109|Lung|Pulmonary
Attribute|Clinical Attribute|Hospital Course|5683,5692|false|false|false|C2707265||Pulmonary
Finding|Finding|Hospital Course|5683,5692|false|false|false|C4522268|Pulmonary (intended site)|Pulmonary
Finding|Body Substance|Hospital Course|5694,5701|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|5694,5701|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|5694,5701|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|Hospital Course|5694,5705|false|false|false|C0332310|Has patient|patient has
Event|Event|Hospital Course|5706,5712|false|false|false|||severe
Finding|Finding|Hospital Course|5706,5712|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Hospital Course|5706,5712|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|Hospital Course|5714,5718|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|5714,5718|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|5714,5718|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|5714,5718|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Functional Concept|Hospital Course|5732,5743|false|false|false|C0549186|Obstructed|obstructive
Event|Event|Hospital Course|5744,5752|false|false|false|||deficits
Event|Event|Hospital Course|5756,5760|false|false|false|||PFTs
Finding|Finding|Hospital Course|5764,5768|false|false|false|C5575035|Well (answer to question)|well
Finding|Finding|Hospital Course|5777,5783|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Hospital Course|5777,5783|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Finding|Hospital Course|5777,5792|false|false|false|C0436345|Symptom severe|severe symptoms
Event|Event|Hospital Course|5784,5792|false|false|false|||symptoms
Finding|Functional Concept|Hospital Course|5784,5792|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Hospital Course|5784,5792|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Functional Concept|Hospital Course|5798,5805|false|false|false|C0443144|At rest (qualifier value)|at rest
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5801,5805|false|false|false|C1742913|REST protein, human|rest
Drug|Biologically Active Substance|Hospital Course|5801,5805|false|false|false|C1742913|REST protein, human|rest
Finding|Daily or Recreational Activity|Hospital Course|5801,5805|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Gene or Genome|Hospital Course|5801,5805|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Molecular Function|Hospital Course|5801,5805|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Finding|Hospital Course|5810,5814|false|false|false|C5575035|Well (answer to question)|well
Event|Event|Hospital Course|5837,5850|false|false|false|||exacerbations
Finding|Finding|Hospital Course|5858,5864|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|5858,5864|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|Hospital Course|5865,5876|false|false|false|||approaching
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5877,5880|false|false|false|C0082420|Endoglin, human|end
Drug|Immunologic Factor|Hospital Course|5877,5880|false|false|false|C0082420|Endoglin, human|end
Finding|Functional Concept|Hospital Course|5877,5880|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Finding|Gene or Genome|Hospital Course|5877,5880|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Attribute|Clinical Attribute|Hospital Course|5881,5886|false|false|false|C1300072|Tumor stage|stage
Disorder|Disease or Syndrome|Hospital Course|5887,5894|false|false|false|C0012634|Disease|disease
Event|Event|Hospital Course|5887,5894|false|false|false|||disease
Event|Event|Hospital Course|5900,5909|false|false|false|||continued
Drug|Organic Chemical|Hospital Course|5910,5916|false|false|false|C0965130|Advair|Advair
Drug|Pharmacologic Substance|Hospital Course|5910,5916|false|false|false|C0965130|Advair|Advair
Disorder|Mental or Behavioral Dysfunction|Hospital Course|5924,5927|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5924,5927|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|5924,5927|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|5924,5927|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|5924,5927|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|5929,5936|false|false|false|C0905678|Spiriva|Spiriva
Drug|Pharmacologic Substance|Hospital Course|5929,5936|false|false|false|C0905678|Spiriva|Spiriva
Event|Event|Hospital Course|5929,5936|false|false|false|||Spiriva
Drug|Pharmacologic Substance|Hospital Course|5947,5957|false|false|false|C2064916|nebulizers (medication)|nebulizers
Event|Event|Hospital Course|5947,5957|false|false|false|||nebulizers
Drug|Organic Chemical|Hospital Course|5964,5976|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|Hospital Course|5964,5976|false|false|false|C0039771|theophylline|theophylline
Event|Event|Hospital Course|5964,5976|false|false|false|||theophylline
Procedure|Laboratory Procedure|Hospital Course|5964,5976|false|false|false|C0039773|Assay of theophylline|theophylline
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5978,5987|false|false|false|C0024109|Lung|Pulmonary
Attribute|Clinical Attribute|Hospital Course|5978,5987|false|false|false|C2707265||Pulmonary
Finding|Finding|Hospital Course|5978,5987|false|false|false|C4522268|Pulmonary (intended site)|Pulmonary
Event|Event|Hospital Course|5988,5999|false|false|false|||recommended
Finding|Functional Concept|Hospital Course|6000,6010|false|false|false|C1524062|Additional|additional
Drug|Organic Chemical|Hospital Course|6011,6021|false|false|false|C0054201|budesonide|budesonide
Drug|Pharmacologic Substance|Hospital Course|6011,6021|false|false|false|C0054201|budesonide|budesonide
Event|Event|Hospital Course|6011,6021|false|false|false|||budesonide
Event|Event|Hospital Course|6023,6031|false|false|false|||inhalers
Finding|Social Behavior|Hospital Course|6035,6040|false|false|false|C0683607|allowing|allow
Event|Event|Hospital Course|6041,6050|false|false|false|||reduction
Finding|Finding|Hospital Course|6041,6050|false|false|false|C0392756|Reduced|reduction
Phenomenon|Natural Phenomenon or Process|Hospital Course|6041,6050|false|false|false|C0301630|Reduction (chemical)|reduction
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6041,6050|false|false|false|C1293152;C4551656|Reduction procedure;Surgical reduction|reduction
Drug|Hormone|Hospital Course|6057,6067|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|Hospital Course|6057,6067|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|Hospital Course|6057,6067|false|false|false|C0032952|prednisone|prednisone
Event|Event|Hospital Course|6068,6072|false|false|false|||dose
Drug|Hormone|Hospital Course|6074,6084|false|false|false|C0032952|prednisone|Prednisone
Drug|Organic Chemical|Hospital Course|6074,6084|false|false|false|C0032952|prednisone|Prednisone
Drug|Pharmacologic Substance|Hospital Course|6074,6084|false|false|false|C0032952|prednisone|Prednisone
Event|Event|Hospital Course|6086,6090|false|false|false|||dose
Event|Event|Hospital Course|6095,6104|false|false|false|||increased
Finding|Body Substance|Hospital Course|6125,6132|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|6125,6132|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|6125,6132|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|6137,6143|false|false|false|||better
Finding|Idea or Concept|Hospital Course|6137,6143|false|false|false|C1550462|Observation Interpretation - better|better
Disorder|Disease or Syndrome|Hospital Course|6153,6157|false|false|false|C0270724|Infantile Neuroaxonal Dystrophy|plan
Event|Event|Hospital Course|6153,6157|false|false|false|||plan
Finding|Functional Concept|Hospital Course|6153,6157|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Intellectual Product|Hospital Course|6153,6157|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Mental Process|Hospital Course|6153,6157|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Finding|Hospital Course|6167,6171|false|false|false|C0043084|Weaning|wean
Finding|Body Substance|Hospital Course|6200,6207|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|6200,6207|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|6200,6207|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|6213,6220|false|false|false|||started
Event|Event|Hospital Course|6224,6231|false|false|false|||chronic
Finding|Intellectual Product|Hospital Course|6224,6231|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Hospital Course|6224,6231|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Drug|Antibiotic|Hospital Course|6232,6244|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|Hospital Course|6232,6244|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|Hospital Course|6232,6244|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Event|Event|Hospital Course|6232,6244|false|false|false|||azithromycin
Finding|Intellectual Product|Hospital Course|6249,6256|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Hospital Course|6249,6256|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Event|Event|Hospital Course|6283,6293|false|false|false|||discussion
Finding|Social Behavior|Hospital Course|6283,6293|false|false|false|C2584313|Discussion (communication)|discussion
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6283,6293|false|false|false|C0557061|Discussion (procedure)|discussion
Event|Event|Hospital Course|6311,6317|false|false|false|||agreed
Event|Event|Hospital Course|6321,6325|false|false|false|||stop
Drug|Antibiotic|Hospital Course|6327,6339|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|Hospital Course|6327,6339|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|Hospital Course|6327,6339|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Event|Event|Hospital Course|6327,6339|false|false|false|||azithromycin
Event|Event|Hospital Course|6343,6352|false|false|false|||discharge
Finding|Body Substance|Hospital Course|6343,6352|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|6343,6352|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|6343,6352|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|6343,6352|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|Hospital Course|6360,6369|false|false|false|||inability
Event|Event|Hospital Course|6373,6380|false|false|false|||monitor
Event|Event|Hospital Course|6389,6393|false|false|false|||week
Finding|Intellectual Product|Hospital Course|6389,6393|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|Hospital Course|6400,6409|false|false|false|||discharge
Finding|Body Substance|Hospital Course|6400,6409|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|6400,6409|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|6400,6409|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|6400,6409|false|false|false|C0030685|Patient Discharge|discharge
Disorder|Disease or Syndrome|Hospital Course|6416,6420|false|false|false|C0270724|Infantile Neuroaxonal Dystrophy|plan
Event|Event|Hospital Course|6416,6420|false|false|false|||plan
Finding|Functional Concept|Hospital Course|6416,6420|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Intellectual Product|Hospital Course|6416,6420|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Mental Process|Hospital Course|6416,6420|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Event|Event|Hospital Course|6424,6431|false|false|false|||restart
Drug|Antibiotic|Hospital Course|6432,6444|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|Hospital Course|6432,6444|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|Hospital Course|6432,6444|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Event|Event|Hospital Course|6432,6444|false|false|false|||azithromycin
Finding|Intellectual Product|Hospital Course|6445,6449|false|false|false|C1720092|Once - dosing instruction fragment|once
Event|Event|Hospital Course|6462,6466|false|false|false|||able
Finding|Finding|Hospital Course|6462,6466|false|false|false|C1299581|Able (qualifier value)|able
Event|Event|Hospital Course|6470,6473|false|false|false|||see
Finding|Body Substance|Hospital Course|6478,6485|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|6478,6485|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|6478,6485|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Body Substance|Hospital Course|6487,6494|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|6487,6494|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|6487,6494|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|6503,6507|true|false|false|||want
Event|Event|Hospital Course|6511,6513|true|false|false|||go
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6518,6527|true|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Hospital Course|6518,6527|true|false|false|C2707265||pulmonary
Finding|Finding|Hospital Course|6518,6527|true|false|false|C4522268|Pulmonary (intended site)|pulmonary
Event|Event|Hospital Course|6528,6533|true|false|false|||rehab
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6528,6533|true|false|false|C0034991|Rehabilitation therapy|rehab
Event|Event|Hospital Course|6543,6547|false|false|false|||seen
Finding|Finding|Hospital Course|6551,6566|false|false|false|C0700049|Encounter due to palliative care|Palliative Care
Procedure|Health Care Activity|Hospital Course|6551,6566|false|false|false|C0030231;C3816218|Palliative Care;Palliative Nursing|Palliative Care
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6551,6566|false|false|false|C0030231;C3816218|Palliative Care;Palliative Nursing|Palliative Care
Event|Activity|Hospital Course|6562,6566|false|false|false|C1947933|care activity|Care
Event|Event|Hospital Course|6562,6566|false|false|false|||Care
Finding|Finding|Hospital Course|6562,6566|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Hospital Course|6562,6566|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Event|Event|Hospital Course|6571,6582|false|false|false|||recommended
Event|Event|Hospital Course|6584,6594|false|false|false|||initiation
Finding|Functional Concept|Hospital Course|6584,6594|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Finding|Genetic Function|Hospital Course|6584,6594|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Finding|Mental Process|Hospital Course|6584,6594|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Drug|Organic Chemical|Hospital Course|6598,6606|false|false|false|C0026549|morphine|morphine
Drug|Pharmacologic Substance|Hospital Course|6598,6606|false|false|false|C0026549|morphine|morphine
Drug|Biomedical or Dental Material|Hospital Course|6607,6613|false|false|false|C0302908;C1697794|Liquid Dosage Form;Liquid substance|liquid
Drug|Substance|Hospital Course|6607,6613|false|false|false|C0302908;C1697794|Liquid Dosage Form;Liquid substance|liquid
Event|Event|Hospital Course|6607,6613|false|false|false|||liquid
Finding|Finding|Hospital Course|6607,6613|false|false|false|C1304698|Liquid (finding)|liquid
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6607,6613|false|false|false|C0301571|Liquid diet|liquid
Drug|Biomedical or Dental Material|Hospital Course|6614,6624|false|false|false|C0038960;C1382107|Suspension substance;Suspensions|suspension
Drug|Substance|Hospital Course|6614,6624|false|false|false|C0038960;C1382107|Suspension substance;Suspensions|suspension
Event|Event|Hospital Course|6614,6624|false|false|false|||suspension
Finding|Functional Concept|Hospital Course|6614,6624|false|false|false|C1705537|Suspension (action)|suspension
Event|Event|Hospital Course|6628,6634|false|false|false|||needed
Event|Event|Hospital Course|6639,6648|false|false|false|||shortness
Finding|Body Substance|Hospital Course|6653,6659|false|false|false|C0225386|Breath|breath
Finding|Intellectual Product|Hospital Course|6664,6669|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Disorder|Disease or Syndrome|Hospital Course|6664,6683|false|false|false|C0022660;C2609414|Acute kidney injury;Kidney Failure, Acute|Acute kidney injury
Disorder|Injury or Poisoning|Hospital Course|6664,6683|false|false|false|C0022660;C2609414|Acute kidney injury;Kidney Failure, Acute|Acute kidney injury
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6670,6676|false|false|false|C0022646;C0227665|Both kidneys;Kidney|kidney
Disorder|Neoplastic Process|Hospital Course|6670,6676|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|kidney
Event|Event|Hospital Course|6670,6676|false|false|false|||kidney
Finding|Sign or Symptom|Hospital Course|6670,6676|false|false|false|C0812426|Kidney problem|kidney
Procedure|Diagnostic Procedure|Hospital Course|6670,6676|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6670,6676|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Disorder|Injury or Poisoning|Hospital Course|6670,6683|false|false|false|C0160420|Injury of kidney|kidney injury
Disorder|Injury or Poisoning|Hospital Course|6677,6683|false|false|false|C3263722;C3263723|Traumatic AND/OR non-traumatic injury;Traumatic injury|injury
Event|Event|Hospital Course|6677,6683|false|false|false|||injury
Drug|Biologically Active Substance|Hospital Course|6685,6695|false|false|false|C0010294|creatinine|Creatinine
Drug|Organic Chemical|Hospital Course|6685,6695|false|false|false|C0010294|creatinine|Creatinine
Event|Event|Hospital Course|6685,6695|false|false|false|||Creatinine
Finding|Physiologic Function|Hospital Course|6685,6695|false|false|false|C4551889|Creatinine metabolic function|Creatinine
Procedure|Laboratory Procedure|Hospital Course|6685,6695|false|false|false|C0201975|Creatinine measurement|Creatinine
Event|Event|Hospital Course|6709,6717|false|false|false|||elevated
Drug|Biomedical or Dental Material|Hospital Course|6733,6741|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|Hospital Course|6733,6741|false|false|false|||baseline
Finding|Idea or Concept|Hospital Course|6733,6741|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Finding|Hospital Course|6754,6760|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|6754,6760|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Intellectual Product|Hospital Course|6765,6769|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Event|Event|Hospital Course|6773,6779|false|false|false|||intake
Finding|Functional Concept|Hospital Course|6773,6779|false|false|false|C1512806|Intake|intake
Procedure|Health Care Activity|Hospital Course|6773,6779|false|false|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|intake
Drug|Biologically Active Substance|Hospital Course|6782,6792|false|false|false|C0010294|creatinine|Creatinine
Drug|Organic Chemical|Hospital Course|6782,6792|false|false|false|C0010294|creatinine|Creatinine
Event|Event|Hospital Course|6782,6792|false|false|false|||Creatinine
Finding|Physiologic Function|Hospital Course|6782,6792|false|false|false|C4551889|Creatinine metabolic function|Creatinine
Procedure|Laboratory Procedure|Hospital Course|6782,6792|false|false|false|C0201975|Creatinine measurement|Creatinine
Event|Event|Hospital Course|6796,6805|false|false|false|||discharge
Finding|Body Substance|Hospital Course|6796,6805|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|6796,6805|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|6796,6805|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|6796,6805|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|Hospital Course|6817,6824|false|false|false|||CHRONIC
Finding|Intellectual Product|Hospital Course|6817,6824|false|false|false|C1547296|Chronic - Admission Level of Care Code|CHRONIC
Procedure|Health Care Activity|Hospital Course|6817,6824|false|false|false|C1555457|Provision of recurring care for chronic illness|CHRONIC
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6858,6865|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|Anxiety
Event|Event|Hospital Course|6858,6865|false|false|false|||Anxiety
Finding|Sign or Symptom|Hospital Course|6858,6865|false|false|false|C0860603|Anxiety symptoms|Anxiety
Drug|Pharmacologic Substance|Hospital Course|6866,6874|false|false|false|C1950154|Insomnia homeopathic medication|Insomnia
Event|Event|Hospital Course|6866,6874|false|false|false|||Insomnia
Finding|Sign or Symptom|Hospital Course|6866,6874|false|false|false|C0917801|Sleeplessness|Insomnia
Event|Event|Hospital Course|6879,6888|false|false|false|||continued
Finding|Idea or Concept|Hospital Course|6889,6893|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|6889,6893|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|6889,6893|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|6894,6903|false|false|false|C0024002|lorazepam|lorazepam
Drug|Pharmacologic Substance|Hospital Course|6894,6903|false|false|false|C0024002|lorazepam|lorazepam
Event|Event|Hospital Course|6894,6903|false|false|false|||lorazepam
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6909,6915|false|false|false|C0018792|Heart Atrium|Atrial
Attribute|Clinical Attribute|Hospital Course|6909,6928|false|false|false|C2926591||Atrial fibrillation
Disorder|Disease or Syndrome|Hospital Course|6909,6928|false|false|false|C0004238|Atrial Fibrillation|Atrial fibrillation
Lab|Laboratory or Test Result|Hospital Course|6909,6928|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Atrial fibrillation
Disorder|Disease or Syndrome|Hospital Course|6916,6928|false|false|false|C0232197|Fibrillation|fibrillation
Event|Event|Hospital Course|6916,6928|false|false|false|||fibrillation
Event|Event|Hospital Course|6933,6942|false|false|false|||continued
Drug|Organic Chemical|Hospital Course|6943,6952|false|false|false|C0012373|diltiazem|diltiazem
Drug|Pharmacologic Substance|Hospital Course|6943,6952|false|false|false|C0012373|diltiazem|diltiazem
Event|Event|Hospital Course|6943,6952|false|false|false|||diltiazem
Event|Activity|Hospital Course|6957,6961|false|false|false|C0871208|Rating (action)|rate
Finding|Idea or Concept|Hospital Course|6957,6961|false|false|false|C1549480|Amount type - Rate|rate
Finding|Functional Concept|Hospital Course|6957,6969|false|false|false|C0489879|rate control|rate control
Drug|Organic Chemical|Hospital Course|6962,6969|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|Hospital Course|6962,6969|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|Hospital Course|6962,6969|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Event|Event|Hospital Course|6962,6969|false|false|false|||control
Finding|Conceptual Entity|Hospital Course|6962,6969|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|Hospital Course|6962,6969|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|Hospital Course|6962,6969|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Drug|Organic Chemical|Hospital Course|6975,6983|false|false|false|C1831808|apixaban|apixaban
Drug|Pharmacologic Substance|Hospital Course|6975,6983|false|false|false|C1831808|apixaban|apixaban
Event|Event|Hospital Course|6975,6983|false|false|false|||apixaban
Event|Event|Hospital Course|6988,7003|false|false|false|||anticoagulation
Finding|Finding|Hospital Course|6988,7003|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|Hospital Course|6988,7003|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6988,7003|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Disorder|Disease or Syndrome|Hospital Course|7011,7023|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|Hospital Course|7011,7023|false|false|false|||Hypertension
Event|Event|Hospital Course|7028,7037|false|false|false|||continued
Finding|Idea or Concept|Hospital Course|7038,7042|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|7038,7042|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|7038,7042|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|7043,7048|false|false|false|C0590690|Imdur|imdur
Drug|Pharmacologic Substance|Hospital Course|7043,7048|false|false|false|C0590690|Imdur|imdur
Event|Event|Hospital Course|7043,7048|false|false|false|||imdur
Drug|Organic Chemical|Hospital Course|7050,7069|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Drug|Pharmacologic Substance|Hospital Course|7050,7069|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Event|Event|Hospital Course|7050,7069|false|false|false|||hydrochlorothiazide
Drug|Organic Chemical|Hospital Course|7076,7085|false|false|false|C0012373|diltiazem|diltiazem
Drug|Pharmacologic Substance|Hospital Course|7076,7085|false|false|false|C0012373|diltiazem|diltiazem
Event|Event|Hospital Course|7076,7085|false|false|false|||diltiazem
Disorder|Disease or Syndrome|Hospital Course|7093,7096|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7093,7096|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|7093,7096|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Hospital Course|7093,7096|false|false|false|||CAD
Finding|Gene or Genome|Hospital Course|7093,7096|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|7093,7096|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|7093,7096|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7093,7096|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7098,7105|true|false|false|C0018787|Heart|Cardiac
Finding|Intellectual Product|Hospital Course|7098,7105|true|false|false|C1314974|Cardiac attachment|Cardiac
Disorder|Injury or Poisoning|Hospital Course|7098,7121|true|false|false|C0261588|Cardiac catheterisation as the cause of abnormal reaction of the patient, or of later complication, without mention of misadventure at the time of the procedure|Cardiac catheterization
Finding|Intellectual Product|Hospital Course|7098,7121|true|false|false|C1547981|Diagnostic Service Section ID - Cardiac Catheterization|Cardiac catheterization
Procedure|Diagnostic Procedure|Hospital Course|7098,7121|true|false|false|C0018795;C1548828|Cardiac Catheterization Procedures;Consent Type - Cardiac Catheterization|Cardiac catheterization
Procedure|Health Care Activity|Hospital Course|7098,7121|true|false|false|C0018795;C1548828|Cardiac Catheterization Procedures;Consent Type - Cardiac Catheterization|Cardiac catheterization
Event|Event|Hospital Course|7106,7121|true|false|false|||catheterization
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7106,7121|true|false|false|C0007430|Catheterization|catheterization
Event|Event|Hospital Course|7129,7135|true|false|false|||showed
Event|Event|Hospital Course|7139,7147|true|false|false|||evidence
Finding|Idea or Concept|Hospital Course|7139,7147|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Hospital Course|7139,7150|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Finding|Idea or Concept|Hospital Course|7152,7163|true|false|false|C0750502|Significant|significant
Event|Event|Hospital Course|7164,7172|true|false|false|||stenosis
Finding|Pathologic Function|Hospital Course|7164,7172|true|false|false|C1261287|Stenosis|stenosis
Event|Event|Hospital Course|7176,7186|true|false|false|||coronaries
Event|Event|Hospital Course|7188,7192|false|false|false|||ECHO
Procedure|Health Care Activity|Hospital Course|7188,7192|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7188,7192|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Event|Event|Hospital Course|7200,7206|true|false|false|||showed
Attribute|Clinical Attribute|Hospital Course|7243,7254|true|false|false|C1980023|Wall motion|wall motion
Phenomenon|Natural Phenomenon or Process|Hospital Course|7248,7254|true|false|false|C0026597|Motion|motion
Disorder|Congenital Abnormality|Hospital Course|7255,7268|true|false|false|C0000768|Congenital Abnormality|abnormalities
Event|Event|Hospital Course|7255,7268|true|false|false|||abnormalities
Finding|Functional Concept|Hospital Course|7255,7268|true|false|false|C0000769|teratologic|abnormalities
Event|Event|Hospital Course|7274,7283|false|false|false|||continued
Finding|Idea or Concept|Hospital Course|7284,7288|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|7284,7288|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|7284,7288|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|7289,7296|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|Hospital Course|7289,7296|false|false|false|C0004057|aspirin|aspirin
Event|Event|Hospital Course|7289,7296|false|false|false|||aspirin
Drug|Organic Chemical|Hospital Course|7301,7313|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|Hospital Course|7301,7313|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|Hospital Course|7301,7313|false|false|false|||atorvastatin
Disorder|Disease or Syndrome|Hospital Course|7319,7325|false|false|false|C0002871|Anemia|Anemia
Event|Event|Hospital Course|7319,7325|false|false|false|||Anemia
Event|Event|Hospital Course|7330,7339|false|false|false|||continued
Finding|Idea or Concept|Hospital Course|7340,7344|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|7340,7344|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|7340,7344|false|false|false|C1553498|home health encounter|home
Drug|Biologically Active Substance|Hospital Course|7345,7349|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|Hospital Course|7345,7349|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|Hospital Course|7345,7349|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Procedure|Laboratory Procedure|Hospital Course|7345,7349|false|false|false|C0337439|Iron measurement|iron
Drug|Inorganic Chemical|Hospital Course|7345,7361|false|false|false|C0721124|Iron Supplement|iron supplements
Drug|Pharmacologic Substance|Hospital Course|7345,7361|false|false|false|C0721124|Iron Supplement|iron supplements
Event|Event|Hospital Course|7350,7361|false|false|false|||supplements
Finding|Idea or Concept|Hospital Course|7368,7380|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Event|Event|Hospital Course|7381,7387|false|false|false|||ISSUES
Event|Event|Hospital Course|7395,7403|false|false|false|||Continue
Finding|Idea or Concept|Hospital Course|7395,7403|false|false|false|C0549178|Continuous|Continue
Drug|Organic Chemical|Hospital Course|7404,7410|false|false|false|C0965130|Advair|Advair
Drug|Pharmacologic Substance|Hospital Course|7404,7410|false|false|false|C0965130|Advair|Advair
Event|Event|Hospital Course|7404,7410|false|false|false|||Advair
Disorder|Mental or Behavioral Dysfunction|Hospital Course|7418,7421|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7418,7421|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|7418,7421|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|7418,7421|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|7418,7421|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|7423,7430|false|false|false|C0905678|Spiriva|Spiriva
Drug|Pharmacologic Substance|Hospital Course|7423,7430|false|false|false|C0905678|Spiriva|Spiriva
Event|Event|Hospital Course|7423,7430|false|false|false|||Spiriva
Drug|Organic Chemical|Hospital Course|7436,7448|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|Hospital Course|7436,7448|false|false|false|C0039771|theophylline|theophylline
Event|Event|Hospital Course|7436,7448|false|false|false|||theophylline
Procedure|Laboratory Procedure|Hospital Course|7436,7448|false|false|false|C0039773|Assay of theophylline|theophylline
Finding|Functional Concept|Hospital Course|7452,7456|false|false|false|C0947322;C1881534|Make - Instruction Imperative;Manufacturer Name|Make
Finding|Intellectual Product|Hospital Course|7452,7456|false|false|false|C0947322;C1881534|Make - Instruction Imperative;Manufacturer Name|Make
Finding|Intellectual Product|Hospital Course|7457,7461|false|false|false|C4724437|SURE Test|sure
Finding|Body Substance|Hospital Course|7462,7469|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|7462,7469|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|7462,7469|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|7470,7478|false|false|false|||receives
Drug|Pharmacologic Substance|Hospital Course|7488,7498|false|false|false|C2064916|nebulizers (medication)|nebulizers
Event|Event|Hospital Course|7488,7498|false|false|false|||nebulizers
Finding|Functional Concept|Hospital Course|7508,7518|false|false|false|C1524062|Additional|additional
Drug|Organic Chemical|Hospital Course|7519,7529|false|false|false|C0054201|budesonide|budesonide
Drug|Pharmacologic Substance|Hospital Course|7519,7529|false|false|false|C0054201|budesonide|budesonide
Event|Event|Hospital Course|7530,7538|false|false|false|||inhalers
Event|Event|Hospital Course|7542,7547|false|false|false|||allow
Event|Event|Hospital Course|7548,7557|false|false|false|||reduction
Finding|Finding|Hospital Course|7548,7557|false|false|false|C0392756|Reduced|reduction
Phenomenon|Natural Phenomenon or Process|Hospital Course|7548,7557|false|false|false|C0301630|Reduction (chemical)|reduction
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7548,7557|false|false|false|C1293152;C4551656|Reduction procedure;Surgical reduction|reduction
Drug|Hormone|Hospital Course|7565,7575|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|Hospital Course|7565,7575|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|Hospital Course|7565,7575|false|false|false|C0032952|prednisone|prednisone
Event|Event|Hospital Course|7576,7580|false|false|false|||dose
Drug|Food|Hospital Course|7584,7589|false|false|false|C0452588|Start brand of breakfast cereal|Start
Event|Event|Hospital Course|7584,7589|false|false|false|||Start
Finding|Intellectual Product|Hospital Course|7584,7589|false|false|false|C1552850|start - HtmlLinkType|Start
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7584,7589|false|false|false|C5447432|Collagen Tile Brachytherapy|Start
Event|Event|Hospital Course|7590,7597|false|false|false|||chronic
Finding|Intellectual Product|Hospital Course|7590,7597|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Hospital Course|7590,7597|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Drug|Antibiotic|Hospital Course|7598,7610|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|Hospital Course|7598,7610|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|Hospital Course|7598,7610|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Event|Event|Hospital Course|7598,7610|false|false|false|||azithromycin
Finding|Intellectual Product|Hospital Course|7615,7622|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Hospital Course|7615,7622|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Finding|Body Substance|Hospital Course|7644,7651|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|7644,7651|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|7644,7651|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|7656,7663|false|false|false|||started
Drug|Antibiotic|Hospital Course|7667,7679|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|Hospital Course|7667,7679|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|Hospital Course|7667,7679|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Event|Event|Hospital Course|7667,7679|false|false|false|||azithromycin
Finding|Idea or Concept|Hospital Course|7687,7695|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|Hospital Course|7728,7738|false|false|false|||discussion
Finding|Social Behavior|Hospital Course|7728,7738|false|false|false|C2584313|Discussion (communication)|discussion
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7728,7738|false|false|false|C0557061|Discussion (procedure)|discussion
Event|Event|Hospital Course|7756,7762|false|false|false|||agreed
Drug|Antibiotic|Hospital Course|7772,7784|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|Hospital Course|7772,7784|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|Hospital Course|7772,7784|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Event|Event|Hospital Course|7772,7784|false|false|false|||azithromycin
Event|Event|Hospital Course|7788,7797|false|false|false|||discharge
Finding|Body Substance|Hospital Course|7788,7797|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|7788,7797|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|7788,7797|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|7788,7797|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|Hospital Course|7805,7814|false|false|false|||inability
Event|Event|Hospital Course|7818,7825|false|false|false|||monitor
Finding|Intellectual Product|Hospital Course|7834,7838|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|Hospital Course|7845,7854|false|false|false|||discharge
Finding|Body Substance|Hospital Course|7845,7854|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|7845,7854|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|7845,7854|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|7845,7854|false|false|false|C0030685|Patient Discharge|discharge
Disorder|Disease or Syndrome|Hospital Course|7865,7869|false|false|false|C0270724|Infantile Neuroaxonal Dystrophy|plan
Event|Event|Hospital Course|7865,7869|false|false|false|||plan
Finding|Functional Concept|Hospital Course|7865,7869|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Intellectual Product|Hospital Course|7865,7869|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Mental Process|Hospital Course|7865,7869|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Drug|Antibiotic|Hospital Course|7881,7893|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|Hospital Course|7881,7893|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|Hospital Course|7881,7893|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Event|Event|Hospital Course|7881,7893|false|false|false|||azithromycin
Finding|Intellectual Product|Hospital Course|7895,7899|false|false|false|C1720092|Once - dosing instruction fragment|once
Event|Event|Hospital Course|7911,7915|false|false|false|||able
Finding|Finding|Hospital Course|7911,7915|false|false|false|C1299581|Able (qualifier value)|able
Event|Event|Hospital Course|7919,7922|false|false|false|||see
Finding|Body Substance|Hospital Course|7927,7934|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|7927,7934|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|7927,7934|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|7945,7954|false|false|false|||recommend
Finding|Intellectual Product|Hospital Course|7955,7964|false|false|false|C1547975;C4554598|Audiology - Clinical Class;Audiology Section ID|audiology
Event|Event|Hospital Course|7965,7972|false|false|false|||testing
Finding|Functional Concept|Hospital Course|7965,7972|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|testing
Finding|Intellectual Product|Hospital Course|7965,7972|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|testing
Finding|Body Substance|Hospital Course|7993,8000|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|7993,8000|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|7993,8000|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|8008,8015|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Hospital Course|8008,8015|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Drug|Antibiotic|Hospital Course|8016,8028|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|Hospital Course|8016,8028|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|Hospital Course|8016,8028|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Event|Event|Hospital Course|8016,8028|false|false|false|||azithromycin
Event|Event|Hospital Course|8031,8039|false|false|false|||Continue
Finding|Functional Concept|Hospital Course|8040,8052|false|false|false|C2348609|Supplement|supplemental
Finding|Finding|Hospital Course|8040,8059|false|false|false|C4534306|Supplemental oxygen|supplemental oxygen
Drug|Biologically Active Substance|Hospital Course|8053,8059|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|Hospital Course|8053,8059|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|Hospital Course|8053,8059|false|false|false|C0030054|oxygen|oxygen
Event|Event|Hospital Course|8053,8059|false|false|false|||oxygen
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8053,8059|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Drug|Organic Chemical|Hospital Course|8064,8071|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Drug|Pharmacologic Substance|Hospital Course|8064,8071|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Event|Event|Hospital Course|8064,8071|false|false|false|||comfort
Finding|Mental Process|Hospital Course|8064,8071|false|false|false|C1331418|Comfort|comfort
Finding|Functional Concept|Hospital Course|8074,8080|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|Follow
Finding|Intellectual Product|Hospital Course|8074,8080|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|Follow
Finding|Finding|Hospital Course|8074,8083|false|false|false|C0589120|Follow-up status|Follow up
Procedure|Health Care Activity|Hospital Course|8074,8083|false|false|false|C1522577|follow-up|Follow up
Event|Event|Hospital Course|8081,8083|false|false|false|||up
Event|Event|Hospital Course|8097,8106|false|false|false|||discharge
Finding|Body Substance|Hospital Course|8097,8106|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|8097,8106|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|8097,8106|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|8097,8106|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|Hospital Course|8110,8118|false|false|false|||Continue
Finding|Idea or Concept|Hospital Course|8110,8118|false|false|false|C0549178|Continuous|Continue
Drug|Organic Chemical|Hospital Course|8119,8126|false|false|false|C0591139|Bactrim|Bactrim
Drug|Pharmacologic Substance|Hospital Course|8119,8126|false|false|false|C0591139|Bactrim|Bactrim
Event|Event|Hospital Course|8127,8130|false|false|false|||PPX
Finding|Gene or Genome|Hospital Course|8127,8130|false|false|false|C1418850|PPP4C gene|PPX
Drug|Biomedical or Dental Material|Hospital Course|8134,8137|false|false|false|C0039225|Tablet Dosage Form|tab
Event|Event|Hospital Course|8138,8140|false|false|false|||SS
Finding|Finding|Hospital Course|8154,8162|false|false|false|C0231448;C5781021|Extended (finding);Extension|extended
Finding|Functional Concept|Hospital Course|8154,8162|false|false|false|C0231448;C5781021|Extended (finding);Extension|extended
Event|Event|Hospital Course|8163,8170|false|false|false|||courses
Drug|Organic Chemical|Hospital Course|8175,8183|false|false|false|C0038317|Steroids|steroids
Drug|Pharmacologic Substance|Hospital Course|8175,8183|false|false|false|C0038317|Steroids|steroids
Event|Event|Hospital Course|8175,8183|false|false|false|||steroids
Finding|Body Substance|Hospital Course|8187,8194|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|8187,8194|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|8187,8194|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|8199,8209|false|false|false|||discharged
Drug|Hormone|Hospital Course|8213,8223|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|Hospital Course|8213,8223|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|Hospital Course|8213,8223|false|false|false|C0032952|prednisone|prednisone
Event|Event|Hospital Course|8213,8223|false|false|false|||prednisone
Disorder|Disease or Syndrome|Hospital Course|8235,8239|false|false|false|C0270724|Infantile Neuroaxonal Dystrophy|plan
Event|Event|Hospital Course|8235,8239|false|false|false|||plan
Finding|Functional Concept|Hospital Course|8235,8239|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Intellectual Product|Hospital Course|8235,8239|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Mental Process|Hospital Course|8235,8239|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Event|Event|Hospital Course|8244,8249|false|false|false|||taper
Procedure|Health Care Activity|Hospital Course|8244,8249|false|false|false|C0441640||taper
Drug|Hormone|Hospital Course|8274,8284|false|false|false|C0032952|prednisone|Prednisone
Drug|Organic Chemical|Hospital Course|8274,8284|false|false|false|C0032952|prednisone|Prednisone
Drug|Pharmacologic Substance|Hospital Course|8274,8284|false|false|false|C0032952|prednisone|Prednisone
Finding|Idea or Concept|Hospital Course|8306,8309|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|Day
Finding|Intellectual Product|Hospital Course|8306,8309|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|Day
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8317,8320|false|false|false|C0082420|Endoglin, human|end
Drug|Immunologic Factor|Hospital Course|8317,8320|false|false|false|C0082420|Endoglin, human|end
Event|Event|Hospital Course|8317,8320|false|false|false|||end
Finding|Functional Concept|Hospital Course|8317,8320|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Finding|Gene or Genome|Hospital Course|8317,8320|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Drug|Hormone|Hospital Course|8327,8337|false|false|false|C0032952|prednisone|Prednisone
Drug|Organic Chemical|Hospital Course|8327,8337|false|false|false|C0032952|prednisone|Prednisone
Drug|Pharmacologic Substance|Hospital Course|8327,8337|false|false|false|C0032952|prednisone|Prednisone
Finding|Idea or Concept|Hospital Course|8359,8362|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|Day
Finding|Intellectual Product|Hospital Course|8359,8362|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|Day
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8370,8373|false|false|false|C0082420|Endoglin, human|end
Drug|Immunologic Factor|Hospital Course|8370,8373|false|false|false|C0082420|Endoglin, human|end
Event|Event|Hospital Course|8370,8373|false|false|false|||end
Finding|Functional Concept|Hospital Course|8370,8373|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Finding|Gene or Genome|Hospital Course|8370,8373|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Drug|Hormone|Hospital Course|8380,8390|false|false|false|C0032952|prednisone|Prednisone
Drug|Organic Chemical|Hospital Course|8380,8390|false|false|false|C0032952|prednisone|Prednisone
Drug|Pharmacologic Substance|Hospital Course|8380,8390|false|false|false|C0032952|prednisone|Prednisone
Finding|Idea or Concept|Hospital Course|8412,8415|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|Day
Finding|Intellectual Product|Hospital Course|8412,8415|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|Day
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8423,8426|false|false|false|C0082420|Endoglin, human|end
Drug|Immunologic Factor|Hospital Course|8423,8426|false|false|false|C0082420|Endoglin, human|end
Event|Event|Hospital Course|8423,8426|false|false|false|||end
Finding|Functional Concept|Hospital Course|8423,8426|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Finding|Gene or Genome|Hospital Course|8423,8426|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Finding|Idea or Concept|Hospital Course|8433,8436|false|false|false|C1548556|Etc.|etc
Event|Activity|Hospital Course|8442,8449|false|false|false|C3812666|Personal Contact|CONTACT
Event|Event|Hospital Course|8442,8449|false|false|false|||CONTACT
Finding|Functional Concept|Hospital Course|8442,8449|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Idea or Concept|Hospital Course|8442,8449|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Intellectual Product|Hospital Course|8442,8449|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Phenomenon|Phenomenon or Process|Hospital Course|8442,8449|false|false|false|C0392367|Physical contact|CONTACT
Disorder|Disease or Syndrome|Hospital Course|8464,8467|false|false|false|C0162531|Hereditary Coproporphyria|HCP
Event|Event|Hospital Course|8464,8467|false|false|false|||HCP
Finding|Gene or Genome|Hospital Course|8464,8467|false|false|false|C1335283;C1412376;C1413681;C1705637;C5780748|AMBP gene;AMBP wt Allele;CPOX gene;PTPN6 gene;PTPN6 wt Allele|HCP
Event|Event|Hospital Course|8476,8480|false|false|false|||CODE
Event|Occupational Activity|Hospital Course|8476,8480|false|false|false|C0009219|Coding|CODE
Finding|Intellectual Product|Hospital Course|8476,8480|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|CODE
Procedure|Health Care Activity|Hospital Course|8476,8487|false|false|false|C0742531|CODE STATUS|CODE STATUS
Attribute|Clinical Attribute|Hospital Course|8481,8487|false|false|false|C5889824||STATUS
Event|Event|Hospital Course|8481,8487|false|false|false|||STATUS
Finding|Idea or Concept|Hospital Course|8481,8487|false|false|false|C1546481|What subject filter - Status|STATUS
Event|Event|Hospital Course|8494,8503|false|false|false|||confirmed
Attribute|Clinical Attribute|Hospital Course|8507,8518|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|8507,8518|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|8507,8518|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|8507,8518|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|8507,8531|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|8522,8531|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|8522,8531|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|Hospital Course|8550,8560|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Hospital Course|8550,8560|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|Hospital Course|8550,8565|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|Hospital Course|8561,8565|false|false|false|||list
Finding|Intellectual Product|Hospital Course|8561,8565|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|Hospital Course|8569,8577|false|false|false|||accurate
Drug|Organic Chemical|Hospital Course|8582,8590|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Hospital Course|8582,8590|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Hospital Course|8582,8590|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|Hospital Course|8582,8590|false|false|false|||complete
Finding|Functional Concept|Hospital Course|8582,8590|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|8582,8590|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|Hospital Course|8595,8608|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|8595,8608|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Hospital Course|8595,8608|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|8595,8608|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|Hospital Course|8623,8626|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|8627,8631|false|false|false|C2598155||Pain
Event|Event|Hospital Course|8627,8631|false|false|false|||Pain
Finding|Functional Concept|Hospital Course|8627,8631|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Hospital Course|8627,8631|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Drug|Organic Chemical|Hospital Course|8636,8645|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|Hospital Course|8636,8645|false|false|false|C0001927|albuterol|albuterol
Event|Event|Hospital Course|8636,8645|false|false|false|||albuterol
Drug|Organic Chemical|Hospital Course|8636,8653|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|Hospital Course|8636,8653|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|Hospital Course|8646,8653|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|Hospital Course|8646,8653|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|Hospital Course|8646,8653|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Event|Event|Hospital Course|8646,8653|false|false|false|||sulfate
Finding|Functional Concept|Hospital Course|8671,8681|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Organism Function|Hospital Course|8671,8681|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Event|Event|Hospital Course|8682,8685|false|false|false|||Q4H
Drug|Organic Chemical|Hospital Course|8690,8698|false|false|false|C1831808|apixaban|Apixaban
Drug|Pharmacologic Substance|Hospital Course|8690,8698|false|false|false|C1831808|apixaban|Apixaban
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8707,8710|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8707,8710|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8707,8710|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|8707,8710|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|8707,8710|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|8715,8722|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Hospital Course|8715,8722|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|Hospital Course|8742,8754|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|8742,8754|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|Hospital Course|8772,8781|false|false|false|C0012373|diltiazem|Diltiazem
Drug|Pharmacologic Substance|Hospital Course|8772,8781|false|false|false|C0012373|diltiazem|Diltiazem
Finding|Finding|Hospital Course|8782,8790|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|8782,8790|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Hospital Course|8791,8798|false|false|false|||Release
Finding|Functional Concept|Hospital Course|8791,8798|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|8791,8798|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8791,8798|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8809,8812|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8809,8812|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8809,8812|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|8809,8812|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|8809,8812|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|8817,8825|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|8817,8825|false|false|false|C1692318|docusate|Docusate
Event|Event|Hospital Course|8817,8825|false|false|false|||Docusate
Drug|Organic Chemical|Hospital Course|8817,8832|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|Hospital Course|8817,8832|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|Hospital Course|8826,8832|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|8826,8832|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|8826,8832|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|8826,8832|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|8826,8832|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|8826,8832|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8843,8846|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8843,8846|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8843,8846|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|8843,8846|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|8843,8846|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|8851,8862|false|false|false|C0165590|dorzolamide|Dorzolamide
Drug|Pharmacologic Substance|Hospital Course|8851,8862|false|false|false|C0165590|dorzolamide|Dorzolamide
Finding|Functional Concept|Hospital Course|8866,8871|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|Hospital Course|8881,8885|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|Hospital Course|8881,8885|false|false|false|C1705648|Dropping|DROP
Event|Event|Hospital Course|8881,8885|false|false|false|||DROP
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8886,8895|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8891,8895|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|Hospital Course|8891,8895|false|false|false|C5848506||EYES
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8896,8899|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8896,8899|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8896,8899|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|8896,8899|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|8896,8899|false|false|false|C1332410|BID gene|BID
Drug|Element, Ion, or Isotope|Hospital Course|8904,8911|false|false|false|C2346592|Ferrous|Ferrous
Drug|Inorganic Chemical|Hospital Course|8904,8919|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Pharmacologic Substance|Hospital Course|8904,8919|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Element, Ion, or Isotope|Hospital Course|8912,8919|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Inorganic Chemical|Hospital Course|8912,8919|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Pharmacologic Substance|Hospital Course|8912,8919|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Event|Event|Hospital Course|8912,8919|false|false|false|||Sulfate
Drug|Organic Chemical|Hospital Course|8941,8952|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|8941,8952|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|Hospital Course|8941,8952|false|false|false|||Fluticasone
Drug|Organic Chemical|Hospital Course|8941,8963|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|Hospital Course|8941,8963|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|Hospital Course|8953,8963|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8964,8969|false|false|false|C0028429||NASAL
Drug|Biomedical or Dental Material|Hospital Course|8964,8969|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Organic Chemical|Hospital Course|8964,8969|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Pharmacologic Substance|Hospital Course|8964,8969|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Finding|Finding|Hospital Course|8964,8969|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Finding|Functional Concept|Hospital Course|8964,8969|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Event|Event|Hospital Course|8972,8976|false|false|false|||SPRY
Event|Event|Hospital Course|8980,8985|false|false|false|||DAILY
Finding|Gene or Genome|Hospital Course|8986,8989|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|8990,8999|false|false|false|C1717415||allergies
Event|Event|Hospital Course|8990,8999|false|false|false|||allergies
Finding|Pathologic Function|Hospital Course|8990,8999|false|false|false|C0020517|Hypersensitivity|allergies
Drug|Organic Chemical|Hospital Course|9005,9016|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|9005,9016|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|9005,9027|false|false|false|C0939232|fluticasone / salmeterol|Fluticasone-Salmeterol
Drug|Organic Chemical|Hospital Course|9005,9034|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Pharmacologic Substance|Hospital Course|9005,9034|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Organic Chemical|Hospital Course|9017,9027|false|false|false|C0073992|salmeterol|Salmeterol
Drug|Pharmacologic Substance|Hospital Course|9017,9027|false|false|false|C0073992|salmeterol|Salmeterol
Event|Event|Hospital Course|9028,9034|false|false|false|||Diskus
Drug|Biomedical or Dental Material|Hospital Course|9047,9050|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Organic Chemical|Hospital Course|9047,9050|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Pharmacologic Substance|Hospital Course|9047,9050|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Event|Event|Hospital Course|9047,9050|false|false|false|||INH
Finding|Functional Concept|Hospital Course|9047,9050|false|false|false|C0205535|Inhalation Route of Administration|INH
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9054,9057|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9054,9057|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9054,9057|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|9054,9057|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|9054,9057|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|9063,9074|false|false|false|C0018305|guaifenesin|Guaifenesin
Drug|Pharmacologic Substance|Hospital Course|9063,9074|false|false|false|C0018305|guaifenesin|Guaifenesin
Finding|Gene or Genome|Hospital Course|9089,9092|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|Hospital Course|9093,9098|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|Hospital Course|9093,9098|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|Hospital Course|9093,9098|false|false|false|||cough
Finding|Sign or Symptom|Hospital Course|9093,9098|false|false|false|C0010200|Coughing|cough
Drug|Organic Chemical|Hospital Course|9104,9123|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Pharmacologic Substance|Hospital Course|9104,9123|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Organic Chemical|Hospital Course|9144,9154|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|Hospital Course|9144,9154|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|Hospital Course|9144,9166|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|Hospital Course|9144,9166|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Event|Event|Hospital Course|9155,9166|false|false|false|||Mononitrate
Finding|Finding|Hospital Course|9168,9176|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|9168,9176|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Hospital Course|9177,9184|false|false|false|||Release
Finding|Functional Concept|Hospital Course|9177,9184|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|9177,9184|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9177,9184|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Hospital Course|9207,9218|false|false|false|C0090306|latanoprost|Latanoprost
Drug|Pharmacologic Substance|Hospital Course|9207,9218|false|false|false|C0090306|latanoprost|Latanoprost
Finding|Functional Concept|Hospital Course|9226,9231|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|Hospital Course|9241,9245|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|Hospital Course|9241,9245|false|false|false|C1705648|Dropping|DROP
Event|Event|Hospital Course|9241,9245|false|false|false|||DROP
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9246,9255|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9251,9255|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|Hospital Course|9251,9255|false|false|false|C5848506||EYES
Drug|Organic Chemical|Hospital Course|9265,9274|false|false|false|C0024002|lorazepam|Lorazepam
Drug|Pharmacologic Substance|Hospital Course|9265,9274|false|false|false|C0024002|lorazepam|Lorazepam
Finding|Gene or Genome|Hospital Course|9289,9292|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Pharmacologic Substance|Hospital Course|9293,9301|false|false|false|C1950154|Insomnia homeopathic medication|Insomnia
Event|Event|Hospital Course|9293,9301|false|false|false|||Insomnia
Finding|Sign or Symptom|Hospital Course|9293,9301|false|false|false|C0917801|Sleeplessness|Insomnia
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9303,9310|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|Hospital Course|9303,9310|false|false|false|||anxiety
Finding|Sign or Symptom|Hospital Course|9303,9310|false|false|false|C0860603|Anxiety symptoms|anxiety
Disorder|Disease or Syndrome|Hospital Course|9312,9319|false|false|false|C1135208|Vertigo as late effect of cerebrovascular disease|vertigo
Event|Event|Hospital Course|9312,9319|false|false|false|||vertigo
Finding|Sign or Symptom|Hospital Course|9312,9319|false|false|false|C0042571|Vertigo|vertigo
Drug|Organic Chemical|Hospital Course|9325,9338|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|Hospital Course|9325,9338|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|Hospital Course|9325,9338|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Event|Event|Hospital Course|9325,9338|false|false|false|||Multivitamins
Drug|Biomedical or Dental Material|Hospital Course|9341,9344|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|Hospital Course|9341,9344|false|false|false|||TAB
Drug|Hormone|Hospital Course|9359,9369|false|false|false|C0032952|prednisone|PredniSONE
Drug|Organic Chemical|Hospital Course|9359,9369|false|false|false|C0032952|prednisone|PredniSONE
Drug|Pharmacologic Substance|Hospital Course|9359,9369|false|false|false|C0032952|prednisone|PredniSONE
Procedure|Health Care Activity|Hospital Course|9386,9393|false|false|false|C0441640||Tapered
Event|Event|Hospital Course|9401,9405|false|false|false|||DOWN
Drug|Organic Chemical|Hospital Course|9411,9421|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Pharmacologic Substance|Hospital Course|9411,9421|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Organic Chemical|Hospital Course|9443,9455|false|false|false|C0039771|theophylline|Theophylline
Drug|Pharmacologic Substance|Hospital Course|9443,9455|false|false|false|C0039771|theophylline|Theophylline
Event|Event|Hospital Course|9443,9455|false|false|false|||Theophylline
Procedure|Laboratory Procedure|Hospital Course|9443,9455|false|false|false|C0039773|Assay of theophylline|Theophylline
Drug|Organic Chemical|Hospital Course|9443,9458|false|false|false|C0939729|Theophylline SR|Theophylline SR
Drug|Pharmacologic Substance|Hospital Course|9443,9458|false|false|false|C0939729|Theophylline SR|Theophylline SR
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9469,9472|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9469,9472|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9469,9472|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|9469,9472|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|9469,9472|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|9478,9488|false|false|false|C0213771|tiotropium|Tiotropium
Drug|Pharmacologic Substance|Hospital Course|9478,9488|false|false|false|C0213771|tiotropium|Tiotropium
Event|Event|Hospital Course|9478,9488|false|false|false|||Tiotropium
Drug|Organic Chemical|Hospital Course|9478,9496|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Pharmacologic Substance|Hospital Course|9478,9496|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Inorganic Chemical|Hospital Course|9489,9496|false|false|false|C0006222|Bromides|Bromide
Event|Event|Hospital Course|9489,9496|false|false|false|||Bromide
Procedure|Laboratory Procedure|Hospital Course|9489,9496|false|false|false|C0202341|Bromides measurement|Bromide
Disorder|Congenital Abnormality|Hospital Course|9499,9502|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|CAP
Drug|Biomedical or Dental Material|Hospital Course|9499,9502|false|false|false|C0006935|capsule (pharmacologic)|CAP
Event|Event|Hospital Course|9499,9502|false|false|false|||CAP
Finding|Gene or Genome|Hospital Course|9499,9502|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|CAP
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9499,9502|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|CAP
Drug|Antibiotic|Hospital Course|9517,9529|false|false|false|C0282386|levofloxacin|Levofloxacin
Drug|Organic Chemical|Hospital Course|9517,9529|false|false|false|C0282386|levofloxacin|Levofloxacin
Drug|Antibiotic|Hospital Course|9561,9573|false|false|false|C0041041|trimethoprim|Trimethoprim
Drug|Organic Chemical|Hospital Course|9561,9573|false|false|false|C0041041|trimethoprim|Trimethoprim
Drug|Biomedical or Dental Material|Hospital Course|9579,9582|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|Hospital Course|9579,9582|false|false|false|||TAB
Event|Event|Hospital Course|9592,9603|false|false|false|||prophylaxis
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9592,9603|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Finding|Idea or Concept|Hospital Course|9614,9618|false|false|false|C0233324;C1705313|Term (lexical);Term Birth|term
Finding|Organism Function|Hospital Course|9614,9618|false|false|false|C0233324;C1705313|Term (lexical);Term Birth|term
Drug|Organic Chemical|Hospital Course|9619,9626|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Drug|Pharmacologic Substance|Hospital Course|9619,9626|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Finding|Individual Behavior|Hospital Course|9619,9630|false|false|false|C0281991|Use of steroids|steroid use
Event|Event|Hospital Course|9627,9630|false|false|false|||use
Finding|Functional Concept|Hospital Course|9627,9630|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|Hospital Course|9627,9630|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Drug|Organic Chemical|Hospital Course|9636,9646|false|false|false|C3464797|Calcitrate|Calcitrate
Drug|Pharmacologic Substance|Hospital Course|9636,9646|false|false|false|C3464797|Calcitrate|Calcitrate
Drug|Organic Chemical|Hospital Course|9647,9654|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|9647,9654|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|9647,9654|false|false|false|C0042890|Vitamins|Vitamin
Event|Event|Hospital Course|9647,9654|false|false|false|||Vitamin
Drug|Hormone|Hospital Course|9647,9656|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|Hospital Course|9647,9656|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|Hospital Course|9647,9656|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|Hospital Course|9647,9656|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|Hospital Course|9647,9656|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|Hospital Course|9655,9656|false|false|false|||D
Drug|Biologically Active Substance|Hospital Course|9658,9665|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Element, Ion, or Isotope|Hospital Course|9658,9665|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Inorganic Chemical|Hospital Course|9658,9665|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Pharmacologic Substance|Hospital Course|9658,9665|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Vitamin|Hospital Course|9658,9665|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Event|Event|Hospital Course|9658,9665|false|false|false|||calcium
Finding|Physiologic Function|Hospital Course|9658,9665|false|false|false|C4553026|Calcium metabolic function|calcium
Procedure|Laboratory Procedure|Hospital Course|9658,9665|false|false|false|C0201925|Calcium measurement|calcium
Drug|Organic Chemical|Hospital Course|9658,9673|false|false|false|C0108101|calcium citrate|calcium citrate
Drug|Pharmacologic Substance|Hospital Course|9658,9673|false|false|false|C0108101|calcium citrate|calcium citrate
Drug|Organic Chemical|Hospital Course|9666,9673|false|false|false|C0008857;C0376259|Citrates;citrate|citrate
Drug|Pharmacologic Substance|Hospital Course|9666,9673|false|false|false|C0008857;C0376259|Citrates;citrate|citrate
Event|Event|Hospital Course|9666,9673|false|false|false|||citrate
Procedure|Laboratory Procedure|Hospital Course|9666,9673|false|false|false|C0201956|Citrate measurement|citrate
Drug|Organic Chemical|Hospital Course|9674,9681|false|false|false|C0042890|Vitamins|vitamin
Drug|Pharmacologic Substance|Hospital Course|9674,9681|false|false|false|C0042890|Vitamins|vitamin
Drug|Vitamin|Hospital Course|9674,9681|false|false|false|C0042890|Vitamins|vitamin
Event|Event|Hospital Course|9674,9681|false|false|false|||vitamin
Drug|Organic Chemical|Hospital Course|9674,9684|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Pharmacologic Substance|Hospital Course|9674,9684|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Vitamin|Hospital Course|9674,9684|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Anatomy|Body Space or Junction|Hospital Course|9707,9711|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|9707,9711|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|9707,9711|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|9707,9711|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|Hospital Course|9712,9717|false|false|false|||DAILY
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9723,9726|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Drug|Food|Hospital Course|9723,9726|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Drug|Immunologic Factor|Hospital Course|9723,9726|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Drug|Pharmacologic Substance|Hospital Course|9723,9726|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Event|Event|Hospital Course|9723,9726|false|false|false|||cod
Finding|Finding|Hospital Course|9723,9726|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|cod
Finding|Gene or Genome|Hospital Course|9723,9726|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|cod
Finding|Pathologic Function|Hospital Course|9723,9726|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|cod
Drug|Food|Hospital Course|9723,9736|false|false|false|C0009213|cod liver oil|cod liver oil
Drug|Organic Chemical|Hospital Course|9723,9736|false|false|false|C0009213|cod liver oil|cod liver oil
Drug|Pharmacologic Substance|Hospital Course|9723,9736|false|false|false|C0009213|cod liver oil|cod liver oil
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9727,9732|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Hospital Course|9727,9732|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Hospital Course|9727,9732|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Hospital Course|9727,9732|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Hospital Course|9727,9732|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Hospital Course|9727,9732|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|Hospital Course|9727,9732|false|false|false|||liver
Finding|Finding|Hospital Course|9727,9732|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Hospital Course|9727,9732|false|false|false|C0872387|Procedures on liver|liver
Drug|Biomedical or Dental Material|Hospital Course|9733,9736|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Food|Hospital Course|9733,9736|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Organic Chemical|Hospital Course|9733,9736|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Pharmacologic Substance|Hospital Course|9733,9736|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Event|Event|Hospital Course|9733,9736|false|false|false|||oil
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9739,9746|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|Hospital Course|9739,9746|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|Hospital Course|9739,9746|false|false|false|C0006935|capsule (pharmacologic)|capsule
Anatomy|Body Space or Junction|Hospital Course|9748,9752|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|9748,9752|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|9748,9752|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|9748,9752|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9753,9756|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9753,9756|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9753,9756|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|9753,9756|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|9753,9756|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|9762,9773|false|false|false|C0027235|ipratropium|Ipratropium
Drug|Pharmacologic Substance|Hospital Course|9762,9773|false|false|false|C0027235|ipratropium|Ipratropium
Event|Event|Hospital Course|9762,9773|false|false|false|||Ipratropium
Drug|Organic Chemical|Hospital Course|9762,9781|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Pharmacologic Substance|Hospital Course|9762,9781|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Inorganic Chemical|Hospital Course|9774,9781|false|false|false|C0006222|Bromides|Bromide
Event|Event|Hospital Course|9774,9781|false|false|false|||Bromide
Procedure|Laboratory Procedure|Hospital Course|9774,9781|false|false|false|C0202341|Bromides measurement|Bromide
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9782,9785|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|Hospital Course|9782,9785|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|Hospital Course|9782,9785|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Event|Event|Hospital Course|9782,9785|false|false|false|||Neb
Finding|Cell Function|Hospital Course|9782,9785|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|Hospital Course|9782,9785|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9788,9791|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|Hospital Course|9788,9791|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|Hospital Course|9788,9791|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|Hospital Course|9788,9791|false|false|false|||NEB
Finding|Cell Function|Hospital Course|9788,9791|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|9788,9791|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|9799,9802|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|9803,9811|false|false|false|||Wheezing
Finding|Sign or Symptom|Hospital Course|9803,9811|false|false|false|C0043144|Wheezing|Wheezing
Event|Event|Hospital Course|9816,9825|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|9816,9825|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|9816,9825|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|9816,9825|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|9816,9825|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|9816,9837|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|9826,9837|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|9826,9837|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|9826,9837|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|9826,9837|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|9842,9855|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|9842,9855|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Hospital Course|9842,9855|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|9842,9855|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|Hospital Course|9870,9873|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|9874,9878|false|false|false|C2598155||Pain
Event|Event|Hospital Course|9874,9878|false|false|false|||Pain
Finding|Functional Concept|Hospital Course|9874,9878|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Hospital Course|9874,9878|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Drug|Organic Chemical|Hospital Course|9883,9893|false|false|false|C3464797|Calcitrate|Calcitrate
Drug|Pharmacologic Substance|Hospital Course|9883,9893|false|false|false|C3464797|Calcitrate|Calcitrate
Drug|Organic Chemical|Hospital Course|9894,9901|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|9894,9901|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|9894,9901|false|false|false|C0042890|Vitamins|Vitamin
Event|Event|Hospital Course|9894,9901|false|false|false|||Vitamin
Drug|Hormone|Hospital Course|9894,9903|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|Hospital Course|9894,9903|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|Hospital Course|9894,9903|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|Hospital Course|9894,9903|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|Hospital Course|9894,9903|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|Hospital Course|9902,9903|false|false|false|||D
Drug|Biologically Active Substance|Hospital Course|9905,9912|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Element, Ion, or Isotope|Hospital Course|9905,9912|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Inorganic Chemical|Hospital Course|9905,9912|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Pharmacologic Substance|Hospital Course|9905,9912|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Vitamin|Hospital Course|9905,9912|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Event|Event|Hospital Course|9905,9912|false|false|false|||calcium
Finding|Physiologic Function|Hospital Course|9905,9912|false|false|false|C4553026|Calcium metabolic function|calcium
Procedure|Laboratory Procedure|Hospital Course|9905,9912|false|false|false|C0201925|Calcium measurement|calcium
Drug|Organic Chemical|Hospital Course|9905,9920|false|false|false|C0108101|calcium citrate|calcium citrate
Drug|Pharmacologic Substance|Hospital Course|9905,9920|false|false|false|C0108101|calcium citrate|calcium citrate
Drug|Organic Chemical|Hospital Course|9913,9920|false|false|false|C0008857;C0376259|Citrates;citrate|citrate
Drug|Pharmacologic Substance|Hospital Course|9913,9920|false|false|false|C0008857;C0376259|Citrates;citrate|citrate
Event|Event|Hospital Course|9913,9920|false|false|false|||citrate
Procedure|Laboratory Procedure|Hospital Course|9913,9920|false|false|false|C0201956|Citrate measurement|citrate
Drug|Organic Chemical|Hospital Course|9921,9928|false|false|false|C0042890|Vitamins|vitamin
Drug|Pharmacologic Substance|Hospital Course|9921,9928|false|false|false|C0042890|Vitamins|vitamin
Drug|Vitamin|Hospital Course|9921,9928|false|false|false|C0042890|Vitamins|vitamin
Event|Event|Hospital Course|9921,9928|false|false|false|||vitamin
Drug|Organic Chemical|Hospital Course|9921,9931|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Pharmacologic Substance|Hospital Course|9921,9931|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Vitamin|Hospital Course|9921,9931|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Anatomy|Body Space or Junction|Hospital Course|9954,9958|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|9954,9958|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|9954,9958|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|9954,9958|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|Hospital Course|9959,9964|false|false|false|||DAILY
Drug|Organic Chemical|Hospital Course|9969,9979|false|false|false|C0213771|tiotropium|Tiotropium
Drug|Pharmacologic Substance|Hospital Course|9969,9979|false|false|false|C0213771|tiotropium|Tiotropium
Event|Event|Hospital Course|9969,9979|false|false|false|||Tiotropium
Drug|Organic Chemical|Hospital Course|9969,9987|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Pharmacologic Substance|Hospital Course|9969,9987|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Inorganic Chemical|Hospital Course|9980,9987|false|false|false|C0006222|Bromides|Bromide
Event|Event|Hospital Course|9980,9987|false|false|false|||Bromide
Procedure|Laboratory Procedure|Hospital Course|9980,9987|false|false|false|C0202341|Bromides measurement|Bromide
Disorder|Congenital Abnormality|Hospital Course|9990,9993|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|CAP
Drug|Biomedical or Dental Material|Hospital Course|9990,9993|false|false|false|C0006935|capsule (pharmacologic)|CAP
Event|Event|Hospital Course|9990,9993|false|false|false|||CAP
Finding|Gene or Genome|Hospital Course|9990,9993|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|CAP
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9990,9993|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|CAP
Drug|Organic Chemical|Hospital Course|10007,10019|false|false|false|C0039771|theophylline|Theophylline
Drug|Pharmacologic Substance|Hospital Course|10007,10019|false|false|false|C0039771|theophylline|Theophylline
Event|Event|Hospital Course|10007,10019|false|false|false|||Theophylline
Procedure|Laboratory Procedure|Hospital Course|10007,10019|false|false|false|C0039773|Assay of theophylline|Theophylline
Drug|Organic Chemical|Hospital Course|10007,10022|false|false|false|C0939729|Theophylline SR|Theophylline SR
Drug|Pharmacologic Substance|Hospital Course|10007,10022|false|false|false|C0939729|Theophylline SR|Theophylline SR
Disorder|Mental or Behavioral Dysfunction|Hospital Course|10033,10036|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10033,10036|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|10033,10036|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|10033,10036|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|10033,10036|false|false|false|C1332410|BID gene|BID
Drug|Antibiotic|Hospital Course|10051,10063|false|false|false|C0041041|trimethoprim|Trimethoprim
Drug|Organic Chemical|Hospital Course|10051,10063|false|false|false|C0041041|trimethoprim|Trimethoprim
Drug|Biomedical or Dental Material|Hospital Course|10069,10072|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|Hospital Course|10069,10072|false|false|false|||TAB
Event|Event|Hospital Course|10082,10093|false|false|false|||prophylaxis
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10082,10093|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Finding|Idea or Concept|Hospital Course|10104,10108|false|false|false|C0233324;C1705313|Term (lexical);Term Birth|term
Finding|Organism Function|Hospital Course|10104,10108|false|false|false|C0233324;C1705313|Term (lexical);Term Birth|term
Drug|Organic Chemical|Hospital Course|10109,10116|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Drug|Pharmacologic Substance|Hospital Course|10109,10116|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Finding|Individual Behavior|Hospital Course|10109,10120|false|false|false|C0281991|Use of steroids|steroid use
Event|Event|Hospital Course|10117,10120|false|false|false|||use
Finding|Functional Concept|Hospital Course|10117,10120|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|Hospital Course|10117,10120|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Drug|Organic Chemical|Hospital Course|10125,10135|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Pharmacologic Substance|Hospital Course|10125,10135|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Hormone|Hospital Course|10156,10166|false|false|false|C0032952|prednisone|PredniSONE
Drug|Organic Chemical|Hospital Course|10156,10166|false|false|false|C0032952|prednisone|PredniSONE
Drug|Pharmacologic Substance|Hospital Course|10156,10166|false|false|false|C0032952|prednisone|PredniSONE
Drug|Organic Chemical|Hospital Course|10186,10195|false|false|false|C0024002|lorazepam|Lorazepam
Drug|Pharmacologic Substance|Hospital Course|10186,10195|false|false|false|C0024002|lorazepam|Lorazepam
Finding|Gene or Genome|Hospital Course|10210,10213|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Pharmacologic Substance|Hospital Course|10214,10222|false|false|false|C1950154|Insomnia homeopathic medication|Insomnia
Event|Event|Hospital Course|10214,10222|false|false|false|||Insomnia
Finding|Sign or Symptom|Hospital Course|10214,10222|false|false|false|C0917801|Sleeplessness|Insomnia
Disorder|Mental or Behavioral Dysfunction|Hospital Course|10224,10231|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|Hospital Course|10224,10231|false|false|false|||anxiety
Finding|Sign or Symptom|Hospital Course|10224,10231|false|false|false|C0860603|Anxiety symptoms|anxiety
Disorder|Disease or Syndrome|Hospital Course|10233,10240|false|false|false|C1135208|Vertigo as late effect of cerebrovascular disease|vertigo
Event|Event|Hospital Course|10233,10240|false|false|false|||vertigo
Finding|Sign or Symptom|Hospital Course|10233,10240|false|false|false|C0042571|Vertigo|vertigo
Drug|Organic Chemical|Hospital Course|10245,10256|false|false|false|C0090306|latanoprost|Latanoprost
Drug|Pharmacologic Substance|Hospital Course|10245,10256|false|false|false|C0090306|latanoprost|Latanoprost
Finding|Functional Concept|Hospital Course|10264,10269|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|Hospital Course|10279,10283|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|Hospital Course|10279,10283|false|false|false|C1705648|Dropping|DROP
Event|Event|Hospital Course|10279,10283|false|false|false|||DROP
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10284,10293|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10289,10293|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|Hospital Course|10289,10293|false|false|false|C5848506||EYES
Drug|Organic Chemical|Hospital Course|10303,10313|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|Hospital Course|10303,10313|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|Hospital Course|10303,10325|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|Hospital Course|10303,10325|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Event|Event|Hospital Course|10314,10325|false|false|false|||Mononitrate
Finding|Finding|Hospital Course|10327,10335|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|10327,10335|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Hospital Course|10336,10343|false|false|false|||Release
Finding|Functional Concept|Hospital Course|10336,10343|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|10336,10343|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10336,10343|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Hospital Course|10366,10377|false|false|false|C0027235|ipratropium|Ipratropium
Drug|Pharmacologic Substance|Hospital Course|10366,10377|false|false|false|C0027235|ipratropium|Ipratropium
Event|Event|Hospital Course|10366,10377|false|false|false|||Ipratropium
Drug|Organic Chemical|Hospital Course|10366,10385|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Pharmacologic Substance|Hospital Course|10366,10385|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Inorganic Chemical|Hospital Course|10378,10385|false|false|false|C0006222|Bromides|Bromide
Event|Event|Hospital Course|10378,10385|false|false|false|||Bromide
Procedure|Laboratory Procedure|Hospital Course|10378,10385|false|false|false|C0202341|Bromides measurement|Bromide
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10386,10389|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|Hospital Course|10386,10389|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|Hospital Course|10386,10389|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Event|Event|Hospital Course|10386,10389|false|false|false|||Neb
Finding|Cell Function|Hospital Course|10386,10389|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|Hospital Course|10386,10389|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10392,10395|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|Hospital Course|10392,10395|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|Hospital Course|10392,10395|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|Hospital Course|10392,10395|false|false|false|||NEB
Finding|Cell Function|Hospital Course|10392,10395|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|10392,10395|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Event|Event|Hospital Course|10403,10411|false|false|false|||Wheezing
Finding|Sign or Symptom|Hospital Course|10403,10411|false|false|false|C0043144|Wheezing|Wheezing
Drug|Organic Chemical|Hospital Course|10417,10436|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Pharmacologic Substance|Hospital Course|10417,10436|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Organic Chemical|Hospital Course|10457,10468|false|false|false|C0018305|guaifenesin|Guaifenesin
Drug|Pharmacologic Substance|Hospital Course|10457,10468|false|false|false|C0018305|guaifenesin|Guaifenesin
Finding|Gene or Genome|Hospital Course|10483,10486|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|Hospital Course|10487,10492|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|Hospital Course|10487,10492|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|Hospital Course|10487,10492|false|false|false|||cough
Finding|Sign or Symptom|Hospital Course|10487,10492|false|false|false|C0010200|Coughing|cough
Drug|Organic Chemical|Hospital Course|10498,10509|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|10498,10509|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|10498,10520|false|false|false|C0939232|fluticasone / salmeterol|Fluticasone-Salmeterol
Drug|Organic Chemical|Hospital Course|10498,10527|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Pharmacologic Substance|Hospital Course|10498,10527|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Organic Chemical|Hospital Course|10510,10520|false|false|false|C0073992|salmeterol|Salmeterol
Drug|Pharmacologic Substance|Hospital Course|10510,10520|false|false|false|C0073992|salmeterol|Salmeterol
Event|Event|Hospital Course|10521,10527|false|false|false|||Diskus
Drug|Biomedical or Dental Material|Hospital Course|10540,10543|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Organic Chemical|Hospital Course|10540,10543|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Pharmacologic Substance|Hospital Course|10540,10543|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Event|Event|Hospital Course|10540,10543|false|false|false|||INH
Finding|Functional Concept|Hospital Course|10540,10543|false|false|false|C0205535|Inhalation Route of Administration|INH
Disorder|Mental or Behavioral Dysfunction|Hospital Course|10547,10550|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10547,10550|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|10547,10550|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|10547,10550|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|10547,10550|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|10556,10567|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|10556,10567|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|Hospital Course|10556,10567|false|false|false|||Fluticasone
Drug|Organic Chemical|Hospital Course|10556,10578|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|Hospital Course|10556,10578|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|Hospital Course|10568,10578|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10579,10584|false|false|false|C0028429||NASAL
Drug|Biomedical or Dental Material|Hospital Course|10579,10584|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Organic Chemical|Hospital Course|10579,10584|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Pharmacologic Substance|Hospital Course|10579,10584|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Finding|Finding|Hospital Course|10579,10584|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Finding|Functional Concept|Hospital Course|10579,10584|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Event|Event|Hospital Course|10587,10591|false|false|false|||SPRY
Event|Event|Hospital Course|10595,10600|false|false|false|||DAILY
Finding|Gene or Genome|Hospital Course|10601,10604|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|10605,10614|false|false|false|C1717415||allergies
Event|Event|Hospital Course|10605,10614|false|false|false|||allergies
Finding|Pathologic Function|Hospital Course|10605,10614|false|false|false|C0020517|Hypersensitivity|allergies
Drug|Element, Ion, or Isotope|Hospital Course|10620,10627|false|false|false|C2346592|Ferrous|Ferrous
Drug|Inorganic Chemical|Hospital Course|10620,10635|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Pharmacologic Substance|Hospital Course|10620,10635|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Element, Ion, or Isotope|Hospital Course|10628,10635|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Inorganic Chemical|Hospital Course|10628,10635|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Pharmacologic Substance|Hospital Course|10628,10635|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Organic Chemical|Hospital Course|10657,10668|false|false|false|C0165590|dorzolamide|Dorzolamide
Drug|Pharmacologic Substance|Hospital Course|10657,10668|false|false|false|C0165590|dorzolamide|Dorzolamide
Event|Event|Hospital Course|10672,10677|false|false|false|||Ophth
Finding|Functional Concept|Hospital Course|10672,10677|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|Hospital Course|10687,10691|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|Hospital Course|10687,10691|false|false|false|C1705648|Dropping|DROP
Event|Event|Hospital Course|10687,10691|false|false|false|||DROP
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10692,10701|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10697,10701|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|Hospital Course|10697,10701|false|false|false|C5848506||EYES
Disorder|Mental or Behavioral Dysfunction|Hospital Course|10702,10705|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10702,10705|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|10702,10705|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|10702,10705|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|10702,10705|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|10711,10720|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|Hospital Course|10711,10720|false|false|false|C0001927|albuterol|albuterol
Event|Event|Hospital Course|10711,10720|false|false|false|||albuterol
Drug|Organic Chemical|Hospital Course|10711,10728|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|Hospital Course|10711,10728|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|Hospital Course|10721,10728|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|Hospital Course|10721,10728|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|Hospital Course|10721,10728|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Event|Event|Hospital Course|10721,10728|false|false|false|||sulfate
Finding|Functional Concept|Hospital Course|10746,10756|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Organism Function|Hospital Course|10746,10756|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Event|Event|Hospital Course|10757,10760|false|false|false|||Q4H
Drug|Organic Chemical|Hospital Course|10766,10774|false|false|false|C1831808|apixaban|Apixaban
Drug|Pharmacologic Substance|Hospital Course|10766,10774|false|false|false|C1831808|apixaban|Apixaban
Disorder|Mental or Behavioral Dysfunction|Hospital Course|10783,10786|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10783,10786|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|10783,10786|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|10783,10786|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|10783,10786|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|10792,10799|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Hospital Course|10792,10799|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|Hospital Course|10820,10832|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|10820,10832|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|Hospital Course|10851,10860|false|false|false|C0012373|diltiazem|Diltiazem
Drug|Pharmacologic Substance|Hospital Course|10851,10860|false|false|false|C0012373|diltiazem|Diltiazem
Finding|Finding|Hospital Course|10861,10869|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|10861,10869|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Hospital Course|10870,10877|false|false|false|||Release
Finding|Functional Concept|Hospital Course|10870,10877|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|10870,10877|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10870,10877|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Disorder|Mental or Behavioral Dysfunction|Hospital Course|10888,10891|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10888,10891|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|10888,10891|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|10888,10891|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|10888,10891|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|10897,10905|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|10897,10905|false|false|false|C1692318|docusate|Docusate
Drug|Organic Chemical|Hospital Course|10897,10912|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|Hospital Course|10897,10912|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|Hospital Course|10906,10912|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|10906,10912|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|10906,10912|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|10906,10912|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|10906,10912|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|10906,10912|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|Hospital Course|10923,10926|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10923,10926|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|10923,10926|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|10923,10926|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|10923,10926|false|false|false|C1332410|BID gene|BID
Drug|Biologically Active Substance|Hospital Course|10932,10938|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|10932,10938|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|10932,10938|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|10932,10938|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|10932,10938|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|10932,10938|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Inorganic Chemical|Hospital Course|10932,10947|false|false|false|C0037494|sodium chloride|Sodium Chloride
Drug|Clinical Drug|Hospital Course|10932,10953|false|false|false|C3213708|Sodium Chloride Nasal Product|Sodium Chloride Nasal
Drug|Element, Ion, or Isotope|Hospital Course|10939,10947|false|false|false|C0008203;C0596019|Chlorides;chloride ion|Chloride
Event|Event|Hospital Course|10939,10947|false|false|false|||Chloride
Finding|Physiologic Function|Hospital Course|10939,10947|false|false|false|C4553021|Chloride metabolic function|Chloride
Procedure|Laboratory Procedure|Hospital Course|10939,10947|false|false|false|C0201952|Chloride measurement|Chloride
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10948,10953|false|false|false|C0028429||Nasal
Drug|Biomedical or Dental Material|Hospital Course|10948,10953|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Organic Chemical|Hospital Course|10948,10953|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Pharmacologic Substance|Hospital Course|10948,10953|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Finding|Finding|Hospital Course|10948,10953|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Functional Concept|Hospital Course|10948,10953|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Event|Event|Hospital Course|10958,10962|false|false|false|||SPRY
Finding|Gene or Genome|Hospital Course|10970,10973|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10974,10979|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|Hospital Course|10974,10979|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|Hospital Course|10974,10979|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|Hospital Course|10974,10979|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|Hospital Course|10974,10979|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|Hospital Course|10974,10979|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Sign or Symptom|Hospital Course|10974,10990|false|false|false|C0858259|Nasal discomfort|nasal discomfort
Event|Event|Hospital Course|10980,10990|false|false|false|||discomfort
Finding|Sign or Symptom|Hospital Course|10980,10990|false|false|false|C2364135|Discomfort|discomfort
Drug|Biologically Active Substance|Hospital Course|10996,11002|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|Hospital Course|10996,11002|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|Hospital Course|10996,11002|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Finding|Physiologic Function|Hospital Course|10996,11002|false|false|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|Hospital Course|10996,11002|false|false|false|C0337443|Sodium measurement|sodium
Drug|Inorganic Chemical|Hospital Course|10996,11011|false|false|false|C0037494|sodium chloride|sodium chloride
Drug|Element, Ion, or Isotope|Hospital Course|11003,11011|false|false|false|C0008203;C0596019|Chlorides;chloride ion|chloride
Event|Event|Hospital Course|11003,11011|false|false|false|||chloride
Finding|Physiologic Function|Hospital Course|11003,11011|false|false|false|C4553021|Chloride metabolic function|chloride
Procedure|Laboratory Procedure|Hospital Course|11003,11011|false|false|false|C0201952|Chloride measurement|chloride
Drug|Biomedical or Dental Material|Hospital Course|11023,11028|false|false|false|C1154182|Spray Dosage Form|spray
Event|Activity|Hospital Course|11023,11028|false|false|false|C2003858|Spray (action)|spray
Event|Event|Hospital Course|11023,11028|false|false|false|||spray
Finding|Functional Concept|Hospital Course|11023,11028|false|false|false|C4521772|Spray (administration method)|spray
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11033,11038|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|Hospital Course|11033,11038|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|Hospital Course|11033,11038|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|Hospital Course|11033,11038|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|Hospital Course|11033,11038|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|Hospital Course|11033,11038|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Sign or Symptom|Hospital Course|11033,11049|false|false|false|C0027424|Nasal congestion (finding)|nasal congestion
Event|Event|Hospital Course|11039,11049|false|false|false|||congestion
Finding|Pathologic Function|Hospital Course|11039,11049|false|false|false|C0700148|Congestion|congestion
Event|Activity|Hospital Course|11050,11054|false|false|false|C1880359|Dispense (activity)|Disp
Finding|Gene or Genome|Hospital Course|11050,11054|false|false|false|C2828567|PRSS30P gene|Disp
Drug|Biomedical or Dental Material|Hospital Course|11060,11065|false|false|false|C1154182|Spray Dosage Form|Spray
Event|Activity|Hospital Course|11060,11065|false|false|false|C2003858|Spray (action)|Spray
Finding|Functional Concept|Hospital Course|11060,11065|false|false|false|C4521772|Spray (administration method)|Spray
Event|Event|Hospital Course|11066,11073|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|11066,11073|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|11081,11089|false|false|false|C0026549|morphine|Morphine
Drug|Pharmacologic Substance|Hospital Course|11081,11089|false|false|false|C0026549|morphine|Morphine
Drug|Organic Chemical|Hospital Course|11081,11097|false|false|false|C0066814|morphine sulfate|Morphine Sulfate
Drug|Pharmacologic Substance|Hospital Course|11081,11097|false|false|false|C0066814|morphine sulfate|Morphine Sulfate
Drug|Element, Ion, or Isotope|Hospital Course|11090,11097|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Inorganic Chemical|Hospital Course|11090,11097|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Pharmacologic Substance|Hospital Course|11090,11097|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Event|Event|Hospital Course|11090,11097|false|false|false|||Sulfate
Anatomy|Body Space or Junction|Hospital Course|11099,11103|false|false|false|C0226896|Oral cavity|Oral
Drug|Biomedical or Dental Material|Hospital Course|11099,11103|false|false|false|C1272919|Oral Dosage Form|Oral
Finding|Finding|Hospital Course|11099,11103|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Finding|Functional Concept|Hospital Course|11099,11103|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Drug|Biomedical or Dental Material|Hospital Course|11099,11112|false|false|false|C0991536|Oral Solution|Oral Solution
Drug|Biomedical or Dental Material|Hospital Course|11104,11112|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|Solution
Drug|Substance|Hospital Course|11104,11112|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|Solution
Event|Event|Hospital Course|11104,11112|false|false|false|||Solution
Finding|Conceptual Entity|Hospital Course|11104,11112|false|false|false|C2699488|Resolution|Solution
Finding|Gene or Genome|Hospital Course|11134,11137|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|11139,11148|false|false|false|||shortness
Attribute|Clinical Attribute|Hospital Course|11139,11158|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|Hospital Course|11139,11158|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|Hospital Course|11152,11158|false|false|false|C0225386|Breath|breath
Drug|Organic Chemical|Hospital Course|11164,11172|false|false|false|C0026549|morphine|morphine
Drug|Pharmacologic Substance|Hospital Course|11164,11172|false|false|false|C0026549|morphine|morphine
Event|Event|Hospital Course|11164,11172|false|false|false|||morphine
Finding|Functional Concept|Hospital Course|11191,11199|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|11194,11199|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|11194,11199|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Event|Hospital Course|11222,11226|false|false|false|||Disp
Finding|Idea or Concept|Hospital Course|11253,11260|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|11268,11278|false|false|false|C0054201|budesonide|Budesonide
Drug|Pharmacologic Substance|Hospital Course|11268,11278|false|false|false|C0054201|budesonide|Budesonide
Drug|Clinical Drug|Hospital Course|11268,11284|false|false|false|C0360546;C3832695|Budesonide Nasal (Brand Name);Budesonide Nasal Product|Budesonide Nasal
Drug|Pharmacologic Substance|Hospital Course|11268,11284|false|false|false|C0360546;C3832695|Budesonide Nasal (Brand Name);Budesonide Nasal Product|Budesonide Nasal
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11279,11284|false|false|false|C0028429||Nasal
Drug|Biomedical or Dental Material|Hospital Course|11279,11284|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Organic Chemical|Hospital Course|11279,11284|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Pharmacologic Substance|Hospital Course|11279,11284|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Finding|Finding|Hospital Course|11279,11284|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Functional Concept|Hospital Course|11279,11284|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Event|Event|Hospital Course|11285,11292|false|false|false|||Inhaler
Finding|Functional Concept|Hospital Course|11285,11292|false|false|false|C4319647|Inhaler (unit of presentation)|Inhaler
Drug|Organic Chemical|Hospital Course|11318,11328|false|false|false|C0054201|budesonide|budesonide
Drug|Pharmacologic Substance|Hospital Course|11318,11328|false|false|false|C0054201|budesonide|budesonide
Event|Event|Hospital Course|11318,11328|false|false|false|||budesonide
Drug|Organic Chemical|Hospital Course|11330,11339|false|false|false|C0678162|Pulmicort|Pulmicort
Drug|Pharmacologic Substance|Hospital Course|11330,11339|false|false|false|C0678162|Pulmicort|Pulmicort
Drug|Organic Chemical|Hospital Course|11330,11349|false|false|false|C1950317|Pulmicort Flexhaler|Pulmicort Flexhaler
Drug|Pharmacologic Substance|Hospital Course|11330,11349|false|false|false|C1950317|Pulmicort Flexhaler|Pulmicort Flexhaler
Event|Event|Hospital Course|11340,11349|false|false|false|||Flexhaler
Event|Event|Hospital Course|11379,11388|false|false|false|||delivered
Drug|Biomedical or Dental Material|Hospital Course|11397,11400|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Organic Chemical|Hospital Course|11397,11400|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Pharmacologic Substance|Hospital Course|11397,11400|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Event|Event|Hospital Course|11397,11400|false|false|false|||INH
Finding|Functional Concept|Hospital Course|11397,11400|false|false|false|C0205535|Inhalation Route of Administration|INH
Event|Event|Hospital Course|11407,11411|false|false|false|||Disp
Finding|Functional Concept|Hospital Course|11416,11423|false|false|false|C4319647|Inhaler (unit of presentation)|Inhaler
Event|Event|Hospital Course|11424,11431|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|11424,11431|false|false|false|C0807726|refill|Refills
Event|Event|Hospital Course|11438,11447|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|11438,11447|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|11438,11447|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|11438,11447|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|11438,11447|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|11438,11459|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|11438,11459|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|11448,11459|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|11448,11459|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|11448,11459|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|Hospital Course|11461,11465|false|false|false|||Home
Finding|Idea or Concept|Hospital Course|11461,11465|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|11461,11465|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|11461,11465|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|Hospital Course|11471,11478|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|Hospital Course|11471,11478|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|Hospital Course|11481,11489|false|false|false|||Facility
Finding|Intellectual Product|Hospital Course|11481,11489|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|Hospital Course|11497,11506|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|11497,11506|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|11497,11506|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|11497,11506|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|11497,11506|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|11497,11516|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|11507,11516|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|11507,11516|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|11507,11516|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|11507,11516|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|11507,11516|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Finding|Principle Diagnosis|11537,11543|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Finding|Intellectual Product|Principle Diagnosis|11537,11543|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Disorder|Disease or Syndrome|Principle Diagnosis|11544,11548|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Principle Diagnosis|11544,11548|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Principle Diagnosis|11544,11548|false|false|false|||COPD
Finding|Gene or Genome|Principle Diagnosis|11544,11548|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Neoplastic Process|Principle Diagnosis|11550,11559|false|false|false|C0027627|Neoplasm Metastasis|SECONDARY
Finding|Functional Concept|Principle Diagnosis|11550,11559|false|false|false|C1522484|metastatic qualifier|SECONDARY
Event|Event|Principle Diagnosis|11560,11569|false|false|false|||DIAGNOSES
Procedure|Diagnostic Procedure|Principle Diagnosis|11560,11569|false|false|false|C0011900|Diagnosis|DIAGNOSES
Disorder|Disease or Syndrome|Principle Diagnosis|11571,11574|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Principle Diagnosis|11571,11574|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Principle Diagnosis|11571,11574|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Principle Diagnosis|11571,11574|false|false|false|||CAD
Finding|Gene or Genome|Principle Diagnosis|11571,11574|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Principle Diagnosis|11571,11574|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Principle Diagnosis|11571,11574|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Principle Diagnosis|11571,11574|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|Principle Diagnosis|11575,11587|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|Principle Diagnosis|11575,11587|false|false|false|||Hypertension
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|11588,11594|false|false|false|C0018792|Heart Atrium|Atrial
Attribute|Clinical Attribute|Principle Diagnosis|11588,11607|false|false|false|C2926591||Atrial fibrillation
Disorder|Disease or Syndrome|Principle Diagnosis|11588,11607|false|false|false|C0004238|Atrial Fibrillation|Atrial fibrillation
Lab|Laboratory or Test Result|Principle Diagnosis|11588,11607|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Atrial fibrillation
Disorder|Disease or Syndrome|Principle Diagnosis|11595,11607|false|false|false|C0232197|Fibrillation|fibrillation
Event|Event|Principle Diagnosis|11595,11607|false|false|false|||fibrillation
Finding|Mental Process|Discharge Condition|11632,11638|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|11632,11645|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|11632,11645|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|11639,11645|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|11639,11645|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|11647,11652|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|11647,11652|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|11657,11665|false|false|false|||coherent
Finding|Finding|Discharge Condition|11657,11665|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|11667,11672|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|11667,11689|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|11667,11689|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|11676,11689|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|11676,11689|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|11676,11689|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|11691,11696|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|11691,11696|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|11691,11696|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|11691,11696|false|false|false|||Alert
Finding|Finding|Discharge Condition|11691,11696|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|11691,11696|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|11691,11696|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|11701,11712|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|11701,11712|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|11714,11722|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|11714,11722|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|11714,11722|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|11723,11729|false|false|false|C5889824||Status
Event|Event|Discharge Condition|11723,11729|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|11723,11729|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|11731,11741|false|false|false|||Ambulatory
Finding|Functional Concept|Discharge Condition|11731,11741|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|11731,11741|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|11731,11741|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|11731,11741|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|11744,11755|false|false|false|||Independent
Finding|Finding|Discharge Condition|11744,11755|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Condition|11744,11755|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Gene or Genome|Discharge Instructions|11784,11788|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Finding|Gene or Genome|Discharge Instructions|11805,11810|false|false|false|C1424898|RXFP2 gene|great
Event|Event|Discharge Instructions|11811,11819|false|false|false|||pleasure
Finding|Intellectual Product|Discharge Instructions|11811,11819|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|Discharge Instructions|11811,11819|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|Discharge Instructions|11827,11831|false|false|false|C1947933|care activity|care
Event|Event|Discharge Instructions|11827,11831|false|false|false|||care
Finding|Finding|Discharge Instructions|11827,11831|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|11827,11831|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|11827,11834|false|false|false|C1555558|care of - AddressPartType|care of
Event|Event|Discharge Instructions|11856,11860|false|false|false|||came
Finding|Idea or Concept|Discharge Instructions|11868,11876|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|Discharge Instructions|11895,11907|false|false|false|||experiencing
Event|Event|Discharge Instructions|11918,11927|false|false|false|||shortness
Attribute|Clinical Attribute|Discharge Instructions|11918,11937|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|Discharge Instructions|11918,11937|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|Discharge Instructions|11931,11937|false|false|false|C0225386|Breath|breath
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|11939,11948|false|false|false|C0024109|Lung|Pulmonary
Attribute|Clinical Attribute|Discharge Instructions|11939,11948|false|false|false|C2707265||Pulmonary
Finding|Finding|Discharge Instructions|11939,11948|false|false|false|C4522268|Pulmonary (intended site)|Pulmonary
Event|Event|Discharge Instructions|11955,11958|false|false|false|||saw
Event|Event|Discharge Instructions|11967,11975|false|false|false|||reviewed
Attribute|Clinical Attribute|Discharge Instructions|11981,11990|false|false|false|C3864998||condition
Disorder|Disease or Syndrome|Discharge Instructions|11981,11990|false|false|false|C0012634|Disease|condition
Event|Event|Discharge Instructions|11981,11990|false|false|false|||condition
Finding|Conceptual Entity|Discharge Instructions|11981,11990|false|false|false|C1705253|Logical Condition|condition
Event|Event|Discharge Instructions|12001,12009|false|false|false|||symptoms
Finding|Functional Concept|Discharge Instructions|12001,12009|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Discharge Instructions|12001,12009|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|Discharge Instructions|12015,12022|false|false|false|||thought
Finding|Idea or Concept|Discharge Instructions|12015,12022|false|false|false|C0039869;C4319827|Thought|thought
Finding|Mental Process|Discharge Instructions|12015,12022|false|false|false|C0039869;C4319827|Thought|thought
Drug|Organic Chemical|Discharge Instructions|12029,12036|false|false|false|C0163712|Relate - vinyl resin|related
Event|Event|Discharge Instructions|12029,12036|false|false|false|||related
Finding|Finding|Discharge Instructions|12029,12036|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|Discharge Instructions|12029,12036|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Event|Event|Discharge Instructions|12040,12046|false|false|false|||severe
Finding|Finding|Discharge Instructions|12040,12046|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Discharge Instructions|12040,12046|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|Discharge Instructions|12047,12051|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Discharge Instructions|12047,12051|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Discharge Instructions|12047,12051|false|false|false|||COPD
Finding|Gene or Genome|Discharge Instructions|12047,12051|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|Discharge Instructions|12065,12072|false|false|false|||changes
Finding|Functional Concept|Discharge Instructions|12065,12072|false|false|false|C0392747|Changing|changes
Attribute|Clinical Attribute|Discharge Instructions|12082,12093|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|12082,12093|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|12082,12093|false|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|12082,12093|false|false|false|C4284232|Medications|medications
Event|Event|Discharge Instructions|12098,12107|false|false|false|||increased
Drug|Hormone|Discharge Instructions|12120,12130|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|Discharge Instructions|12120,12130|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|Discharge Instructions|12120,12130|false|false|false|C0032952|prednisone|prednisone
Event|Event|Discharge Instructions|12120,12130|false|false|false|||prednisone
Finding|Finding|Discharge Instructions|12137,12152|false|false|false|C0700049|Encounter due to palliative care|Palliative Care
Procedure|Health Care Activity|Discharge Instructions|12137,12152|false|false|false|C0030231;C3816218|Palliative Care;Palliative Nursing|Palliative Care
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|12137,12152|false|false|false|C0030231;C3816218|Palliative Care;Palliative Nursing|Palliative Care
Event|Activity|Discharge Instructions|12148,12152|false|false|false|C1947933|care activity|Care
Finding|Finding|Discharge Instructions|12148,12152|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Discharge Instructions|12148,12152|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Attribute|Clinical Attribute|Discharge Instructions|12148,12157|false|false|false|C4321316||Care team
Finding|Finding|Discharge Instructions|12148,12157|false|false|false|C4321315|Care team|Care team
Event|Event|Discharge Instructions|12153,12157|false|false|false|||team
Event|Event|Discharge Instructions|12162,12171|false|false|false|||consulted
Event|Event|Discharge Instructions|12176,12183|false|false|false|||started
Drug|Organic Chemical|Discharge Instructions|12191,12199|false|false|false|C0026549|morphine|morphine
Drug|Pharmacologic Substance|Discharge Instructions|12191,12199|false|false|false|C0026549|morphine|morphine
Event|Event|Discharge Instructions|12191,12199|false|false|false|||morphine
Drug|Biomedical or Dental Material|Discharge Instructions|12201,12207|false|false|false|C0302908;C1697794|Liquid Dosage Form;Liquid substance|liquid
Drug|Substance|Discharge Instructions|12201,12207|false|false|false|C0302908;C1697794|Liquid Dosage Form;Liquid substance|liquid
Event|Event|Discharge Instructions|12201,12207|false|false|false|||liquid
Finding|Finding|Discharge Instructions|12201,12207|false|false|false|C1304698|Liquid (finding)|liquid
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|12201,12207|false|false|false|C0301571|Liquid diet|liquid
Drug|Biomedical or Dental Material|Discharge Instructions|12208,12218|false|false|false|C0038960;C1382107|Suspension substance;Suspensions|suspension
Drug|Substance|Discharge Instructions|12208,12218|false|false|false|C0038960;C1382107|Suspension substance;Suspensions|suspension
Event|Event|Discharge Instructions|12208,12218|false|false|false|||suspension
Finding|Functional Concept|Discharge Instructions|12208,12218|false|false|false|C1705537|Suspension (action)|suspension
Event|Event|Discharge Instructions|12222,12226|false|false|false|||help
Attribute|Clinical Attribute|Discharge Instructions|12237,12246|false|false|false|C5885990||breathing
Finding|Finding|Discharge Instructions|12237,12246|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|Discharge Instructions|12237,12246|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|Discharge Instructions|12237,12246|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|Discharge Instructions|12237,12246|false|false|false|C1160636|respiratory system process|breathing
Finding|Sign or Symptom|Discharge Instructions|12237,12255|false|false|false|C0424805|breath symptom|breathing symptoms
Event|Event|Discharge Instructions|12247,12255|false|false|false|||symptoms
Finding|Functional Concept|Discharge Instructions|12247,12255|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Discharge Instructions|12247,12255|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Attribute|Clinical Attribute|Discharge Instructions|12279,12290|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|12279,12290|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|12279,12290|false|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|12279,12290|false|false|false|C4284232|Medications|medications
Finding|Finding|Discharge Instructions|12294,12298|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Discharge Instructions|12294,12298|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Discharge Instructions|12294,12298|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|Discharge Instructions|12303,12309|false|false|false|||follow
Event|Event|Discharge Instructions|12324,12331|false|false|false|||doctors
Procedure|Health Care Activity|Discharge Instructions|12371,12379|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|12380,12392|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|12380,12392|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|12380,12392|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

