 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Procedure|Health Care Activity|SIMPLE_SEGMENT|47,56|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|47,61|false|false|false|C2598112||Admission Date
Finding|Body Substance|SIMPLE_SEGMENT|81,90|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|81,90|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|81,90|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|81,90|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|81,95|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|113,118|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|113,118|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|113,118|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|137,140|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|137,140|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|137,140|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|137,140|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|137,140|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|148,155|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|148,155|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Finding|Finding|SIMPLE_SEGMENT|157,164|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Finding|Functional Concept|SIMPLE_SEGMENT|157,164|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Finding|Idea or Concept|SIMPLE_SEGMENT|157,164|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|157,164|false|false|false|C0543467|Operative Surgical Procedures|SURGERY
Attribute|Clinical Attribute|SIMPLE_SEGMENT|167,176|false|false|false|C1717415||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|167,176|false|false|false|C0020517|Hypersensitivity|Allergies
Attribute|Clinical Attribute|SIMPLE_SEGMENT|188,197|false|false|false|C1717415||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|188,197|false|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|200,222|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|208,212|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|SIMPLE_SEGMENT|208,212|false|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|SIMPLE_SEGMENT|208,222|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Finding|Functional Concept|SIMPLE_SEGMENT|225,234|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|243,258|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|249,258|false|false|false|C3864418||Complaint
Finding|Finding|SIMPLE_SEGMENT|249,258|false|false|false|C5441521|Complaint (finding)|Complaint
Disorder|Neoplastic Process|SIMPLE_SEGMENT|260,294|false|false|false|C5206813|Locally Advanced Gastric Carcinoma|Locally advanced gastric carcinoma
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|277,284|false|false|false|C0038351|Stomach|gastric
Disorder|Neoplastic Process|SIMPLE_SEGMENT|277,294|false|false|false|C0699791|Stomach Carcinoma|gastric carcinoma
Disorder|Neoplastic Process|SIMPLE_SEGMENT|285,294|false|false|false|C0007097|Carcinoma|carcinoma
Finding|Classification|SIMPLE_SEGMENT|297,302|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|303,311|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|303,311|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|315,333|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|324,333|false|false|false|C0945766||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|324,333|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|324,333|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|324,333|false|false|false|C0184661|Interventional procedure|Procedure
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|335,345|false|false|false|C0010702|Cystoscopy|Cystoscopy
Finding|Intellectual Product|SIMPLE_SEGMENT|356,364|false|true|false|C1546572||catheter
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|356,374|false|true|false|C0883301|Catheter placement|catheter placement
Procedure|Health Care Activity|SIMPLE_SEGMENT|365,374|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|365,374|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|376,387|false|false|false|C0031150;C1883297|Laparoscopy;Therapeutic Laparoscopy|Laparoscopy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|376,387|false|false|false|C0031150;C1883297|Laparoscopy;Therapeutic Laparoscopy|Laparoscopy
Finding|Finding|SIMPLE_SEGMENT|394,400|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Finding|Intellectual Product|SIMPLE_SEGMENT|394,400|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|394,400|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Procedure|Health Care Activity|SIMPLE_SEGMENT|394,400|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|402,413|false|false|false|C0017195|Endoscopy of stomach|Gastroscopy
Finding|Conceptual Entity|SIMPLE_SEGMENT|417,424|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|417,424|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|417,424|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|417,427|false|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|417,443|false|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|417,443|false|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|428,435|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|428,435|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|428,443|false|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|436,443|false|false|false|C0221423|Illness (finding)|Illness
Finding|Idea or Concept|SIMPLE_SEGMENT|462,466|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|SIMPLE_SEGMENT|462,466|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Finding|SIMPLE_SEGMENT|471,475|false|false|false|C1706180|Male Gender|male
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|498,505|false|false|false|C0038351|Stomach|gastric
Disorder|Neoplastic Process|SIMPLE_SEGMENT|507,513|false|false|false|C0006826|Malignant Neoplasms|cancer
Attribute|Clinical Attribute|SIMPLE_SEGMENT|515,520|false|false|false|C1300072|Tumor stage|stage
Finding|Conceptual Entity|SIMPLE_SEGMENT|556,564|false|false|false|C1880198|Cure (remedy)|curative
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|556,564|false|false|false|C1276305|Curative - procedure intent|curative
Finding|Idea or Concept|SIMPLE_SEGMENT|565,571|false|false|false|C0162425;C1550453|Act Mood - intent|intent
Finding|Mental Process|SIMPLE_SEGMENT|565,571|false|false|false|C0162425;C1550453|Act Mood - intent|intent
Procedure|Health Care Activity|SIMPLE_SEGMENT|572,580|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|572,580|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|572,590|false|false|false|C0015252;C0728940|Excision;removal technique|surgical resection
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|581,590|false|false|false|C0015252;C0728940|Excision;removal technique|resection
Finding|Functional Concept|SIMPLE_SEGMENT|611,620|false|false|false|C0205263|Induce (action)|induction
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|611,620|false|false|false|C0857127|Induction procedure|induction
Finding|Functional Concept|SIMPLE_SEGMENT|622,634|false|false|false|C0013217|pharmacotherapeutic|chemotherapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|622,634|false|false|false|C0013216;C0392920;C3665472|Chemotherapy;Chemotherapy Regimen;Pharmacotherapy|chemotherapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|656,667|false|false|false|C0600558|Neoadjuvant Therapy|neoadjuvant
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|656,680|false|false|false|C5392214|Neoadjuvant Chemotherapy|neoadjuvant chemotherapy
Finding|Functional Concept|SIMPLE_SEGMENT|668,680|false|false|false|C0013217|pharmacotherapeutic|chemotherapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|668,680|false|false|false|C0013216;C0392920;C3665472|Chemotherapy;Chemotherapy Regimen;Pharmacotherapy|chemotherapy
Finding|Intellectual Product|SIMPLE_SEGMENT|700,707|false|false|false|C0282416|Overall Publication Type|Overall
Finding|Functional Concept|SIMPLE_SEGMENT|725,737|false|false|false|C0013217|pharmacotherapeutic|chemotherapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|725,737|false|false|false|C0013216;C0392920;C3665472|Chemotherapy;Chemotherapy Regimen;Pharmacotherapy|chemotherapy
Finding|Finding|SIMPLE_SEGMENT|738,742|false|false|false|C5575035|Well (answer to question)|well
Finding|Idea or Concept|SIMPLE_SEGMENT|756,767|false|false|false|C0750502|Significant|significant
Finding|Functional Concept|SIMPLE_SEGMENT|768,780|false|false|false|C0001688;C0879626|Adverse effects;aspects of adverse effects|side effects
Finding|Pathologic Function|SIMPLE_SEGMENT|768,780|false|false|false|C0001688;C0879626|Adverse effects;aspects of adverse effects|side effects
Finding|Idea or Concept|SIMPLE_SEGMENT|796,801|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|SIMPLE_SEGMENT|796,801|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Functional Concept|SIMPLE_SEGMENT|815,820|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|815,836|false|false|false|C0230329|Right upper extremity|right upper extremity
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|821,836|false|false|false|C1140618|Upper Extremity|upper extremity
Finding|Pathologic Function|SIMPLE_SEGMENT|821,842|false|false|false|C0522035|Edema of the upper extremity|upper extremity edema
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|827,836|false|false|false|C0015385|Limb structure|extremity
Finding|Pathologic Function|SIMPLE_SEGMENT|827,842|false|false|false|C0085649|Peripheral edema|extremity edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|837,842|false|false|false|C1717255||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|837,842|false|false|false|C0013604|Edema|edema
Finding|Pathologic Function|SIMPLE_SEGMENT|867,877|false|false|false|C0040053|Thrombosis|thrombosis
Drug|Organic Chemical|SIMPLE_SEGMENT|910,917|false|false|false|C0728963|Lovenox|Lovenox
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|910,917|false|false|false|C0728963|Lovenox|Lovenox
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|927,930|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|927,930|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|927,930|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|927,930|false|false|false|C1332410|BID gene|BID
Finding|Individual Behavior|SIMPLE_SEGMENT|944,953|false|false|false|C1321605|Compliance behavior|compliant
Finding|Finding|SIMPLE_SEGMENT|971,976|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|971,976|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Attribute|Clinical Attribute|SIMPLE_SEGMENT|978,984|true|false|false|C4255480||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|978,984|true|false|false|C0027497|Nausea|nausea
Finding|Body Substance|SIMPLE_SEGMENT|986,992|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Physiologic Function|SIMPLE_SEGMENT|986,992|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Sign or Symptom|SIMPLE_SEGMENT|986,992|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Sign or Symptom|SIMPLE_SEGMENT|994,1000|false|false|false|C0085593|Chills|chills
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1002,1008|false|false|false|C0944911||weight
Finding|Finding|SIMPLE_SEGMENT|1002,1008|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|1002,1008|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|1002,1008|false|false|false|C1305866|Weighing patient|weight
Finding|Finding|SIMPLE_SEGMENT|1002,1013|false|false|false|C1262477;C3540682|Losing Weight (question);Weight Loss|weight loss
Finding|Intellectual Product|SIMPLE_SEGMENT|1002,1013|false|false|false|C1262477;C3540682|Losing Weight (question);Weight Loss|weight loss
Finding|Finding|SIMPLE_SEGMENT|1009,1013|false|false|false|C5890125|Loss (adaptation)|loss
Finding|Pathologic Function|SIMPLE_SEGMENT|1015,1021|false|false|false|C0025222|Melena|melena
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1023,1035|false|false|false|C0018932|Hematochezia|hematochezia
Finding|Sign or Symptom|SIMPLE_SEGMENT|1023,1035|false|false|false|C1321898|Blood in stool|hematochezia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1039,1048|false|false|false|C0018965|Hematuria|hematuria
Finding|Functional Concept|SIMPLE_SEGMENT|1074,1080|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Finding|Functional Concept|SIMPLE_SEGMENT|1081,1088|false|false|false|C0332305|With staging|staging
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1109,1113|false|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Finding|Idea or Concept|SIMPLE_SEGMENT|1131,1139|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|1131,1142|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1143,1150|true|false|false|C0012634|Disease|disease
Finding|Finding|SIMPLE_SEGMENT|1179,1188|false|false|false|C4738506|Operating|operating
Finding|Finding|SIMPLE_SEGMENT|1221,1229|false|false|false|C0332149|Possible|possibly
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|1235,1242|false|false|false|C0302912|Radicals (chemistry)|radical
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1243,1249|false|false|false|C4522154|Distal Resection Margin|distal
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1243,1261|false|false|false|C0176758;C0192440|Billroth I Procedure;Partial gastrectomy with anastomosis to duodenum|distal gastrectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1250,1261|false|false|false|C0017118|Gastrectomy|gastrectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1267,1282|false|false|false|C0024203|Lymph node excision|lymphadenectomy
Finding|Idea or Concept|SIMPLE_SEGMENT|1289,1294|false|false|false|C0035647|Risk|risks
Finding|Finding|SIMPLE_SEGMENT|1311,1318|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|1311,1318|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|1311,1318|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1311,1318|false|false|false|C0543467|Operative Surgical Procedures|surgery
Finding|Body Substance|SIMPLE_SEGMENT|1348,1355|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1348,1355|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1348,1355|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|SIMPLE_SEGMENT|1359,1365|false|false|false|C1561567|detail - Response Level|detail
Finding|Finding|SIMPLE_SEGMENT|1418,1438|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Finding|Functional Concept|SIMPLE_SEGMENT|1423,1430|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|1423,1430|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|1423,1430|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1423,1430|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|1423,1438|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1431,1438|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1431,1438|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1431,1438|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1440,1460|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Finding|Functional Concept|SIMPLE_SEGMENT|1445,1452|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|1445,1452|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|1445,1452|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1445,1452|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|1445,1460|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1453,1460|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1453,1460|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1453,1460|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1462,1470|false|false|false|C0033572;C4266527|Prostate;Structure of prostate (body structure)|Prostate
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1462,1470|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|Prostate
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1462,1470|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|Prostate
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1462,1477|false|false|false|C0376358;C0600139|Malignant neoplasm of prostate;Prostate carcinoma|Prostate cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1471,1477|false|false|false|C0006826|Malignant Neoplasms|cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1471,1486|false|false|false|C0549473|Thyroid carcinoma|cancer, Thyroid
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1479,1486|false|false|false|C0040132|Thyroid Gland|Thyroid
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1479,1486|false|false|false|C0040128|Thyroid Diseases|Thyroid
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1479,1486|false|false|false|C0040134;C3540038;C5781115|THYROID;THYROID DIAGNOSTIC RADIOPHARMACEUTICALS;thyroid (USP)|Thyroid
Drug|Hormone|SIMPLE_SEGMENT|1479,1486|false|false|false|C0040134;C3540038;C5781115|THYROID;THYROID DIAGNOSTIC RADIOPHARMACEUTICALS;thyroid (USP)|Thyroid
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|1479,1486|false|false|false|C0040134;C3540038;C5781115|THYROID;THYROID DIAGNOSTIC RADIOPHARMACEUTICALS;thyroid (USP)|Thyroid
Drug|Organic Chemical|SIMPLE_SEGMENT|1479,1486|false|false|false|C0040134;C3540038;C5781115|THYROID;THYROID DIAGNOSTIC RADIOPHARMACEUTICALS;thyroid (USP)|Thyroid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1479,1486|false|false|false|C0040134;C3540038;C5781115|THYROID;THYROID DIAGNOSTIC RADIOPHARMACEUTICALS;thyroid (USP)|Thyroid
Procedure|Health Care Activity|SIMPLE_SEGMENT|1479,1486|false|false|false|C2228489|examination of thyroid|Thyroid
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1479,1493|false|false|false|C0040137|Thyroid Nodule|Thyroid nodule
Finding|Finding|SIMPLE_SEGMENT|1479,1493|false|false|false|C2116082||Thyroid nodule
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1495,1506|false|false|false|C0020676|Hypothyroidism|Hypothyroid
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1508,1512|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Finding|Intellectual Product|SIMPLE_SEGMENT|1513,1517|false|false|false|C1547225|Mild Severity of Illness Code|mild
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1519,1533|false|false|false|C1510475|Diverticulosis|Diverticulosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1537,1548|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Procedure|Health Care Activity|SIMPLE_SEGMENT|1537,1548|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1553,1559|false|false|false|C0002871|Anemia|anemia
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1560,1564|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|1560,1564|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1560,1564|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1560,1564|false|false|false|C0337439|Iron measurement|iron
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|1565,1568|false|false|false|C0054282|butyl phosphorotrithioate|def
Drug|Organic Chemical|SIMPLE_SEGMENT|1565,1568|false|false|false|C0054282|butyl phosphorotrithioate|def
Finding|Gene or Genome|SIMPLE_SEGMENT|1565,1568|false|false|false|C1823727|UTP25 gene|def
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1570,1576|false|false|false|C0002871|Anemia|anemia
Finding|Finding|SIMPLE_SEGMENT|1607,1628|false|false|false|C0455610|History of surgery|Past Surgical History
Procedure|Health Care Activity|SIMPLE_SEGMENT|1612,1620|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1612,1620|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Finding|Finding|SIMPLE_SEGMENT|1612,1628|false|false|false|C0744961|history of prior surgery|Surgical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1621,1628|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1621,1628|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1621,1628|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1630,1638|false|false|false|C0033572;C4266527|Prostate;Structure of prostate (body structure)|Prostate
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1630,1638|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|Prostate
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1630,1638|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|Prostate
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1630,1645|false|false|false|C0376358;C0600139|Malignant neoplasm of prostate;Prostate carcinoma|Prostate cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1639,1645|false|false|false|C0006826|Malignant Neoplasms|cancer
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1646,1654|false|false|false|C1548801|Body Site Modifier - External|external
Finding|Functional Concept|SIMPLE_SEGMENT|1646,1654|false|false|false|C0521134|External route|external
Drug|Organic Chemical|SIMPLE_SEGMENT|1655,1659|false|false|false|C4521565|Beam -- chemical|beam
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1655,1659|false|false|false|C4521565|Beam -- chemical|beam
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|1655,1659|false|false|false|C2347880|Beam - rays of radiation or stream of particles|beam
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1655,1659|false|false|false|C0338248|carmustine/cytarabine/etoposide/melphalan regimen|beam
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1665,1673|false|false|false|C0001074|Structure of achilles tendon|Achilles
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1665,1680|false|false|false|C0001074;C1305378|Structure of achilles tendon|Achilles tendon
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1665,1687|false|false|false|C0407029|Repair of Achilles tendon|Achilles tendon repair
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1674,1680|false|false|false|C0039508|Tendon structure|tendon
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1674,1687|false|false|false|C0565350|Plastic repair of tendon|tendon repair
Finding|Functional Concept|SIMPLE_SEGMENT|1681,1687|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Finding|Organism Function|SIMPLE_SEGMENT|1681,1687|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Procedure|Health Care Activity|SIMPLE_SEGMENT|1681,1687|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1681,1687|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Finding|Functional Concept|SIMPLE_SEGMENT|1703,1708|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1703,1714|false|false|false|C0817321|Right tibia|right tibia
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1709,1714|false|false|false|C0040184|Bone structure of tibia|tibia
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1709,1725|false|false|false|C0947635|tibia and fibula|tibia and fibula
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1719,1725|false|false|false|C0016068|Fibula|fibula
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1727,1740|false|false|false|C0040423|Tonsillectomy|Tonsillectomy
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1741,1744|false|false|false|C1114365||age
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1741,1744|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|SIMPLE_SEGMENT|1741,1744|false|false|false|C0162574|Glycation End Products, Advanced|age
Finding|Functional Concept|SIMPLE_SEGMENT|1752,1758|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|1752,1766|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1759,1766|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1759,1766|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1759,1766|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|1772,1778|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|1772,1778|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|1772,1778|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|1772,1778|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|1772,1786|false|false|false|C0241889|Family Medical History|Family History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1779,1786|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1779,1786|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1779,1786|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1788,1794|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|SIMPLE_SEGMENT|1788,1794|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1812,1820|false|false|false|C0024299|Lymphoma|Lymphoma
Finding|Idea or Concept|SIMPLE_SEGMENT|1822,1828|false|false|false|C1546508|Relationship - Mother|Mother
Finding|Gene or Genome|SIMPLE_SEGMENT|1846,1850|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Intellectual Product|SIMPLE_SEGMENT|1846,1850|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1859,1867|false|false|false|C0011265;C0497327|Dementia;Presenile dementia|Dementia
Finding|Finding|SIMPLE_SEGMENT|1873,1881|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|1873,1881|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1873,1881|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|1873,1886|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1873,1886|false|false|false|C0031809|Physical Examination|Physical Exam
Finding|Functional Concept|SIMPLE_SEGMENT|1882,1886|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1882,1886|false|false|false|C0582103|Medical Examination|Exam
Finding|Idea or Concept|SIMPLE_SEGMENT|1898,1902|false|false|false|C1511726|Data|Data
Finding|Gene or Genome|SIMPLE_SEGMENT|1933,1937|false|false|false|C1823816|C1orf210 gene|Temp
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1933,1937|false|false|false|C0279848|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Temp
Finding|Finding|SIMPLE_SEGMENT|2038,2046|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Finding|Functional Concept|SIMPLE_SEGMENT|2038,2046|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Finding|Organism Function|SIMPLE_SEGMENT|2038,2046|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2038,2046|false|false|false|C0011209|Obstetric Delivery|delivery
Finding|Classification|SIMPLE_SEGMENT|2053,2056|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|GEN
Finding|Gene or Genome|SIMPLE_SEGMENT|2053,2056|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|GEN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2065,2068|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2065,2068|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2065,2068|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|2065,2068|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2065,2068|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Finding|Finding|SIMPLE_SEGMENT|2065,2068|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2091,2096|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2110,2116|false|false|false|C0036410|Sclera|sclera
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2110,2116|false|false|false|C0036412|Scleral Diseases|sclera
Procedure|Health Care Activity|SIMPLE_SEGMENT|2110,2116|false|false|false|C2228481|examination of sclera|sclera
Finding|Finding|SIMPLE_SEGMENT|2117,2126|false|false|false|C0205180|Anicteric|anicteric
Procedure|Health Care Activity|SIMPLE_SEGMENT|2135,2139|false|false|false|C1315068|Pulmonary ventilator management|PULM
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2144,2155|true|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|SIMPLE_SEGMENT|2144,2155|true|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|SIMPLE_SEGMENT|2144,2155|true|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|SIMPLE_SEGMENT|2144,2155|true|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Sign or Symptom|SIMPLE_SEGMENT|2144,2164|true|false|false|C0476273|Respiratory distress|respiratory distress
Finding|Finding|SIMPLE_SEGMENT|2156,2164|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|SIMPLE_SEGMENT|2156,2164|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2165,2168|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|ABD
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|2165,2168|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|ABD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2170,2174|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Finding|Finding|SIMPLE_SEGMENT|2198,2206|true|false|false|C0427198|Protective muscle spasm|guarding
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|2208,2211|false|false|false|C0015306|Hereditary Multiple Exostoses|EXT
Finding|Gene or Genome|SIMPLE_SEGMENT|2208,2211|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|EXT
Finding|Finding|SIMPLE_SEGMENT|2213,2217|false|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2213,2217|false|false|false|C0687712|warming process|warm
Finding|Finding|SIMPLE_SEGMENT|2219,2223|false|false|false|C5575035|Well (answer to question)|well
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2237,2242|true|false|false|C1717255||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|2237,2242|true|false|false|C0013604|Edema|edema
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2244,2249|false|false|false|C0004936;C1306597|Mental disorders;Psychiatric problem|PSYCH
Finding|Mental Process|SIMPLE_SEGMENT|2258,2265|false|false|false|C0233820|Insight|insight
Finding|Finding|SIMPLE_SEGMENT|2267,2273|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Intellectual Product|SIMPLE_SEGMENT|2267,2273|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Mental Process|SIMPLE_SEGMENT|2267,2273|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2279,2283|false|false|false|C2713234||mood
Finding|Conceptual Entity|SIMPLE_SEGMENT|2279,2283|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|mood
Finding|Finding|SIMPLE_SEGMENT|2279,2283|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|mood
Finding|Mental Process|SIMPLE_SEGMENT|2279,2283|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|mood
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|2284,2289|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|WOUND
Finding|Body Substance|SIMPLE_SEGMENT|2284,2289|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|WOUND
Finding|Functional Concept|SIMPLE_SEGMENT|2284,2289|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|WOUND
Finding|Intellectual Product|SIMPLE_SEGMENT|2284,2289|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|WOUND
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2294,2302|false|false|false|C2338258|Cranial incision point|Incision
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|2294,2302|false|false|false|C0332803|Surgical wound|Incision
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2294,2302|false|false|false|C0184898|Surgical incisions|Incision
Finding|Intellectual Product|SIMPLE_SEGMENT|2311,2316|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|2317,2325|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2317,2332|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|2317,2332|false|false|false|C0489547|Hospital course|Hospital Course
Finding|Idea or Concept|SIMPLE_SEGMENT|2351,2355|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|SIMPLE_SEGMENT|2351,2355|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Finding|SIMPLE_SEGMENT|2360,2364|false|false|false|C1706180|Male Gender|Male
Finding|Finding|SIMPLE_SEGMENT|2424,2432|false|false|false|C0332149|Possible|possibly
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|2438,2445|false|false|false|C0302912|Radicals (chemistry)|radical
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2446,2452|false|false|false|C4522154|Distal Resection Margin|distal
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2454,2465|false|false|false|C0017118|Gastrectomy|gastrectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2471,2486|false|false|false|C0024203|Lymph node excision|lymphadenectomy
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2508,2515|false|false|false|C0038351|Stomach|gastric
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2517,2526|false|false|false|C0007097|Carcinoma|carcinoma
Finding|Functional Concept|SIMPLE_SEGMENT|2533,2545|false|false|false|C0013217|pharmacotherapeutic|chemotherapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2533,2545|false|false|false|C0013216;C0392920;C3665472|Chemotherapy;Chemotherapy Regimen;Pharmacotherapy|chemotherapy
Procedure|Health Care Activity|SIMPLE_SEGMENT|2553,2562|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2553,2562|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Finding|Functional Concept|SIMPLE_SEGMENT|2570,2575|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Drug|Food|SIMPLE_SEGMENT|2592,2596|false|false|false|C0452253|Port - alcoholic beverage|port
Finding|Functional Concept|SIMPLE_SEGMENT|2598,2610|false|false|false|C4281791|Insufflation route|insufflation
Procedure|Health Care Activity|SIMPLE_SEGMENT|2598,2610|false|false|false|C0021634|Insufflation|insufflation
Finding|Functional Concept|SIMPLE_SEGMENT|2624,2629|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2624,2644|false|false|false|C0230177|Structure of right upper quadrant of abdomen|right upper quadrant
Drug|Food|SIMPLE_SEGMENT|2646,2650|false|false|false|C0452253|Port - alcoholic beverage|port
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2673,2680|false|false|false|C0028977|Omentum|omentum
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2707,2727|false|false|false|C0230254|Structure of transverse mesocolon|transverse mesocolon
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2718,2727|false|false|false|C0025483|Mesocolon|mesocolon
Finding|Finding|SIMPLE_SEGMENT|2731,2735|false|false|false|C5575035|Well (answer to question)|well
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2743,2748|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2743,2748|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2743,2748|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Finding|Finding|SIMPLE_SEGMENT|2743,2748|false|false|false|C0750873|COLON PROBLEM|colon
Finding|Finding|SIMPLE_SEGMENT|2769,2776|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|2769,2776|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|2769,2776|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2769,2776|false|false|false|C0543467|Operative Surgical Procedures|surgery
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2806,2816|false|false|false|C0031153;C0442034|Peritoneum;peritoneal|peritoneal
Anatomy|Tissue|SIMPLE_SEGMENT|2806,2816|false|false|false|C0031153;C0442034|Peritoneum;peritoneal|peritoneal
Finding|Functional Concept|SIMPLE_SEGMENT|2817,2825|false|false|false|C0333562|Deposition (morphologic abnormality)|deposits
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2834,2844|false|false|false|C0031153;C0442034|Peritoneum;peritoneal|peritoneal
Anatomy|Tissue|SIMPLE_SEGMENT|2834,2844|false|false|false|C0031153;C0442034|Peritoneum;peritoneal|peritoneal
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2908,2922|false|false|false|C0205699;C2007060|Carcinomatosis;carcinomatosis of unspecified behavior|carcinomatosis
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2947,2961|false|false|false|C0001418;C5551397|Adenocarcinoma;Malignant adenomatous neoplasm|adenocarcinoma
Anatomy|Tissue|SIMPLE_SEGMENT|2977,2987|false|false|false|C0031153;C0230198;C4482223|Abdomen>Peritoneum;Peritoneum;Serous layer of peritoneum|peritoneum
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2977,2987|false|false|false|C0496874;C0496954|Benign neoplasm of peritoneum;Neoplasm of uncertain or unknown behavior of peritoneum|peritoneum
Finding|Idea or Concept|SIMPLE_SEGMENT|2998,3004|false|false|false|C0392360|Indication of (contextual qualifier)|reason
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3010,3019|false|false|false|C0945766||procedure
Event|Occupational Activity|SIMPLE_SEGMENT|3010,3019|false|false|false|C1546467|Act Class - procedure|procedure
Finding|Functional Concept|SIMPLE_SEGMENT|3010,3019|false|false|false|C2700391|Procedure (set of actions)|procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3010,3019|false|false|false|C0184661|Interventional procedure|procedure
Finding|Intellectual Product|SIMPLE_SEGMENT|3025,3029|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Body Substance|SIMPLE_SEGMENT|3060,3067|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|3060,3067|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|3060,3067|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|3097,3103|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Intellectual Product|SIMPLE_SEGMENT|3108,3112|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Intellectual Product|SIMPLE_SEGMENT|3144,3150|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Idea or Concept|SIMPLE_SEGMENT|3158,3162|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|3158,3162|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|3158,3162|false|false|false|C1553498|home health encounter|home
Finding|Body Substance|SIMPLE_SEGMENT|3178,3185|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|3178,3185|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|3178,3185|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3190,3195|false|false|false|C5890168||alert
Drug|Organic Chemical|SIMPLE_SEGMENT|3190,3195|false|false|false|C0718338|Alert brand of caffeine|alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3190,3195|false|false|false|C0718338|Alert brand of caffeine|alert
Finding|Finding|SIMPLE_SEGMENT|3190,3195|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Functional Concept|SIMPLE_SEGMENT|3190,3195|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Intellectual Product|SIMPLE_SEGMENT|3190,3195|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Finding|SIMPLE_SEGMENT|3200,3208|false|false|false|C1961028|Oriented to place|oriented
Procedure|Health Care Activity|SIMPLE_SEGMENT|3221,3236|false|false|false|C0019993|Hospitalization|hospitalization
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3238,3242|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|3238,3242|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|3238,3242|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|3270,3278|false|false|false|C0728755|Dilaudid|dilaudid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3270,3278|false|false|false|C0728755|Dilaudid|dilaudid
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3279,3282|false|false|false|C0149576|Structure of posterior cerebral artery|PCA
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3279,3282|false|false|false|C0268398;C4275079|Familial lichen amyloidosis;Posterior cortical atrophy syndrome|PCA
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3279,3282|false|false|false|C0030131;C0034330|p-Chloroamphetamine;pyrrolidonecarboxylic acid|PCA
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3279,3282|false|false|false|C0030131;C0034330|p-Chloroamphetamine;pyrrolidonecarboxylic acid|PCA
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|3279,3282|false|false|false|C0030131;C0034330|p-Chloroamphetamine;pyrrolidonecarboxylic acid|PCA
Drug|Organic Chemical|SIMPLE_SEGMENT|3279,3282|false|false|false|C0030131;C0034330|p-Chloroamphetamine;pyrrolidonecarboxylic acid|PCA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3279,3282|false|false|false|C0030131;C0034330|p-Chloroamphetamine;pyrrolidonecarboxylic acid|PCA
Finding|Finding|SIMPLE_SEGMENT|3279,3282|false|false|false|C0220723;C1549860;C1836722|CHOANAL ATRESIA, POSTERIOR;FLVCR1 gene;PCA Message Structure|PCA
Finding|Gene or Genome|SIMPLE_SEGMENT|3279,3282|false|false|false|C0220723;C1549860;C1836722|CHOANAL ATRESIA, POSTERIOR;FLVCR1 gene;PCA Message Structure|PCA
Finding|Intellectual Product|SIMPLE_SEGMENT|3279,3282|false|false|false|C0220723;C1549860;C1836722|CHOANAL ATRESIA, POSTERIOR;FLVCR1 gene;PCA Message Structure|PCA
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3279,3282|false|false|false|C0030625;C0078944;C5968782|Passive Cutaneous Anaphylaxis;Patient controlled intravenous analgesia;Patient-Controlled Analgesia|PCA
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3279,3282|false|false|false|C0030625;C0078944;C5968782|Passive Cutaneous Anaphylaxis;Patient controlled intravenous analgesia;Patient-Controlled Analgesia|PCA
Finding|Intellectual Product|SIMPLE_SEGMENT|3311,3315|false|false|false|C1720594|Then - dosing instruction fragment|then
Drug|Organic Chemical|SIMPLE_SEGMENT|3332,3340|false|false|false|C0040610|tramadol|tramadol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3332,3340|false|false|false|C0040610|tramadol|tramadol
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3332,3340|false|false|false|C1266765|Tramadol measurement (procedure)|tramadol
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3370,3374|false|false|false|C2598155||Pain
Finding|Functional Concept|SIMPLE_SEGMENT|3370,3374|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|3370,3374|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Finding|SIMPLE_SEGMENT|3379,3388|false|false|false|C5202951;C5202952;C5202953|Can Do Very Well;Describes Very Well;Very Well|very well
Finding|Finding|SIMPLE_SEGMENT|3384,3388|false|false|false|C5575035|Well (answer to question)|well
Finding|Body Substance|SIMPLE_SEGMENT|3411,3418|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|3411,3418|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|3411,3418|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|3428,3434|false|false|false|C1547311|Patient Condition Code - Stable|stable
Anatomy|Body System|SIMPLE_SEGMENT|3442,3456|false|false|false|C0007226;C3887460|Cardiovascular;Cardiovascular system|cardiovascular
Drug|Food|SIMPLE_SEGMENT|3470,3475|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|vital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3470,3481|false|false|false|C0488614;C0518766|Vital signs|vital signs
Procedure|Health Care Activity|SIMPLE_SEGMENT|3470,3481|false|false|false|C0150404|Taking vital signs|vital signs
Finding|Finding|SIMPLE_SEGMENT|3476,3481|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|3476,3481|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3512,3521|false|false|false|C0024109|Lung|PULMONARY
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3512,3521|false|false|false|C2707265||PULMONARY
Finding|Finding|SIMPLE_SEGMENT|3512,3521|false|false|false|C4522268|Pulmonary (intended site)|PULMONARY
Finding|Body Substance|SIMPLE_SEGMENT|3527,3534|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|3527,3534|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|3527,3534|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|3544,3550|false|false|false|C1547311|Patient Condition Code - Stable|stable
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3558,3567|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3558,3567|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|3558,3567|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Drug|Food|SIMPLE_SEGMENT|3581,3586|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|vital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3581,3592|false|false|false|C0488614;C0518766|Vital signs|vital signs
Procedure|Health Care Activity|SIMPLE_SEGMENT|3581,3592|false|false|false|C0150404|Taking vital signs|vital signs
Finding|Finding|SIMPLE_SEGMENT|3587,3592|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|3587,3592|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Idea or Concept|SIMPLE_SEGMENT|3619,3623|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|Good
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3624,3633|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3624,3633|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|3624,3633|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3635,3641|false|false|false|C0184958|Toilet procedure|toilet
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3643,3659|false|false|false|C0013457|Early Ambulation|early ambulation
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|3649,3659|false|false|false|C0080331;C0945826|Ambulation;Walking (function)|ambulation
Finding|Functional Concept|SIMPLE_SEGMENT|3649,3659|false|false|false|C0080331;C0945826|Ambulation;Walking (function)|ambulation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3664,3684|false|false|false|C0454512|Incentive spirometry|incentive spirometry
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3674,3684|false|false|false|C0037981|Spirometry|spirometry
Procedure|Health Care Activity|SIMPLE_SEGMENT|3713,3728|false|false|false|C0019993|Hospitalization|hospitalization
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3756,3765|false|false|false|C0945766||procedure
Event|Occupational Activity|SIMPLE_SEGMENT|3756,3765|false|false|false|C1546467|Act Class - procedure|procedure
Finding|Functional Concept|SIMPLE_SEGMENT|3756,3765|false|false|false|C2700391|Procedure (set of actions)|procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3756,3765|false|false|false|C0184661|Interventional procedure|procedure
Finding|Finding|SIMPLE_SEGMENT|3788,3794|false|false|false|C1299582|Unable|unable
Finding|Finding|SIMPLE_SEGMENT|3799,3803|false|false|false|C2828386|Pass (indicator)|pass
Event|Event|SIMPLE_SEGMENT|3816,3823|false|false|false|C1516084|Attempt|attempt
Finding|Idea or Concept|SIMPLE_SEGMENT|3829,3837|false|false|false|C1548173;C2828392|Standard (document);Type of Agreement - Standard|standard
Finding|Intellectual Product|SIMPLE_SEGMENT|3829,3837|false|false|false|C1548173;C2828392|Standard (document);Type of Agreement - Standard|standard
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3829,3837|false|false|false|C3873211|Standard base excess calculation technique|standard
Finding|Gene or Genome|SIMPLE_SEGMENT|3848,3852|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Intellectual Product|SIMPLE_SEGMENT|3848,3852|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Finding|SIMPLE_SEGMENT|3874,3881|false|false|false|C0021359;C4074771|Infertility;Sterility, Reproductive|sterile
Finding|Pathologic Function|SIMPLE_SEGMENT|3874,3881|false|false|false|C0021359;C4074771|Infertility;Sterility, Reproductive|sterile
Finding|Functional Concept|SIMPLE_SEGMENT|3882,3891|false|false|false|C0449851|Techniques|technique
Procedure|Health Care Activity|SIMPLE_SEGMENT|3913,3922|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3913,3922|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Finding|Functional Concept|SIMPLE_SEGMENT|3941,3952|false|false|false|C0870325;C1547755;C1947919;C2347934;C4048755|Application Document;Apply;Computer Application;HL7 Version 2.5 - Application;Regulatory Application|application
Finding|Idea or Concept|SIMPLE_SEGMENT|3941,3952|false|false|false|C0870325;C1547755;C1947919;C2347934;C4048755|Application Document;Apply;Computer Application;HL7 Version 2.5 - Application;Regulatory Application|application
Finding|Intellectual Product|SIMPLE_SEGMENT|3941,3952|false|false|false|C0870325;C1547755;C1947919;C2347934;C4048755|Application Document;Apply;Computer Application;HL7 Version 2.5 - Application;Regulatory Application|application
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3941,3952|false|false|false|C0185125|Application procedure|application
Finding|Gene or Genome|SIMPLE_SEGMENT|3977,3981|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Intellectual Product|SIMPLE_SEGMENT|3977,3981|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Finding|SIMPLE_SEGMENT|4005,4011|false|false|false|C1299582|Unable|unable
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4031,4039|false|false|false|C0033572;C4266527|Prostate;Structure of prostate (body structure)|prostate
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4031,4039|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|prostate
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4031,4039|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|prostate
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4128,4135|false|false|false|C0041967|Urethra|urethra
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4128,4135|false|false|false|C0041969;C0153620;C0154019;C0496929|Benign neoplasm of urethra;Malignant neoplasm of urethra;Neoplasm of uncertain or unknown behavior of urethra;Urethral Diseases|urethra
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4128,4135|false|false|false|C0041969;C0153620;C0154019;C0496929|Benign neoplasm of urethra;Malignant neoplasm of urethra;Neoplasm of uncertain or unknown behavior of urethra;Urethral Diseases|urethra
Finding|Body Substance|SIMPLE_SEGMENT|4128,4135|false|false|false|C1547951;C1550675|Urethra specimen;Urethra specimen code|urethra
Finding|Intellectual Product|SIMPLE_SEGMENT|4128,4135|false|false|false|C1547951;C1550675|Urethra specimen;Urethra specimen code|urethra
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4128,4135|false|false|false|C0810170|Procedure on urethra|urethra
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4199,4206|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4199,4206|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4199,4206|false|false|false|C0872388|Procedures on bladder|bladder
Finding|Conceptual Entity|SIMPLE_SEGMENT|4212,4217|false|false|false|C1710028|Scope|scope
Finding|Gene or Genome|SIMPLE_SEGMENT|4273,4277|false|false|false|C1823858|WIPF2 gene|wire
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4291,4299|false|false|false|C0033572;C4266527|Prostate;Structure of prostate (body structure)|prostate
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4291,4299|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|prostate
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4291,4299|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|prostate
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4313,4320|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4313,4320|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4313,4320|false|false|false|C0872388|Procedures on bladder|bladder
Finding|Body Substance|SIMPLE_SEGMENT|4326,4333|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|4326,4333|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|4326,4333|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Activity|SIMPLE_SEGMENT|4368,4373|false|false|false|C1882509|put - instruction imperative|place
Finding|Functional Concept|SIMPLE_SEGMENT|4368,4373|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|SIMPLE_SEGMENT|4368,4373|false|false|false|C1533810||place
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4379,4391|false|false|false|C3263700||instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|4379,4391|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|instructions
Finding|Classification|SIMPLE_SEGMENT|4422,4432|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|4422,4432|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Functional Concept|SIMPLE_SEGMENT|4455,4462|false|false|false|C0042034;C4067975|Urination;Voids|voiding
Finding|Organism Function|SIMPLE_SEGMENT|4455,4462|false|false|false|C0042034;C4067975|Urination;Voids|voiding
Procedure|Research Activity|SIMPLE_SEGMENT|4463,4468|false|false|false|C0008976|Clinical Trials|trial
Drug|Antibiotic|SIMPLE_SEGMENT|4473,4484|true|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Finding|Body Substance|SIMPLE_SEGMENT|4508,4515|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|4508,4515|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|4508,4515|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|4534,4546|false|false|false|C0184625||regular diet
Drug|Food|SIMPLE_SEGMENT|4542,4546|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Finding|Functional Concept|SIMPLE_SEGMENT|4542,4546|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|SIMPLE_SEGMENT|4542,4546|false|false|false|C0012159|Diet therapy|diet
Finding|Body Substance|SIMPLE_SEGMENT|4556,4565|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|4556,4565|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|4556,4565|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|4556,4565|false|false|false|C0030685|Patient Discharge|discharge
Finding|Body Substance|SIMPLE_SEGMENT|4578,4585|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|4578,4585|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|4578,4585|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|SIMPLE_SEGMENT|4588,4593|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|4588,4593|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Finding|SIMPLE_SEGMENT|4626,4631|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|4626,4631|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4636,4645|false|false|false|C0009450|Communicable Diseases|infection
Finding|Pathologic Function|SIMPLE_SEGMENT|4636,4645|false|false|false|C3714514|Infection|infection
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4677,4681|false|false|false|C0018966|Heme|HEME
Drug|Organic Chemical|SIMPLE_SEGMENT|4677,4681|false|false|false|C0018966|Heme|HEME
Finding|Body Substance|SIMPLE_SEGMENT|4683,4690|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|4683,4690|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|4683,4690|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|4700,4703|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4700,4703|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4700,4703|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|4700,4703|false|false|false|C1332410|BID gene|BID
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4712,4715|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4712,4715|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4712,4715|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4712,4727|false|false|false|C0853245|DVT prophylaxis|DVT prophylaxis
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4716,4727|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Finding|Functional Concept|SIMPLE_SEGMENT|4732,4740|false|false|false|C0332287;C1883712|Add - instruction imperative;In addition to|addition
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4757,4773|false|false|false|C0013457|Early Ambulation|early ambulation
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|4763,4773|false|false|false|C0080331;C0945826|Ambulation;Walking (function)|ambulation
Finding|Functional Concept|SIMPLE_SEGMENT|4763,4773|false|false|false|C0080331;C0945826|Ambulation;Walking (function)|ambulation
Finding|Functional Concept|SIMPLE_SEGMENT|4787,4798|false|false|false|C0332459;C4551657|Compressed structure|compression
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|4787,4798|false|false|false|C0728907|Compression|compression
Procedure|Machine Activity|SIMPLE_SEGMENT|4787,4798|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4787,4798|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Finding|Gene or Genome|SIMPLE_SEGMENT|4812,4816|false|false|false|C1420638;C1539127;C1710283|CORO7 gene;TCF21 gene;TCF21 wt Allele|POD1
Finding|Body Substance|SIMPLE_SEGMENT|4821,4828|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|4821,4828|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|4821,4828|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|4850,4854|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|4850,4854|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|4850,4854|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|4856,4866|false|false|false|C0206460|enoxaparin|enoxaparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4856,4866|false|false|false|C0206460|enoxaparin|enoxaparin
Finding|Body Substance|SIMPLE_SEGMENT|4874,4883|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|4874,4883|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|4874,4883|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|4874,4883|false|false|false|C0030685|Patient Discharge|discharge
Finding|Idea or Concept|SIMPLE_SEGMENT|4887,4899|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Finding|Finding|SIMPLE_SEGMENT|4936,4940|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|4936,4940|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|4936,4940|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Body Substance|SIMPLE_SEGMENT|4944,4953|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|4944,4953|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|4944,4953|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|4944,4953|false|false|false|C0030685|Patient Discharge|discharge
Finding|Body Substance|SIMPLE_SEGMENT|4959,4966|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|4959,4966|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|4959,4966|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|SIMPLE_SEGMENT|4977,4981|false|false|false|C5575035|Well (answer to question)|well
Finding|Finding|SIMPLE_SEGMENT|4983,4991|false|false|false|C0277797|Apyrexial|afebrile
Finding|Intellectual Product|SIMPLE_SEGMENT|4998,5004|false|false|false|C1547311|Patient Condition Code - Stable|stable
Drug|Food|SIMPLE_SEGMENT|5005,5010|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|vital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5005,5016|false|false|false|C0488614;C0518766|Vital signs|vital signs
Procedure|Health Care Activity|SIMPLE_SEGMENT|5005,5016|false|false|false|C0150404|Taking vital signs|vital signs
Finding|Finding|SIMPLE_SEGMENT|5011,5016|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|5011,5016|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Body Substance|SIMPLE_SEGMENT|5022,5029|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|5022,5029|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|5022,5029|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Food|SIMPLE_SEGMENT|5045,5049|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Finding|Functional Concept|SIMPLE_SEGMENT|5045,5049|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|SIMPLE_SEGMENT|5045,5049|false|false|false|C0012159|Diet therapy|diet
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5064,5068|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5064,5068|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|5064,5068|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|5064,5068|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5086,5090|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|5086,5090|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|5086,5090|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|SIMPLE_SEGMENT|5095,5099|false|false|false|C5575035|Well (answer to question)|well
Finding|Body Substance|SIMPLE_SEGMENT|5117,5124|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|5117,5124|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|5117,5124|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|5140,5144|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|5140,5144|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|5140,5144|false|false|false|C1553498|home health encounter|home
Finding|Intellectual Product|SIMPLE_SEGMENT|5160,5168|false|false|false|C1546572||catheter
Finding|Intellectual Product|SIMPLE_SEGMENT|5187,5195|false|false|false|C1548344|Visit User Code - Teaching|teaching
Procedure|Educational Activity|SIMPLE_SEGMENT|5187,5195|false|false|false|C0039401;C0220924|Education (procedure);Teaching aspects|teaching
Event|Activity|SIMPLE_SEGMENT|5200,5204|false|false|false|C1947933|care activity|care
Finding|Finding|SIMPLE_SEGMENT|5200,5204|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|5200,5204|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Body Substance|SIMPLE_SEGMENT|5210,5217|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|5210,5217|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|5210,5217|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Body Substance|SIMPLE_SEGMENT|5227,5236|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|5227,5236|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|5227,5236|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|5227,5236|false|false|false|C0030685|Patient Discharge|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|5238,5246|false|false|false|C1548344|Visit User Code - Teaching|teaching
Procedure|Educational Activity|SIMPLE_SEGMENT|5238,5246|false|false|false|C0039401;C0220924|Education (procedure);Teaching aspects|teaching
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5261,5273|false|false|false|C3263700||instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|5261,5273|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|instructions
Finding|Mental Process|SIMPLE_SEGMENT|5279,5292|false|false|false|C0162340|Comprehension|understanding
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5309,5318|false|false|false|C4255433||agreement
Finding|Intellectual Product|SIMPLE_SEGMENT|5309,5318|false|false|false|C0680240;C4255373|Agreement;Agreement (document)|agreement
Finding|Social Behavior|SIMPLE_SEGMENT|5309,5318|false|false|false|C0680240;C4255373|Agreement;Agreement (document)|agreement
Finding|Body Substance|SIMPLE_SEGMENT|5328,5337|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|5328,5337|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|5328,5337|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|5328,5337|false|false|false|C0030685|Patient Discharge|discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5328,5342|false|false|false|C2745873||discharge plan
Finding|Intellectual Product|SIMPLE_SEGMENT|5328,5342|false|false|false|C2735970|Discharge plan|discharge plan
Procedure|Health Care Activity|SIMPLE_SEGMENT|5328,5342|false|false|false|C0012622|Discharge Planning|discharge plan
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5338,5342|false|false|false|C0270724|Infantile Neuroaxonal Dystrophy|plan
Finding|Functional Concept|SIMPLE_SEGMENT|5338,5342|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Intellectual Product|SIMPLE_SEGMENT|5338,5342|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Mental Process|SIMPLE_SEGMENT|5338,5342|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5346,5357|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5346,5357|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|5346,5357|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|5346,5370|false|false|false|C1627937|Medications on admission|Medications on Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|5361,5370|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5372,5383|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5372,5383|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|5372,5383|false|false|false|C4284232|Medications|Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5386,5398|false|false|false|C5886759|Prescription (attribute)|Prescription
Finding|Intellectual Product|SIMPLE_SEGMENT|5386,5398|false|false|false|C1521941|prescription document|Prescription
Procedure|Health Care Activity|SIMPLE_SEGMENT|5386,5398|false|false|false|C0033080|Prescription (procedure)|Prescription
Drug|Hormone|SIMPLE_SEGMENT|5399,5409|false|false|false|C1878933|Bio-Throid|BIO-THROID
Drug|Organic Chemical|SIMPLE_SEGMENT|5399,5409|false|false|false|C1878933|Bio-Throid|BIO-THROID
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5399,5409|false|false|false|C1878933|Bio-Throid|BIO-THROID
Drug|Hormone|SIMPLE_SEGMENT|5412,5422|false|false|false|C1878933|Bio-Throid|Bio-Throid
Drug|Organic Chemical|SIMPLE_SEGMENT|5412,5422|false|false|false|C1878933|Bio-Throid|Bio-Throid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5412,5422|false|false|false|C1878933|Bio-Throid|Bio-Throid
Finding|Intellectual Product|SIMPLE_SEGMENT|5433,5437|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5433,5443|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|SIMPLE_SEGMENT|5440,5443|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|5440,5443|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Functional Concept|SIMPLE_SEGMENT|5469,5477|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|Provider
Finding|Intellectual Product|SIMPLE_SEGMENT|5469,5477|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|Provider
Drug|Organic Chemical|SIMPLE_SEGMENT|5479,5489|false|false|false|C0206460|enoxaparin|ENOXAPARIN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5479,5489|false|false|false|C0206460|enoxaparin|ENOXAPARIN
Drug|Organic Chemical|SIMPLE_SEGMENT|5492,5502|false|false|false|C0206460|enoxaparin|enoxaparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5492,5502|false|false|false|C0206460|enoxaparin|enoxaparin
Finding|Functional Concept|SIMPLE_SEGMENT|5517,5529|false|false|false|C1522438|Subcutaneous Route of Administration|subcutaneous
Drug|Organic Chemical|SIMPLE_SEGMENT|5556,5566|false|false|false|C0028978|omeprazole|OMEPRAZOLE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5556,5566|false|false|false|C0028978|omeprazole|OMEPRAZOLE
Drug|Organic Chemical|SIMPLE_SEGMENT|5569,5579|false|false|false|C0028978|omeprazole|omeprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5569,5579|false|false|false|C0028978|omeprazole|omeprazole
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5586,5593|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|5586,5593|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5586,5593|false|false|false|C0006935|capsule (pharmacologic)|capsule
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5614,5621|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|5614,5621|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5614,5621|false|false|false|C0006935|capsule (pharmacologic)|capsule
Finding|Functional Concept|SIMPLE_SEGMENT|5625,5633|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5628,5633|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5628,5633|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Organic Chemical|SIMPLE_SEGMENT|5646,5655|false|false|false|C0077656|ubiquinol|UBIQUINOL
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5646,5655|false|false|false|C0077656|ubiquinol|UBIQUINOL
Drug|Organic Chemical|SIMPLE_SEGMENT|5658,5667|false|false|false|C0077656|ubiquinol|ubiquinol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5658,5667|false|false|false|C0077656|ubiquinol|ubiquinol
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5687,5692|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5687,5692|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|SIMPLE_SEGMENT|5701,5704|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|5701,5704|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Functional Concept|SIMPLE_SEGMENT|5730,5738|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|Provider
Finding|Intellectual Product|SIMPLE_SEGMENT|5730,5738|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|Provider
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5742,5753|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5742,5753|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|5742,5753|false|false|false|C4284232|Medications|Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5756,5759|false|false|false|C0013231|Drugs, Non-Prescription|OTC
Finding|Gene or Genome|SIMPLE_SEGMENT|5756,5759|false|false|false|C1418193|OTC gene|OTC
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|5760,5767|false|false|false|C2346592|Ferrous|FERROUS
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5760,5775|false|false|false|C0060282|ferrous sulfate|FERROUS SULFATE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5760,5775|false|false|false|C0060282|ferrous sulfate|FERROUS SULFATE
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|5768,5775|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|SULFATE
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5768,5775|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|SULFATE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5768,5775|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|SULFATE
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|5778,5785|false|false|false|C2346592|Ferrous|ferrous
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5778,5793|false|false|false|C0060282|ferrous sulfate|ferrous sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5778,5793|false|false|false|C0060282|ferrous sulfate|ferrous sulfate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|5786,5793|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5786,5793|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5786,5793|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5808,5812|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|5808,5812|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5808,5812|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5808,5812|false|false|false|C0337439|Iron measurement|iron
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5825,5831|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|SIMPLE_SEGMENT|5835,5843|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5838,5843|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5838,5843|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|SIMPLE_SEGMENT|5852,5855|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|5852,5855|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Functional Concept|SIMPLE_SEGMENT|5880,5888|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|Provider
Finding|Intellectual Product|SIMPLE_SEGMENT|5880,5888|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|Provider
Finding|Finding|SIMPLE_SEGMENT|5904,5915|false|false|false|C3811910|combination - answer to question|COMBINATION
Finding|Finding|SIMPLE_SEGMENT|5942,5951|false|false|false|C0087130|Uncertainty|uncertain
Finding|Functional Concept|SIMPLE_SEGMENT|5977,5985|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|Provider
Finding|Intellectual Product|SIMPLE_SEGMENT|5977,5985|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|Provider
Finding|Body Substance|SIMPLE_SEGMENT|5996,6005|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|5996,6005|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|5996,6005|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|5996,6005|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|5996,6017|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6006,6017|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6006,6017|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|6006,6017|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|6023,6036|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6023,6036|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6023,6036|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Organic Chemical|SIMPLE_SEGMENT|6058,6066|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6058,6066|false|false|false|C1692318|docusate|Docusate
Drug|Organic Chemical|SIMPLE_SEGMENT|6058,6073|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6058,6073|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6067,6073|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|6067,6073|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6067,6073|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|6067,6073|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6067,6073|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|6084,6087|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6084,6087|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6084,6087|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|6084,6087|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|6094,6099|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6094,6099|false|false|false|C3489575|sennosides, USP|Senna
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|6110,6113|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6110,6113|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6110,6113|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|6110,6113|false|false|false|C1332410|BID gene|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|6114,6117|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Sign or Symptom|SIMPLE_SEGMENT|6118,6130|false|false|false|C0009806|Constipation|Constipation
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6139,6143|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|6139,6143|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Drug|Substance|SIMPLE_SEGMENT|6139,6143|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Finding|Intellectual Product|SIMPLE_SEGMENT|6139,6143|false|false|false|C1546701|line source specimen code|Line
Drug|Organic Chemical|SIMPLE_SEGMENT|6150,6158|false|false|false|C0040610|tramadol|TraMADol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6150,6158|false|false|false|C0040610|tramadol|TraMADol
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6150,6158|false|false|false|C1266765|Tramadol measurement (procedure)|TraMADol
Finding|Gene or Genome|SIMPLE_SEGMENT|6172,6175|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6176,6180|false|false|false|C2598155||Pain
Finding|Functional Concept|SIMPLE_SEGMENT|6176,6180|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6176,6180|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Finding|SIMPLE_SEGMENT|6183,6191|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|6183,6191|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6198,6208|false|false|false|C0013227|Pharmaceutical Preparations|medication
Finding|Intellectual Product|SIMPLE_SEGMENT|6198,6208|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Finding|Finding|SIMPLE_SEGMENT|6214,6217|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|SIMPLE_SEGMENT|6214,6217|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|6223,6231|false|false|false|C0027415|Narcotics|narcotic
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6223,6231|false|false|false|C0027415|Narcotics|narcotic
Finding|Conceptual Entity|SIMPLE_SEGMENT|6240,6245|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Finding|Functional Concept|SIMPLE_SEGMENT|6240,6245|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Finding|Sign or Symptom|SIMPLE_SEGMENT|6247,6259|false|false|false|C0009806|Constipation|constipation
Drug|Organic Chemical|SIMPLE_SEGMENT|6266,6274|false|false|false|C0040610|tramadol|tramadol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6266,6274|false|false|false|C0040610|tramadol|tramadol
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6266,6274|false|false|false|C1266765|Tramadol measurement (procedure)|tramadol
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6289,6295|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|SIMPLE_SEGMENT|6299,6307|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6302,6307|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6302,6307|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6339,6345|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|SIMPLE_SEGMENT|6346,6353|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|6362,6372|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6362,6372|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Organic Chemical|SIMPLE_SEGMENT|6362,6379|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6362,6379|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6373,6379|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|6373,6379|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6373,6379|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|6373,6379|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6373,6379|false|false|false|C0337443|Sodium measurement|Sodium
Finding|Body Substance|SIMPLE_SEGMENT|6401,6410|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6401,6410|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6401,6410|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6401,6410|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6401,6422|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|6401,6422|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6411,6422|false|false|false|C2926604||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|6411,6422|false|false|false|C0184758|Patient disposition|Disposition
Finding|Idea or Concept|SIMPLE_SEGMENT|6424,6428|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|6424,6428|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|6424,6428|false|false|false|C1553498|home health encounter|Home
Finding|Body Substance|SIMPLE_SEGMENT|6431,6440|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6431,6440|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6431,6440|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6431,6440|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|6431,6450|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6441,6450|false|false|false|C0945731||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|6441,6450|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|6441,6450|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6441,6450|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|6452,6462|false|false|false|C0036525;C1522484|Metastatic to;metastatic qualifier|Metastatic
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6452,6477|false|false|false|C0278498|Malignant neoplasm of stomach stage IV|Metastatic gastric cancer
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6463,6470|false|false|false|C0038351|Stomach|gastric
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6463,6477|false|false|false|C0024623;C0699791|Malignant neoplasm of stomach;Stomach Carcinoma|gastric cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6471,6477|false|false|false|C0006826|Malignant Neoplasms|cancer
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6479,6484|false|false|false|C1300072|Tumor stage|stage
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6498,6506|false|false|false|C0041967|Urethra|Urethral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6498,6506|false|false|false|C2349082|Urethral Dosage Form|Urethral
Finding|Functional Concept|SIMPLE_SEGMENT|6498,6506|false|false|false|C1522518|Intraurethral Route of Administration|Urethral
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6498,6516|false|false|false|C0041974|Urethral Stenosis|Urethral stricture
Finding|Pathologic Function|SIMPLE_SEGMENT|6498,6516|false|false|false|C4551691|Urethral stricture|Urethral stricture
Finding|Pathologic Function|SIMPLE_SEGMENT|6507,6516|false|false|false|C1261287|Stenosis|stricture
Finding|Body Substance|SIMPLE_SEGMENT|6519,6528|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6519,6528|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6519,6528|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6519,6528|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6529,6538|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6529,6538|false|false|false|C0012634|Disease|Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|6529,6538|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|6540,6546|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6540,6553|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|6540,6553|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6547,6553|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|6547,6553|false|false|false|C1546481|What subject filter - Status|Status
Finding|Idea or Concept|SIMPLE_SEGMENT|6555,6560|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Finding|SIMPLE_SEGMENT|6565,6573|false|false|false|C4068804|Coherent|coherent
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6575,6597|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|6575,6597|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|6584,6597|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|6584,6597|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6599,6604|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|6599,6604|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6599,6604|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|SIMPLE_SEGMENT|6599,6604|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|6599,6604|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|6599,6604|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|6609,6620|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|6622,6630|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|6622,6630|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|6622,6630|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6631,6637|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|6631,6637|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|SIMPLE_SEGMENT|6639,6649|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|6639,6649|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|6639,6649|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|6639,6649|false|false|false|C1561560|ambulatory encounter|Ambulatory
Finding|Finding|SIMPLE_SEGMENT|6652,6663|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|SIMPLE_SEGMENT|6652,6663|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Body Substance|SIMPLE_SEGMENT|6668,6677|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6668,6677|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6668,6677|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6668,6677|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6668,6690|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|6668,6690|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|6668,6690|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6678,6690|false|false|false|C3263700||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|6678,6690|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Finding|Gene or Genome|SIMPLE_SEGMENT|6692,6696|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Finding|Intellectual Product|SIMPLE_SEGMENT|6716,6724|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|SIMPLE_SEGMENT|6716,6724|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|SIMPLE_SEGMENT|6732,6736|false|false|false|C1947933|care activity|care
Finding|Finding|SIMPLE_SEGMENT|6732,6736|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|6732,6736|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|6732,6739|false|false|false|C1555558|care of - AddressPartType|care of
Finding|Idea or Concept|SIMPLE_SEGMENT|6787,6795|false|false|false|C1547192|Organization unit type - Hospital|hospital
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6801,6808|false|false|false|C0038351|Stomach|gastric
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6801,6815|false|false|false|C0024623;C0699791|Malignant neoplasm of stomach;Stomach Carcinoma|gastric cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6809,6815|false|false|false|C0006826|Malignant Neoplasms|cancer
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6853,6865|false|false|false|C0031150|Laparoscopy|laparoscopic
Finding|Idea or Concept|SIMPLE_SEGMENT|6867,6874|false|false|false|C1550516|Target Awareness - partial|partial
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6867,6886|false|false|false|C0030600|Subtotal gastrectomy|partial gastrectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6875,6886|false|false|false|C0017118|Gastrectomy|gastrectomy
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6891,6902|false|false|false|C0017195|Endoscopy of stomach|gastroscopy
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6919,6932|true|false|false|C0802632||complications
Finding|Functional Concept|SIMPLE_SEGMENT|6919,6932|true|false|false|C0009566;C1171258|Complication;complication aspects|complications
Finding|Pathologic Function|SIMPLE_SEGMENT|6919,6932|true|false|false|C0009566;C1171258|Complication;complication aspects|complications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6952,6961|false|false|false|C0945766||procedure
Event|Occupational Activity|SIMPLE_SEGMENT|6952,6961|false|false|false|C1546467|Act Class - procedure|procedure
Finding|Functional Concept|SIMPLE_SEGMENT|6952,6961|false|false|false|C2700391|Procedure (set of actions)|procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6952,6961|false|false|false|C0184661|Interventional procedure|procedure
Finding|Finding|SIMPLE_SEGMENT|6962,6966|false|false|false|C5575035|Well (answer to question)|well
Finding|Body Substance|SIMPLE_SEGMENT|6988,6996|false|false|false|C0015733|Feces|stooling
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|7011,7023|false|false|false|C0184625||regular diet
Drug|Food|SIMPLE_SEGMENT|7019,7023|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Finding|Functional Concept|SIMPLE_SEGMENT|7019,7023|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|SIMPLE_SEGMENT|7019,7023|false|false|false|C0012159|Diet therapy|diet
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7034,7038|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|7034,7038|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|7034,7038|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7057,7061|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|7057,7061|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|7057,7061|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7062,7073|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7062,7073|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|SIMPLE_SEGMENT|7062,7073|false|false|false|C4284232|Medications|medications
Finding|Functional Concept|SIMPLE_SEGMENT|7074,7082|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7077,7082|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|7077,7082|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|SIMPLE_SEGMENT|7123,7127|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|7123,7127|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|7123,7127|false|false|false|C1553498|home health encounter|home
Finding|Idea or Concept|SIMPLE_SEGMENT|7147,7162|false|false|false|C0034866|Recommendation|recommendations
Finding|Finding|SIMPLE_SEGMENT|7193,7203|false|false|false|C5453124|Uneventful|uneventful
Event|Activity|SIMPLE_SEGMENT|7204,7212|false|false|false|C0237820||recovery
Finding|Organism Function|SIMPLE_SEGMENT|7204,7212|false|false|false|C2004454|Recovery - healing process|recovery
Event|Activity|SIMPLE_SEGMENT|7216,7224|false|false|false|C0441655|Activities|ACTIVITY
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|7216,7224|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|ACTIVITY
Finding|Finding|SIMPLE_SEGMENT|7216,7224|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|ACTIVITY
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7271,7275|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|7271,7275|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|7271,7275|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|7271,7284|false|false|false|C0002771|Analgesics|pain medicine
Drug|Organic Chemical|SIMPLE_SEGMENT|7271,7284|false|false|false|C0002771|Analgesics|pain medicine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7271,7284|false|false|false|C0002771|Analgesics|pain medicine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7276,7284|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Finding|Finding|SIMPLE_SEGMENT|7319,7328|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Idea or Concept|SIMPLE_SEGMENT|7319,7328|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Intellectual Product|SIMPLE_SEGMENT|7319,7328|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Pathologic Function|SIMPLE_SEGMENT|7319,7328|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|7319,7328|false|false|false|C0013956|Emergency Situation|emergency
Procedure|Health Care Activity|SIMPLE_SEGMENT|7319,7328|false|false|false|C1553500|emergency encounter|emergency
Finding|Finding|SIMPLE_SEGMENT|7346,7352|false|false|false|C4300351|Prior functioning.stairs|stairs
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7391,7396|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|SIMPLE_SEGMENT|7399,7402|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|7399,7402|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7482,7489|false|false|false|C5444295||surgeon
Finding|Idea or Concept|SIMPLE_SEGMENT|7498,7502|false|false|false|C1552851|next - HtmlLinkType|next
Finding|Social Behavior|SIMPLE_SEGMENT|7503,7508|false|false|false|C0545082|Visit|visit
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7532,7537|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7532,7537|false|false|false|C1570446|TNFSF14 protein, human|light
Finding|Finding|SIMPLE_SEGMENT|7532,7537|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|SIMPLE_SEGMENT|7532,7537|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|SIMPLE_SEGMENT|7532,7537|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|7532,7537|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7532,7537|false|false|false|C0031765|Phototherapy|light
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|7532,7546|false|false|false|C1517883|Light Exercise|light exercise
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|7538,7546|false|false|false|C0015259|Exercise|exercise
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7538,7546|false|false|false|C1522704|Exercise Pain Management|exercise
Finding|Finding|SIMPLE_SEGMENT|7561,7572|false|false|false|C5546696|Feeling comfortable|comfortable
Event|Activity|SIMPLE_SEGMENT|7596,7604|false|false|false|C0441655|Activities|activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|7596,7604|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Finding|Finding|SIMPLE_SEGMENT|7596,7604|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7618,7626|false|false|false|C0168634|BaseLine dental cement|baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|7618,7626|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|7650,7658|false|false|false|C0015259|Exercise|exercise
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7650,7658|false|false|false|C1522704|Exercise Pain Management|exercise
Finding|Functional Concept|SIMPLE_SEGMENT|7697,7703|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Finding|Intellectual Product|SIMPLE_SEGMENT|7697,7703|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|7705,7710|false|false|false|C0036658|Sensory perception|sense
Event|Activity|SIMPLE_SEGMENT|7747,7754|true|false|false|C0206244|Lifting|lifting
Finding|Finding|SIMPLE_SEGMENT|7756,7765|true|false|false|C3845310|10 pounds|10 pounds
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7798,7805|false|false|false|C5444295||surgeon
Finding|Finding|SIMPLE_SEGMENT|7807,7814|false|false|false|C3888388|Usually|usually
Finding|Behavior|SIMPLE_SEGMENT|7848,7854|false|false|false|C0036864|Sex Behavior|sexual
Finding|Behavior|SIMPLE_SEGMENT|7848,7863|false|false|false|C0036864;C5575036|Sex Behavior;Sexual Activity|sexual activity
Finding|Individual Behavior|SIMPLE_SEGMENT|7848,7863|false|false|false|C0036864;C5575036|Sex Behavior;Sexual Activity|sexual activity
Event|Activity|SIMPLE_SEGMENT|7855,7863|false|false|false|C0441655|Activities|activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|7855,7863|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Finding|Finding|SIMPLE_SEGMENT|7855,7863|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Finding|Intellectual Product|SIMPLE_SEGMENT|7876,7882|false|false|false|C2348314|Doctor - Title|doctor
Finding|Mental Process|SIMPLE_SEGMENT|7921,7925|false|false|false|C1527305|Feelings|FEEL
Finding|Intellectual Product|SIMPLE_SEGMENT|7938,7947|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|feel weak
Finding|Sign or Symptom|SIMPLE_SEGMENT|7938,7947|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|feel weak
Finding|Intellectual Product|SIMPLE_SEGMENT|7943,7947|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|weak
Finding|Sign or Symptom|SIMPLE_SEGMENT|7943,7947|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|weak
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|7996,7999|false|false|false|C4283878|Neutrophil Activation Probe Imaging Agent|nap
Finding|Gene or Genome|SIMPLE_SEGMENT|7996,7999|false|false|false|C0870935;C1423800|CTNNBL1 gene;Napping|nap
Finding|Physiologic Function|SIMPLE_SEGMENT|7996,7999|false|false|false|C0870935;C1423800|CTNNBL1 gene;Napping|nap
Finding|Intellectual Product|SIMPLE_SEGMENT|8000,8005|false|false|false|C4050225|Often - answer to question|often
Finding|Gene or Genome|SIMPLE_SEGMENT|8007,8013|false|false|false|C1424587|LITAF gene|Simple
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|8024,8031|false|false|false|C0178629|exhaust|exhaust
Finding|Sign or Symptom|SIMPLE_SEGMENT|8054,8058|false|false|false|C0234233;C1442877|Sore skin;Sore to touch|sore
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8054,8065|false|false|false|C0031350|Pharyngitis|sore throat
Drug|Organic Chemical|SIMPLE_SEGMENT|8054,8065|false|false|false|C0723402;C3244654|Sore Throat brand of Phenol;Sore Throat brand of benzocaine & menthol|sore throat
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8054,8065|false|false|false|C0723402;C3244654|Sore Throat brand of Phenol;Sore Throat brand of benzocaine & menthol|sore throat
Finding|Sign or Symptom|SIMPLE_SEGMENT|8054,8065|false|false|false|C0242429|Sore Throat|sore throat
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8059,8065|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8059,8065|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8059,8065|false|false|false|C1950455|Throat Homeopathic Medication|throat
Finding|Body Substance|SIMPLE_SEGMENT|8059,8065|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Finding|Intellectual Product|SIMPLE_SEGMENT|8059,8065|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Finding|Functional Concept|SIMPLE_SEGMENT|8079,8083|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Finding|Gene or Genome|SIMPLE_SEGMENT|8079,8083|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8102,8108|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8102,8108|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8102,8108|false|false|false|C1950455|Throat Homeopathic Medication|throat
Finding|Body Substance|SIMPLE_SEGMENT|8102,8108|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Finding|Intellectual Product|SIMPLE_SEGMENT|8102,8108|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Finding|Finding|SIMPLE_SEGMENT|8120,8127|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|8120,8127|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|8120,8127|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8120,8127|false|false|false|C0543467|Operative Surgical Procedures|surgery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8135,8141|false|false|false|C0021853|Intestines|BOWELS
Finding|Sign or Symptom|SIMPLE_SEGMENT|8145,8157|false|false|false|C0009806|Constipation|Constipation
Finding|Functional Concept|SIMPLE_SEGMENT|8163,8169|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Finding|Intellectual Product|SIMPLE_SEGMENT|8163,8169|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Finding|Pathologic Function|SIMPLE_SEGMENT|8170,8181|false|false|false|C0879626|Adverse effects|side effect
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|8185,8193|false|false|false|C0027415|Narcotics|narcotic
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8185,8193|false|false|false|C0027415|Narcotics|narcotic
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8194,8198|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|8194,8198|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|8194,8198|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|8194,8207|false|false|false|C0002771|Analgesics|pain medicine
Drug|Organic Chemical|SIMPLE_SEGMENT|8194,8207|false|false|false|C0002771|Analgesics|pain medicine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8194,8207|false|false|false|C0002771|Analgesics|pain medicine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8199,8207|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Drug|Organic Chemical|SIMPLE_SEGMENT|8217,8226|false|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8217,8226|false|false|false|C0030049|oxycodone|oxycodone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8217,8226|false|false|false|C0524222|Oxycodone measurement|oxycodone
Finding|Body Substance|SIMPLE_SEGMENT|8254,8259|false|false|false|C0015733|Feces|stool
Drug|Organic Chemical|SIMPLE_SEGMENT|8254,8268|false|false|false|C0301470;C1154263|Stool Softener;Stool Softener brand of docusate sodium|stool softener
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8254,8268|false|false|false|C0301470;C1154263|Stool Softener;Stool Softener brand of docusate sodium|stool softener
Drug|Organic Chemical|SIMPLE_SEGMENT|8279,8285|false|false|false|C0282139|Colace|Colace
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8279,8285|false|false|false|C0282139|Colace|Colace
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8291,8298|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|8291,8298|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8291,8298|false|false|false|C0006935|capsule (pharmacologic)|capsule
Drug|Organic Chemical|SIMPLE_SEGMENT|8303,8309|false|false|false|C0720654|Gentle|gentle
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8303,8309|false|false|false|C0720654|Gentle|gentle
Drug|Organic Chemical|SIMPLE_SEGMENT|8303,8318|false|false|false|C0720655|Gentle Laxative|gentle laxative
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8303,8318|false|false|false|C0720655|Gentle Laxative|gentle laxative
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8310,8318|false|false|false|C0282090|Laxatives|laxative
Drug|Food|SIMPLE_SEGMENT|8328,8332|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|milk
Drug|Immunologic Factor|SIMPLE_SEGMENT|8328,8332|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|milk
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8328,8332|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|milk
Drug|Substance|SIMPLE_SEGMENT|8328,8332|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|milk
Finding|Body Substance|SIMPLE_SEGMENT|8328,8332|false|false|false|C0026131;C1546713|Milk (body substance);Milk Specimen Code|milk
Finding|Intellectual Product|SIMPLE_SEGMENT|8328,8332|false|false|false|C0026131;C1546713|Milk (body substance);Milk Specimen Code|milk
Drug|Inorganic Chemical|SIMPLE_SEGMENT|8337,8345|false|false|false|C0024477|magnesium oxide|magnesia
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8337,8345|false|false|false|C0024477|magnesium oxide|magnesia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8349,8352|false|false|false|C0265246|Townes syndrome|tbs
Finding|Finding|SIMPLE_SEGMENT|8349,8352|false|false|false|C1419808;C5780809;C5958753|SALL1 gene;SALL1 wt Allele;Toxicity Burden Score|tbs
Finding|Gene or Genome|SIMPLE_SEGMENT|8349,8352|false|false|false|C1419808;C5780809;C5958753|SALL1 gene;SALL1 wt Allele;Toxicity Burden Score|tbs
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8349,8352|false|false|false|C5889868|theta-burst stimulation|tbs
Finding|Idea or Concept|SIMPLE_SEGMENT|8362,8365|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|8362,8365|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8394,8403|false|false|false|C0013227|Pharmaceutical Preparations|medicines
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8414,8426|true|false|false|C5886759|Prescription (attribute)|prescription
Finding|Intellectual Product|SIMPLE_SEGMENT|8414,8426|true|false|false|C1521941|prescription document|prescription
Procedure|Health Care Activity|SIMPLE_SEGMENT|8414,8426|true|false|false|C0033080|Prescription (procedure)|prescription
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8459,8464|false|false|false|C0021853|Intestines|bowel
Finding|Organism Function|SIMPLE_SEGMENT|8459,8473|true|false|false|C0011135|Defecation|bowel movement
Finding|Organism Function|SIMPLE_SEGMENT|8465,8473|true|false|false|C0026649|Movement|movement
Finding|Intellectual Product|SIMPLE_SEGMENT|8478,8487|false|false|false|C2984058|Have Pain|have pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8483,8487|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|8483,8487|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|8483,8487|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8500,8506|false|false|false|C0021853|Intestines|bowels
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8518,8525|false|false|false|C5444295||surgeon
Event|Activity|SIMPLE_SEGMENT|8540,8550|false|false|false|C3241922|Operation Activity|operations
Finding|Functional Concept|SIMPLE_SEGMENT|8540,8550|false|false|false|C0038895;C3244305;C3244306|ActInformationPrivacyReason - operations;HL7PublishingSubSection - operations;Surgical aspects|operations
Finding|Intellectual Product|SIMPLE_SEGMENT|8540,8550|false|false|false|C0038895;C3244305;C3244306|ActInformationPrivacyReason - operations;HL7PublishingSubSection - operations;Surgical aspects|operations
Finding|Finding|SIMPLE_SEGMENT|8552,8560|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|8552,8560|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Finding|SIMPLE_SEGMENT|8584,8592|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|8584,8592|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Drug|Organic Chemical|SIMPLE_SEGMENT|8605,8618|false|false|false|C0718564|Anti-Diarrhea|anti-diarrhea
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8605,8618|false|false|false|C0718564|Anti-Diarrhea|anti-diarrhea
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8619,8628|false|false|false|C0013227|Pharmaceutical Preparations|medicines
Drug|Substance|SIMPLE_SEGMENT|8647,8653|false|false|false|C0302908|Liquid substance|fluids
Finding|Body Substance|SIMPLE_SEGMENT|8647,8653|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8647,8653|false|false|false|C0016286|Fluid Therapy|fluids
Finding|Finding|SIMPLE_SEGMENT|8710,8716|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|8710,8716|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|8725,8733|false|false|false|C0231218;C0557911;C2987492|Feel Ill Question;Feeling bad emotionally;Malaise|feel ill
Finding|Sign or Symptom|SIMPLE_SEGMENT|8725,8733|false|false|false|C0231218;C0557911;C2987492|Feel Ill Question;Feeling bad emotionally;Malaise|feel ill
Finding|Sign or Symptom|SIMPLE_SEGMENT|8730,8733|false|false|false|C0231218|Malaise|ill
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8752,8759|false|false|false|C5444295||surgeon
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8762,8766|false|false|false|C2598155||PAIN
Finding|Functional Concept|SIMPLE_SEGMENT|8762,8766|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|PAIN
Finding|Sign or Symptom|SIMPLE_SEGMENT|8762,8766|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|PAIN
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8762,8777|false|false|false|C0002766|Pain management (procedure)|PAIN MANAGEMENT
Event|Occupational Activity|SIMPLE_SEGMENT|8767,8777|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|MANAGEMENT
Procedure|Health Care Activity|SIMPLE_SEGMENT|8767,8777|false|false|false|C0376636|Disease Management|MANAGEMENT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8813,8825|false|false|false|C5886759|Prescription (attribute)|prescription
Finding|Intellectual Product|SIMPLE_SEGMENT|8813,8825|false|false|false|C1521941|prescription document|prescription
Procedure|Health Care Activity|SIMPLE_SEGMENT|8813,8825|false|false|false|C0033080|Prescription (procedure)|prescription
Drug|Organic Chemical|SIMPLE_SEGMENT|8832,8841|false|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8832,8841|false|false|false|C0030049|oxycodone|oxycodone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8832,8841|false|false|false|C0524222|Oxycodone measurement|oxycodone
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8847,8851|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|8847,8851|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|8847,8851|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|SIMPLE_SEGMENT|8847,8859|false|false|false|C5548091|Demonstrates adequate pain control|pain control
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8847,8859|false|false|false|C0002766;C1304888|Pain control;Pain management (procedure)|pain control
Drug|Organic Chemical|SIMPLE_SEGMENT|8852,8859|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8852,8859|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|SIMPLE_SEGMENT|8852,8859|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Finding|Conceptual Entity|SIMPLE_SEGMENT|8852,8859|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|SIMPLE_SEGMENT|8852,8859|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|SIMPLE_SEGMENT|8852,8859|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Drug|Organic Chemical|SIMPLE_SEGMENT|8874,8881|false|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8874,8881|false|false|false|C0699142|Tylenol|Tylenol
Finding|Finding|SIMPLE_SEGMENT|8967,8974|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|8967,8974|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|8967,8974|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8967,8974|false|false|false|C0543467|Operative Surgical Procedures|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|9002,9010|false|true|false|C0442805|Increase|increase
Finding|Finding|SIMPLE_SEGMENT|9011,9015|false|true|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|9011,9015|false|true|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|9011,9015|false|true|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9053,9057|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9053,9057|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9053,9057|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|9105,9114|false|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9105,9114|false|false|false|C0030049|oxycodone|oxycodone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9105,9114|false|false|false|C0524222|Oxycodone measurement|oxycodone
Finding|Finding|SIMPLE_SEGMENT|9119,9127|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|9119,9127|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Finding|SIMPLE_SEGMENT|9132,9138|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|9132,9138|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Finding|SIMPLE_SEGMENT|9132,9143|false|false|false|C0278140;C4050465;C4521229|Neck Pain Score 6;Severe Extremity Pain;Severe pain|severe pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9139,9143|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9139,9143|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9139,9143|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|9167,9174|false|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9167,9174|false|false|false|C0699142|Tylenol|Tylenol
Finding|Body Substance|SIMPLE_SEGMENT|9191,9196|false|false|false|C0015733|Feces|stool
Drug|Organic Chemical|SIMPLE_SEGMENT|9191,9205|false|false|false|C0301470;C1154263|Stool Softener;Stool Softener brand of docusate sodium|stool softener
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9191,9205|false|false|false|C0301470;C1154263|Stool Softener;Stool Softener brand of docusate sodium|stool softener
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|9215,9224|false|false|false|C0027415|Narcotics|narcotics
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9215,9224|false|false|false|C0027415|Narcotics|narcotics
Finding|Sign or Symptom|SIMPLE_SEGMENT|9246,9258|false|false|false|C0009806|Constipation|constipation
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9303,9314|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9303,9314|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|SIMPLE_SEGMENT|9303,9314|false|false|false|C4284232|Medications|medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9337,9341|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9337,9341|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9337,9341|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Idea or Concept|SIMPLE_SEGMENT|9353,9359|false|false|false|C1550462|Observation Interpretation - better|better
Finding|Idea or Concept|SIMPLE_SEGMENT|9360,9363|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|9360,9363|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Idea or Concept|SIMPLE_SEGMENT|9367,9370|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|9367,9370|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9388,9392|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9388,9392|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9388,9392|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|SIMPLE_SEGMENT|9405,9410|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Idea or Concept|SIMPLE_SEGMENT|9405,9410|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Idea or Concept|SIMPLE_SEGMENT|9422,9428|false|false|false|C1550462|Observation Interpretation - better|better
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9450,9457|false|false|false|C5444295||surgeon
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9521,9528|false|false|false|C5444295||surgeon
Finding|Finding|SIMPLE_SEGMENT|9533,9538|false|false|false|C1444775;C1539835;C3890003|SPEN gene;SPEN wt Allele;Sharp sensation quality|sharp
Finding|Gene or Genome|SIMPLE_SEGMENT|9533,9538|false|false|false|C1444775;C1539835;C3890003|SPEN gene;SPEN wt Allele;Sharp sensation quality|sharp
Finding|Sign or Symptom|SIMPLE_SEGMENT|9533,9543|false|false|false|C0455270|Sharp pain|sharp pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9539,9543|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9539,9543|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9539,9543|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|SIMPLE_SEGMENT|9551,9557|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|9551,9557|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Finding|SIMPLE_SEGMENT|9551,9562|false|false|false|C0278140;C4050465;C4521229|Neck Pain Score 6;Severe Extremity Pain;Severe pain|severe pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9558,9562|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9558,9562|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9558,9562|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9590,9595|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|9590,9595|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9590,9600|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9590,9600|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9596,9600|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9596,9600|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9596,9600|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|SIMPLE_SEGMENT|9602,9610|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|9602,9610|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|9602,9610|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|9602,9610|false|false|false|C0033095||pressure
Drug|Organic Chemical|SIMPLE_SEGMENT|9638,9643|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9638,9643|false|false|false|C3815497|Cough (guaifenesin)|cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|9638,9643|false|false|false|C0010200|Coughing|cough
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9645,9664|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|SIMPLE_SEGMENT|9645,9664|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|SIMPLE_SEGMENT|9658,9664|false|false|false|C0225386|Breath|breath
Finding|Sign or Symptom|SIMPLE_SEGMENT|9666,9674|false|false|false|C0043144|Wheezing|wheezing
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9677,9681|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9677,9681|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9677,9681|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|SIMPLE_SEGMENT|9698,9703|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Idea or Concept|SIMPLE_SEGMENT|9698,9703|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Finding|SIMPLE_SEGMENT|9709,9713|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|9709,9713|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|9709,9713|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9717,9721|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9717,9721|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9717,9721|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|SIMPLE_SEGMENT|9727,9732|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|9727,9732|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|9743,9749|false|false|false|C0085593|Chills|chills
Finding|Finding|SIMPLE_SEGMENT|9751,9756|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|9751,9756|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Functional Concept|SIMPLE_SEGMENT|9786,9792|false|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9786,9792|false|false|false|C4319952|Change - procedure|change
Finding|Functional Concept|SIMPLE_SEGMENT|9786,9795|false|false|false|C0392747|Changing|change in
Finding|Functional Concept|SIMPLE_SEGMENT|9796,9802|false|false|false|C0349590;C1262865|Nature;Natures|nature
Finding|Idea or Concept|SIMPLE_SEGMENT|9796,9802|false|false|false|C0349590;C1262865|Nature;Natures|nature
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9822,9826|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9822,9826|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9822,9826|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9829,9835|false|false|false|C4255480||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|9829,9835|false|false|false|C0027497|Nausea|nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|9829,9848|false|false|false|C0027498|Nausea and vomiting|nausea and vomiting
Finding|Sign or Symptom|SIMPLE_SEGMENT|9840,9848|false|false|false|C0042963|Vomiting|vomiting
Drug|Substance|SIMPLE_SEGMENT|9872,9878|false|false|false|C0302908|Liquid substance|fluids
Finding|Body Substance|SIMPLE_SEGMENT|9872,9878|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9872,9878|false|false|false|C0016286|Fluid Therapy|fluids
Drug|Food|SIMPLE_SEGMENT|9880,9884|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Drug|Immunologic Factor|SIMPLE_SEGMENT|9880,9884|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9880,9884|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9895,9906|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9895,9906|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|SIMPLE_SEGMENT|9895,9906|false|false|false|C4284232|Medications|medications
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9928,9938|false|false|false|C0011175|Dehydration|dehydrated
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9940,9949|false|false|false|C0043352|Xerostomia|dry mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9944,9949|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|9944,9949|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Finding|SIMPLE_SEGMENT|9951,9967|false|false|false|C0039231|Tachycardia|rapid heart beat
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9957,9962|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|9957,9962|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|9957,9962|false|false|false|C0795691|HEART PROBLEM|heart
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|9957,9967|false|false|false|C0425583|Heart beat|heart beat
Finding|Sign or Symptom|SIMPLE_SEGMENT|9970,9983|false|false|false|C0849959|feeling dizzy|feeling dizzy
Finding|Sign or Symptom|SIMPLE_SEGMENT|9978,9983|false|false|false|C0012833|Dizziness|dizzy
Finding|Finding|SIMPLE_SEGMENT|9987,9992|false|false|false|C0039070;C4554554|Faint - appearance;Syncope|faint
Finding|Sign or Symptom|SIMPLE_SEGMENT|9987,9992|false|false|false|C0039070;C4554554|Faint - appearance;Syncope|faint
Finding|Functional Concept|SIMPLE_SEGMENT|10025,10031|false|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10025,10031|false|false|false|C4319952|Change - procedure|change
Finding|Functional Concept|SIMPLE_SEGMENT|10025,10034|false|false|false|C0392747|Changing|change in
Finding|Functional Concept|SIMPLE_SEGMENT|10040,10048|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|10040,10048|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|10056,10064|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|10056,10064|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|10083,10093|false|false|false|C1524062|Additional|Additional
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10099,10103|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|10099,10103|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|10099,10103|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|SIMPLE_SEGMENT|10120,10125|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Idea or Concept|SIMPLE_SEGMENT|10120,10125|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Finding|SIMPLE_SEGMENT|10131,10135|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|10131,10135|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|10131,10135|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10154,10159|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|10154,10159|false|false|false|C0741025|Chest problem|chest
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10172,10179|false|false|false|C0042027|Urinary tract|urinary
Finding|Sign or Symptom|SIMPLE_SEGMENT|10182,10189|false|false|false|C0085624|Burning sensation|burning
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10193,10198|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|SIMPLE_SEGMENT|10193,10198|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Body Substance|SIMPLE_SEGMENT|10207,10212|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|SIMPLE_SEGMENT|10207,10212|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|SIMPLE_SEGMENT|10207,10212|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10243,10254|false|false|false|C0802604;C2598133||MEDICATIONS
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10243,10254|false|false|false|C0013227|Pharmaceutical Preparations|MEDICATIONS
Finding|Intellectual Product|SIMPLE_SEGMENT|10243,10254|false|false|false|C4284232|Medications|MEDICATIONS
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10271,10280|false|false|false|C0013227|Pharmaceutical Preparations|medicines
Event|Activity|SIMPLE_SEGMENT|10304,10313|false|false|false|C3241922|Operation Activity|operation
Procedure|Machine Activity|SIMPLE_SEGMENT|10304,10313|false|false|false|C0543467;C1880161|Computer Operation;Operative Surgical Procedures|operation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10304,10313|false|false|false|C0543467;C1880161|Computer Operation;Operative Surgical Procedures|operation
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10417,10425|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Procedure|Health Care Activity|SIMPLE_SEGMENT|10445,10449|false|false|false|C1515187|Take|take
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10468,10475|false|false|false|C5444295||surgeon
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|10479,10484|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|WOUND
Finding|Body Substance|SIMPLE_SEGMENT|10479,10484|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|WOUND
Finding|Functional Concept|SIMPLE_SEGMENT|10479,10484|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|WOUND
Finding|Intellectual Product|SIMPLE_SEGMENT|10479,10484|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|WOUND
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10479,10489|false|false|false|C0886052;C1272654|Wound care management;wound care|WOUND CARE
Event|Activity|SIMPLE_SEGMENT|10485,10489|false|false|false|C1947933|care activity|CARE
Finding|Finding|SIMPLE_SEGMENT|10485,10489|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|CARE
Finding|Intellectual Product|SIMPLE_SEGMENT|10485,10489|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|CARE
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10494,10502|false|false|false|C1705365|Dressing Dosage Form|dressing
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|10494,10502|false|false|false|C0518459;C1305428|Ability to dress|dressing
Finding|Finding|SIMPLE_SEGMENT|10494,10502|false|false|false|C0518459;C1305428|Ability to dress|dressing
Procedure|Health Care Activity|SIMPLE_SEGMENT|10494,10502|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10494,10502|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Event|Activity|SIMPLE_SEGMENT|10503,10510|false|false|false|C1883720|Removing (action)|removal
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10503,10510|false|false|false|C0015252;C0185115;C0728940|Excision;Extraction;removal technique|removal
Finding|Idea or Concept|SIMPLE_SEGMENT|10579,10582|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|10579,10582|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10592,10599|false|false|false|C2346961|Bandage Dosage Form|bandage
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|10673,10677|false|false|false|C0039003|Swimming|swim
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10683,10686|false|false|false|C0030587|Paroxysmal atrial tachycardia|pat
Drug|Organic Chemical|SIMPLE_SEGMENT|10683,10686|false|false|false|C2825250|Fenamole|pat
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10683,10686|false|false|false|C2825250|Fenamole|pat
Finding|Molecular Function|SIMPLE_SEGMENT|10683,10686|false|false|false|C2247344;C2247346;C2248827|aspartate-prephenate aminotransferase activity;glutamate-prephenate aminotransferase activity;protein acetyltransferase activity|pat
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10683,10686|false|false|false|C3897364|Thermoacoustic Computed Tomography|pat
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10692,10700|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|10692,10700|false|false|false|C0332803|Surgical wound|incision
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10692,10700|false|false|false|C0184898|Surgical incisions|incision
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10791,10796|false|false|false|C1410088|Still|still
Procedure|Health Care Activity|SIMPLE_SEGMENT|10890,10895|false|false|false|C0150141|Bathing|baths
Finding|Functional Concept|SIMPLE_SEGMENT|10897,10901|false|false|false|C1549544|Soak Administration|soak
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10897,10901|false|false|false|C0204774|Soak (procedure)|soak
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|10906,10910|false|false|false|C0039003|Swimming|swim
Finding|Finding|SIMPLE_SEGMENT|10923,10936|false|false|false|C0241311|post operative (finding)|after surgery
Finding|Finding|SIMPLE_SEGMENT|10929,10936|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|10929,10936|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|10929,10936|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10929,10936|false|false|false|C0543467|Operative Surgical Procedures|surgery
Procedure|Health Care Activity|SIMPLE_SEGMENT|10968,10976|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10968,10976|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10997,11004|false|false|false|C5444295||surgeon
Finding|Finding|SIMPLE_SEGMENT|11019,11027|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Finding|Idea or Concept|SIMPLE_SEGMENT|11019,11027|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Finding|Organism Function|SIMPLE_SEGMENT|11034,11042|false|false|false|C0037361|Smell Perception|smelling
Finding|Finding|SIMPLE_SEGMENT|11045,11051|false|false|false|C4554530|Bloody|bloody
Drug|Substance|SIMPLE_SEGMENT|11053,11056|false|false|false|C0444185|Pus specimen|pus
Finding|Body Substance|SIMPLE_SEGMENT|11053,11056|false|false|false|C0034161;C1546758|Pus;Pus Specimen Code|pus
Finding|Intellectual Product|SIMPLE_SEGMENT|11053,11056|false|false|false|C0034161;C1546758|Pus;Pus Specimen Code|pus
Finding|Idea or Concept|SIMPLE_SEGMENT|11058,11061|false|false|false|C1548556|Etc.|etc
Finding|Body Substance|SIMPLE_SEGMENT|11076,11084|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|SIMPLE_SEGMENT|11076,11084|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11076,11084|false|false|false|C0013103|Drainage procedure|drainage
Anatomy|Body Location or Region|SIMPLE_SEGMENT|11095,11103|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|11095,11103|false|false|false|C0332803|Surgical wound|incision
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11095,11103|false|false|false|C0184898|Surgical incisions|incision
Anatomy|Body Location or Region|SIMPLE_SEGMENT|11104,11108|false|false|false|C1515974|Anatomic Site|site
Finding|Intellectual Product|SIMPLE_SEGMENT|11104,11108|false|false|false|C1546778||site
Anatomy|Body Location or Region|SIMPLE_SEGMENT|11127,11135|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|11127,11135|false|false|false|C0332803|Surgical wound|incision
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11127,11135|false|false|false|C0184898|Surgical incisions|incision
Finding|Finding|SIMPLE_SEGMENT|11140,11149|false|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Functional Concept|SIMPLE_SEGMENT|11140,11149|false|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Sign or Symptom|SIMPLE_SEGMENT|11140,11154|false|false|false|C5141269|Increased pain|increased pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11150,11154|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|11150,11154|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|11150,11154|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|11158,11166|false|false|false|C0009938|Contusions|bruising
Finding|Finding|SIMPLE_SEGMENT|11158,11166|false|false|false|C2136686|reported bruising (history)|bruising
Finding|Finding|SIMPLE_SEGMENT|11179,11184|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|11179,11184|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11188,11197|false|false|false|C0009450|Communicable Diseases|infection
Finding|Pathologic Function|SIMPLE_SEGMENT|11188,11197|false|false|false|C3714514|Infection|infection
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11206,11213|false|false|false|C0041834|Erythema|redness
Finding|Finding|SIMPLE_SEGMENT|11206,11213|false|false|false|C0332575|Redness|redness
Anatomy|Body System|SIMPLE_SEGMENT|11233,11237|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11233,11237|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|11233,11237|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Finding|Body Substance|SIMPLE_SEGMENT|11233,11237|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|SIMPLE_SEGMENT|11233,11237|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Finding|SIMPLE_SEGMENT|11240,11248|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|11240,11248|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Finding|SIMPLE_SEGMENT|11250,11259|false|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Functional Concept|SIMPLE_SEGMENT|11250,11259|false|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Sign or Symptom|SIMPLE_SEGMENT|11250,11264|false|false|false|C5141269|Increased pain|increased pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11260,11264|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|11260,11264|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|11260,11264|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Body Substance|SIMPLE_SEGMENT|11279,11287|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|SIMPLE_SEGMENT|11279,11287|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11279,11287|false|false|false|C0013103|Drainage procedure|drainage
Event|Activity|SIMPLE_SEGMENT|11385,11389|false|false|false|C1947933|care activity|care
Finding|Finding|SIMPLE_SEGMENT|11385,11389|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|11385,11389|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Idea or Concept|SIMPLE_SEGMENT|11438,11442|false|false|false|C0376558|Life|life
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|11438,11442|false|false|false|C1522684|Laser-Induced Fluorescence Endoscopy|life
Event|Activity|SIMPLE_SEGMENT|11447,11457|false|false|false|C0441655|Activities|activities
Finding|Finding|SIMPLE_SEGMENT|11447,11457|false|false|false|C2239122|activities (history)|activities
Finding|Idea or Concept|SIMPLE_SEGMENT|11460,11464|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|11460,11464|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|11460,11464|false|false|false|C1553498|home health encounter|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|11491,11499|false|false|false|C1546572||catheter
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11508,11515|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|11508,11515|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11508,11515|false|false|false|C0872388|Procedures on bladder|bladder
Finding|Idea or Concept|SIMPLE_SEGMENT|11542,11545|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|11542,11545|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Finding|SIMPLE_SEGMENT|11554,11561|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|11554,11561|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|11554,11561|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11554,11561|false|false|false|C0543467|Operative Surgical Procedures|surgery
Finding|Finding|SIMPLE_SEGMENT|11568,11578|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Finding|Intellectual Product|SIMPLE_SEGMENT|11617,11625|false|false|false|C1546572||catheter
Event|Activity|SIMPLE_SEGMENT|11637,11648|false|false|false|C0003629|Appointments|appointment
Finding|Idea or Concept|SIMPLE_SEGMENT|11690,11696|false|false|false|C1554106|MDF AttributeType - Number|number
Event|Activity|SIMPLE_SEGMENT|11721,11732|false|false|false|C0003629|Appointments|appointment
Event|Event|SIMPLE_SEGMENT|11776,11783|false|false|false|C1516084|Attempt|attempt
Finding|Finding|SIMPLE_SEGMENT|11817,11821|false|false|false|C1299581|Able (qualifier value)|able
Finding|Functional Concept|SIMPLE_SEGMENT|11832,11837|false|false|false|C5848602|Exhausted|Empty
Finding|Intellectual Product|SIMPLE_SEGMENT|11842,11845|false|false|false|C1552710|Bag Data Type|bag
Finding|Organism Function|SIMPLE_SEGMENT|11879,11886|false|false|false|C0006147|Breast Feeding|nursing
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11879,11886|false|false|false|C0028678|RNAx nursing therapy actions|nursing
Finding|Finding|SIMPLE_SEGMENT|11887,11892|false|false|false|C1551040|Encounter Special Courtesy - staff|staff
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11915,11918|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Intellectual Product|SIMPLE_SEGMENT|11919,11922|false|false|false|C1552710|Bag Data Type|bag
Finding|Body Substance|SIMPLE_SEGMENT|11935,11944|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|11935,11944|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|11935,11944|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|11935,11944|false|false|false|C0030685|Patient Discharge|discharge
Finding|Functional Concept|SIMPLE_SEGMENT|11960,11963|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|SIMPLE_SEGMENT|11960,11963|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|11974,11979|false|false|false|C0221188|Tripping|trips
Finding|Intellectual Product|SIMPLE_SEGMENT|11999,12002|false|false|false|C1552710|Bag Data Type|bag
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12024,12027|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Idea or Concept|SIMPLE_SEGMENT|12037,12041|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|12037,12041|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|12037,12041|false|false|false|C1553498|home health encounter|home
Finding|Idea or Concept|SIMPLE_SEGMENT|12086,12090|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|12086,12090|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|12086,12090|false|false|false|C1553498|home health encounter|home
Finding|Intellectual Product|SIMPLE_SEGMENT|12113,12119|false|false|false|C1561574|Amount class - Amount|amount
Finding|Intellectual Product|SIMPLE_SEGMENT|12129,12132|false|false|false|C1552710|Bag Data Type|bag
Finding|Intellectual Product|SIMPLE_SEGMENT|12179,12184|false|false|false|C4050225|Often - answer to question|often
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12232,12235|false|false|false|C4522181|Brachial Amyotrophic Diplegia|bad
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12232,12235|false|false|false|C1530798|BAD protein, human|bad
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12232,12235|false|false|false|C1530798|BAD protein, human|bad
Finding|Gene or Genome|SIMPLE_SEGMENT|12232,12235|false|false|false|C1366450|BAD gene|bad
Finding|Finding|SIMPLE_SEGMENT|12250,12257|false|false|false|C4534363|At home|at home
Finding|Idea or Concept|SIMPLE_SEGMENT|12253,12257|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|12253,12257|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|12253,12257|false|false|false|C1553498|home health encounter|home
Event|Activity|SIMPLE_SEGMENT|12295,12299|false|false|false|C1947933|care activity|Care
Finding|Finding|SIMPLE_SEGMENT|12295,12299|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|SIMPLE_SEGMENT|12295,12299|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12295,12304|false|false|false|C4321316||Care Team
Finding|Finding|SIMPLE_SEGMENT|12295,12304|false|false|false|C4321315|Care team|Care Team
Procedure|Health Care Activity|SIMPLE_SEGMENT|12307,12315|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12316,12328|false|false|false|C3263700||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|12316,12328|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

