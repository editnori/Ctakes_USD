CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Neurology speciality|Title|false|false||NEUROLOGYnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Known|Modifier|false|false||Knownnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Adverse reaction to drug|Finding|true|false||Adverse Drug Reactionsnull|Adverse reaction to drug|Finding|true|false||Drug Reactionsnull|Pharmaceutical Preparations|Drug|false|false||Drug
null|Pharmacologic Substance|Drug|false|false||Drugnull|Drug problem|Finding|false|false||Drugnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Chief complaint (finding)|Finding|false|false||Chief Complaintnull|Complaint (finding)|Finding|false|false||Complaintnull|null|Attribute|false|false||Complaintnull|Speech|Finding|false|false||speechnull|Speech assessment|Procedure|false|false||speechnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|History of present illness (finding)|Finding|false|false||History of Present Illnessnull|null|Attribute|false|false||History of Present Illnessnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Present illness|Finding|false|false||Present Illnessnull|Present|Finding|false|false||Present
null|Presentation|Finding|false|false||Presentnull|Illness (finding)|Finding|false|false||Illnessnull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Old|Time|false|false||oldnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Woman|Subject|false|false||woman
null|Human, Female adult|Subject|false|false||womannull|Atrial Fibrillation|Disorder|false|false||Atrial fibrillationnull|null|Attribute|false|false||Atrial fibrillationnull|Atrial Fibrillation by ECG Finding|Lab|false|false||Atrial fibrillationnull|Heart Atrium|Anatomy|false|false||Atrialnull|Fibrillation|Disorder|false|false||fibrillationnull|Eliquis|Drug|false|false||Eliquis
null|Eliquis|Drug|false|false||Eliquisnull|Once daily|Time|false|false||once dailynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Daily|Time|false|false||dailynull|Hypertensive disease|Disorder|false|false||hypertensionnull|Hyperlipidemia|Disorder|false|false||hyperlipidemia
null|Hyperlipoproteinemias|Disorder|false|false||hyperlipidemianull|Serum lipids high (finding)|Finding|false|false||hyperlipidemianull|Congestive heart failure|Disorder|false|false||CHFnull|Choroidal fissure|Anatomy|false|false||CHFnull|Transfer - product ownership|Finding|false|false||transfer
null|Transfer Technique|Finding|false|false||transfer
null|ActClass - transfer|Finding|false|false||transfer
null|null|Finding|false|false||transfernull|Transfer (immobility management)|Procedure|false|false||transfernull|Sudden onset (contextual qualifier) (qualifier value)|Finding|false|false||acute onsetnull|Sudden onset (attribute)|Time|false|false||acute onset
null|acute|Time|false|false||acute onsetnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Onset of (contextual qualifier)|Modifier|false|false||onsetnull|Age of Onset|LabModifier|false|false||onsetnull|Dysarthria|Disorder|false|false||dysarthrianull|Cancer/Testis Antigen|Drug|false|false||CTAnull|PCYT1A wt Allele|Finding|false|false||CTA
null|CERNA3 gene|Finding|false|false||CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false||CTAnull|Possible|Finding|false|false||possiblenull|Possible diagnosis|Modifier|false|false||possible
null|Possibly Related to Intervention|Modifier|false|false||possiblenull|Target Awareness - partial|Finding|false|false||partialnull|Partial|LabModifier|false|false||partialnull|Thrombus|Finding|false|false||thrombus
null|Blood Clot|Finding|false|false||thrombusnull|Thrombus <Thrombidae>|Entity|false|false||thrombusnull|Stenosis|Finding|false|false||stenosisnull|Stenosis <Pimeliinae>|Entity|false|false||stenosisnull|Stenosis Morphology|Modifier|false|false||stenosisnull|Upper|Modifier|false|false||superiornull|Organization Unit Type - Division|Finding|false|false||divisionnull|Division (surgical procedure)|Procedure|false|false||division
null|Transection (procedure)|Procedure|false|false||divisionnull|Division (action)|Event|false|false||divisionnull|Administrative Division|Entity|false|false||divisionnull|Preventive monitoring|Procedure|false|false||monitoringnull|null|Event|false|false||monitoringnull|Possible|Finding|false|false||possiblenull|Possible diagnosis|Modifier|false|false||possible
null|Possibly Related to Intervention|Modifier|false|false||possiblenull|Thrombectomy|Procedure|false|false||thrombectomynull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Daughter|Subject|false|false||daughternull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Excellent - LanguageAbilityProficiency|Modifier|false|false||excellent
null|Excellent - Specimen Quality|Modifier|false|false||excellent
null|Excellent (qualifier value)|Modifier|false|false||excellentnull|Historian|Subject|false|false||historiannull|Dinner|Finding|false|false||dinnernull|With dinner|Time|false|false||dinnernull|Friends (Religious Affiliation)|Subject|false|false||friends
null|friend|Subject|false|false||friendsnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Residential flat|Device|false|false||apartmentnull|Computers|Device|false|false||computernull|Last|Modifier|false|false||Lastnull|Known|Modifier|false|false||knownnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Then - dosing instruction fragment|Finding|false|false||Thennull|Then|Time|false|false||Thennull|Oppositional Defiant Disorder|Disorder|false|false||oddnull|GJA1 gene|Finding|false|false||odd
null|OSR1 gene|Finding|false|false||oddnull|Observation of Sensation|Finding|false|false||sensation
null|Sensory perception|Finding|false|false||sensationnull|sensory exam|Procedure|false|false||sensationnull|Sensation quality|Modifier|false|false||sensationnull|Alveolar rhabdomyosarcoma|Disorder|false|false||armsnull|Adherence to Refills and Medications Scale|Finding|false|false||arms
null|KIDINS220 gene|Finding|false|false||armsnull|Upper arm|Anatomy|false|false||armsnull|null|Attribute|false|false||armsnull|Room - Patient location type|Modifier|false|false||room
null|Room|Modifier|false|false||roomnull|Very|Modifier|false|false||verynull|Then - dosing instruction fragment|Finding|false|false||Thennull|Then|Time|false|false||Thennull|Family member|Subject|false|false||family membersnull|Entity Name Part Type - family|Finding|false|false||family
null|Last Name|Finding|false|false||family
null|Living Arrangement - Family|Finding|false|false||family
null|Family (taxonomic)|Finding|false|false||family
null|Family Collection|Finding|false|false||familynull|Family|Subject|false|false||familynull|member|Subject|false|false||membersnull|Door (physical object)|Device|false|false||doornull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Open|Modifier|false|false||opennull|Door (physical object)|Device|false|false||doornull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|RXFP2 gene|Finding|false|false||greatnull|Greater|LabModifier|false|false||great
null|Large|LabModifier|false|false||greatnull|Has difficulty doing (qualifier value)|Finding|false|false||difficultynull|Walkers|Device|false|false||walkernull|Usually|Finding|false|false||usuallynull|Usual|Modifier|false|false||usuallynull|Walkers|Device|false|false||walkernull|Knee Replacement Arthroplasty|Procedure|false|false||knee replacementnull|null|Attribute|false|false||knee replacementnull|Examination of knee joint|Procedure|false|false||kneenull|Knee region structure|Anatomy|false|false||knee
null|Knee|Anatomy|false|false||knee
null|Lower extremity>Knee|Anatomy|false|false||knee
null|Knee joint|Anatomy|false|false||kneenull|Replacement|Finding|false|false||replacementnull|Replacement - supply|Procedure|false|false||replacement
null|Surgical Replantation|Procedure|false|false||replacementnull|Chairs|Device|false|false||chairnull|Chairperson|Subject|false|false||chairnull|Walkers|Device|false|false||walkernull|Door (physical object)|Device|false|false||doornull|Unlock|Finding|false|false||unlocknull|Problems - What subject filter|Finding|false|false||problemsnull|Family member|Subject|false|false||family membersnull|Entity Name Part Type - family|Finding|false|false||family
null|Last Name|Finding|false|false||family
null|Living Arrangement - Family|Finding|false|false||family
null|Family (taxonomic)|Finding|false|false||family
null|Family Collection|Finding|false|false||familynull|Family|Subject|false|false||familynull|member|Subject|false|false||membersnull|Has difficulty doing (qualifier value)|Finding|false|false||difficultynull|Term (lexical)|Finding|false|false||wordnull|Experimental Finding|Finding|true|false||finding
null|Signs and Symptoms|Finding|true|false||finding
null|Finding|Finding|true|false||findingnull|Has difficulty doing (qualifier value)|Finding|false|false||difficultynull|Person Info|Finding|false|false||personnull|null|Attribute|false|false||personnull|Persons|Subject|false|false||personnull|Too much|Finding|false|false||too muchnull|Much|Finding|false|false||muchnull|Very|Modifier|false|false||verynull|Awareness|Finding|false|false||awarenull|Dysarthria|Disorder|false|false||dysarthrianull|Daughter|Subject|false|false||daughtersnull|Cerebrovascular accident|Disorder|false|false||strokenull|Stroke (heart beat)|Finding|false|false||strokenull|Then - dosing instruction fragment|Finding|false|false||Thennull|Then|Time|false|false||Thennull|Idea|Entity|true|false||ideanull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|Walkers|Device|false|false||walkernull|Unsteady|Modifier|false|false||unsteadynull|Nearly|Modifier|false|false||almostnull|Visual changes|Finding|true|false||visual changesnull|Visual|Finding|false|false||visualnull|Changing|Finding|true|false||changesnull|Changed status|LabModifier|false|false||changesnull|Numbness|Finding|true|false||numbness
null|Hypesthesia|Finding|true|false||numbnessnull|Paresthesia|Disorder|false|false||tinglingnull|Has tingling sensation|Finding|false|false||tinglingnull|Focal|Modifier|false|false||focalnull|Weakness|Finding|true|false||weakness
null|Asthenia|Finding|true|false||weaknessnull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|Door (physical object)|Device|false|false||doornull|Issue (document)|Finding|true|false||issue
null|Problem|Finding|true|false||issuenull|Issue (action)|Event|true|false||issuenull|Shakes|Finding|false|false||shakynull|Ethyl Methanesulfonate|Drug|false|false||EMS
null|Ethyl Methanesulfonate|Drug|false|false||EMS
null|Ethyl Methanesulfonate|Drug|false|false||EMSnull|EMSLR gene|Finding|false|false||EMSnull|Emergency Medical Services|Procedure|false|false||EMSnull|NIH stroke scale|Finding|false|false||NIHSSnull|Speech|Finding|false|false||speechnull|Speech assessment|Procedure|false|false||speechnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Paramedic (occupation)|Subject|false|false||Paramedicsnull|Speech|Finding|false|false||speechnull|Speech assessment|Procedure|false|false||speechnull|Rapid|Modifier|false|false||rapidlynull|Route|Modifier|false|false||routenull|Past 30 days|Time|false|false||Last monthnull|Last|Modifier|false|false||Lastnull|Transaction counts and value totals - month|Finding|false|false||month
null|Precision - month|Finding|false|false||monthnull|month|Time|false|false||month
null|Monthly (qualifier value)|Time|false|false||monthnull|N-(4-aminophenethyl)spiroperidol|Drug|false|false||napsnull|outcomes otolaryngology hearing|Finding|false|false||hearing
null|Hearing finding|Finding|false|false||hearing
null|Hearing|Finding|false|false||hearingnull|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group|Finding|false|false||poor
null|Patient Condition Code - Poor|Finding|false|false||poornull|Poverty|Subject|false|false||poornull|Language Proficiency - Poor|Modifier|false|false||poor
null|Specimen Quality - Poor|Modifier|false|false||poor
null|Poor - grade|Modifier|false|false||poor
null|Poor - qualifier|Modifier|false|false||poornull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Hearing Aids|Device|false|false||hearing aidsnull|outcomes otolaryngology hearing|Finding|false|false||hearing
null|Hearing finding|Finding|false|false||hearing
null|Hearing|Finding|false|false||hearingnull|Acquired Immunodeficiency Syndrome|Disorder|false|false||aidsnull|month|Time|false|false||monthsnull|Dysuria|Finding|false|false||dysurianull|More|LabModifier|false|false||morenull|Frequent headache|Finding|false|false||frequent headachesnull|Frequently|Time|false|false||frequentnull|Headache|Finding|false|false||headachesnull|month|Time|false|false||monthsnull|Last|Modifier|false|false||Lastnull|Headache|Finding|false|false||headachenull|tramadol|Drug|false|false||tramadol
null|tramadol|Drug|false|false||tramadolnull|Tramadol measurement (procedure)|Procedure|false|false||tramadolnull|Acetaminophen [EPC]|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophennull|Acetaminophen measurement|Procedure|false|false||acetaminophennull|Couple (action)|Finding|false|false||couplenull|Couples (persons)|Subject|false|false||couplenull|Night time|Time|false|false||nightnull|Headache|Finding|false|false||headachesnull|Night time|Time|false|false||at nightnull|Night time|Time|false|false||nightnull|Headache|Finding|false|false||headachenull|positional|Finding|false|false||positionalnull|Gradual|Modifier|false|false||gradualnull|Weight Loss|Finding|false|false||weight loss
null|Losing Weight (question)|Finding|false|false||weight lossnull|Measured weight loss (observable entity)|LabModifier|false|false||weight lossnull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|Loss (adaptation)|Finding|false|false||lossnull|Loss (quantitative)|LabModifier|false|false||lossnull|12 Months|Time|false|false||12 monthsnull|month|Time|false|false||monthsnull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|Nearly|Modifier|false|false||almostnull|liquid-based cytology (procedure)|Procedure|false|false||lbsnull|Pounds|LabModifier|false|false||lbsnull|liquid-based cytology (procedure)|Procedure|false|false||lbsnull|Pounds|LabModifier|false|false||lbsnull|Desire for food|Finding|false|false||appetitenull|Still|Disorder|false|false||stillnull|Language Ability Proficiency - Good|Finding|false|false||good
null|Language Proficiency - Good|Finding|false|false||goodnull|Specimen Quality - Good|Modifier|false|false||good
null|Good|Modifier|false|false||goodnull|Smaller|Modifier|false|false||lessnull|Less Than|LabModifier|false|false||lessnull|Hunger|Finding|false|false||hungrynull|Daughter|Subject|false|false||Daughternull|Marked|Modifier|false|false||marked
null|Massive|Modifier|false|false||markednull|Memory observations|Finding|false|false||memory
null|Memory G-code|Finding|false|false||memory
null|Memory|Finding|false|false||memorynull|Memory Device|Device|false|false||memorynull|week|Time|false|false||weeksnull|year|Time|false|false||yearsnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Dinner|Finding|false|false||dinnernull|With dinner|Time|false|false||dinnernull|week|Time|false|false||weeksnull|Entity Name Part Type - family|Finding|false|false||family
null|Last Name|Finding|false|false||family
null|Living Arrangement - Family|Finding|false|false||family
null|Family (taxonomic)|Finding|false|false||family
null|Family Collection|Finding|false|false||familynull|Family|Subject|false|false||familynull|Visit|Finding|false|false||visitnull|MELTF-AS1 gene|Finding|false|false||planenull|Airplanes|Device|false|false||planenull|Anatomic Plane|Modifier|false|false||planenull|Pillow|Device|false|false||pillownull|sleeping upright or using specific number of extra pillows (orthopnea)|Finding|false|false||orthopnea
null|Orthopnea|Finding|false|false||orthopneanull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Atrial Fibrillation|Disorder|false|false||Atrial fibrillationnull|null|Attribute|false|false||Atrial fibrillationnull|Atrial Fibrillation by ECG Finding|Lab|false|false||Atrial fibrillationnull|Heart Atrium|Anatomy|false|false||Atrialnull|Fibrillation|Disorder|false|false||fibrillationnull|Eliquis|Drug|false|false||Eliquis
null|Eliquis|Drug|false|false||Eliquisnull|Congestive heart failure|Disorder|false|false||CHFnull|Choroidal fissure|Anatomy|false|false||CHFnull|Hypercholesterolemia|Disorder|false|false||Hypercholesterolemianull|Hypercholesterolemia result|Finding|false|false||Hypercholesterolemianull|Hypertensive disease|Disorder|false|false||Hypertensionnull|Social and personal history|Finding|false|false||Social History
null|Social History|Finding|false|false||Social Historynull|Social|Finding|false|false||Socialnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Family Medical History|Finding|false|false||Family Historynull|Entity Name Part Type - family|Finding|false|false||Family
null|Last Name|Finding|false|false||Family
null|Living Arrangement - Family|Finding|false|false||Family
null|Family (taxonomic)|Finding|false|false||Family
null|Family Collection|Finding|false|false||Familynull|Family|Subject|false|false||Familynull|History of present illness (finding)|Finding|false|true||History
null|History of previous events|Finding|false|true||History
null|Historical aspects qualifier|Finding|false|true||History
null|Medical History|Finding|false|true||History
null|Concept History|Finding|false|true||Historynull|History|Subject|false|false||Historynull|Indirect exposure mechanism - Father|Finding|false|false||Father
null|Relationship - Father|Finding|false|false||Father
null|Father - courtesy title|Finding|false|false||Fathernull|Father (person)|Subject|false|false||Fathernull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Alcoholics|Subject|false|false||alcoholicnull|Schizophrenia|Disorder|false|false||schizophrenianull|Relationship - Mother|Finding|false|false||Mothernull|Mother (person)|Subject|false|false||Mothernull|Congestive heart failure|Disorder|false|false||CHFnull|Choroidal fissure|Anatomy|false|false||CHFnull|Brother - courtesy title|Finding|false|false||Brother
null|Relationship - Brother|Finding|false|false||Brothernull|Brothers|Subject|false|false||Brothernull|Cerebrovascular accident|Disorder|false|false||strokenull|Stroke (heart beat)|Finding|false|false||strokenull|Carotid Stenosis|Disorder|false|false||carotid stenosisnull|Carotid Arteries|Anatomy|false|false||carotidnull|Stenosis|Finding|false|false||stenosisnull|Stenosis <Pimeliinae>|Entity|false|false||stenosisnull|Stenosis Morphology|Modifier|false|false||stenosisnull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Generalnull|General medical service|Procedure|false|false||Generalnull|Generalized|Modifier|false|false||Generalnull|Awake (finding)|Finding|false|false||Awakenull|Awakening (time frame)|Time|false|false||Awakenull|cooperative|Entity|false|false||cooperativenull|Elderly woman|Subject|false|false||elderly womannull|Elderly (population group)|Subject|false|false||elderlynull|Old age|Time|false|false||elderlynull|Woman|Subject|false|false||woman
null|Human, Female adult|Subject|false|false||womannull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|HEENT|Anatomy|false|false||HEENTnull|Scleral icterus|Finding|true|false||scleral icterusnull|Sclera|Anatomy|false|false||scleralnull|Icterus|Finding|true|false||icterusnull|Icterus <Icteridae>|Entity|true|false||icterusnull|null|LabModifier|false|false||icterusnull|Myelofibrosis|Disorder|false|false||MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false||MMMnull|Lesion|Finding|true|false||lesionsnull|Oropharyngeal|Anatomy|false|false||oropharynxnull|Passive joint movement of neck (finding)|Finding|false|false||Neck
null|Neck problem|Finding|false|false||Necknull|dendritic spine neck|Anatomy|false|false||Neck
null|Neck|Anatomy|false|false||Necknull|Supple|Finding|false|false||Supplenull|Nuchal Rigidity|Finding|true|false||nuchal rigiditynull|nuchal|Modifier|false|false||nuchalnull|Muscle Rigidity|Finding|true|false||rigiditynull|plastic property - rigidity|Phenomenon|true|false||rigiditynull|Pulmonary (intended site)|Finding|false|false||Pulmonarynull|Lung|Anatomy|false|false||Pulmonarynull|null|Attribute|false|false||Pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||Pulmonarynull|Work of Breathing|Finding|false|false||work of breathingnull|Work|Event|false|false||worknull|outcomes otolaryngology breathing|Finding|false|false||breathing
null|Inspiration (function)|Finding|false|false||breathing
null|Respiration|Finding|false|false||breathingnull|null|Attribute|false|false||breathingnull|respiratory system process|Phenomenon|false|false||breathingnull|Cardiac attachment|Finding|false|false||Cardiacnull|Heart|Anatomy|false|false||Cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||Cardiacnull|Feels warm|Finding|false|false||warmnull|warming process|Phenomenon|false|false||warmnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Malignant neoplasm of abdomen|Disorder|false|false||Abdomennull|Abdomen problem|Finding|false|false||Abdomennull|Abdomen|Anatomy|false|false||Abdomen
null|Abdominal Cavity|Anatomy|false|false||Abdomennull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|All extremities|Anatomy|false|false||Extremities
null|Limb structure|Anatomy|false|false||Extremitiesnull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||Skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false||Skinnull|Skin Specimen Source Code|Finding|false|false||Skin
null|Skin Specimen|Finding|false|false||Skinnull|Skin, Human|Anatomy|false|false||Skin
null|Skin|Anatomy|false|false||Skinnull|Ecchymosis|Finding|false|false||ecchymosesnull|Shin|Anatomy|false|false||shinnull|More|LabModifier|false|false||morenull|Extensive|Modifier|false|false||extensivenull|Shin|Anatomy|false|false||shinnull|Neurologic (qualifier value)|Modifier|false|false||Neurologicnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Able (qualifier value)|Finding|false|false||Ablenull|Ability|Subject|false|false||Ablenull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|MDF Attribute Type - Name|Finding|false|false||name
null|Person Name|Finding|false|false||name
null|Name|Finding|false|false||namenull|Name (property) (qualifier value)|Modifier|false|false||namenull|Backward (qualifier value)|Modifier|false|false||backward
null|Retrograde direction|Modifier|false|false||backwardnull|Programming Languages|Finding|true|false||Languagenull|null|Attribute|true|false||Languagenull|Languages|Entity|true|false||Languagenull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|speech fluency repetition (physical finding)|Finding|false|false||repetition
null|Repeat|Finding|false|false||repetitionnull|Comprehension|Finding|false|false||comprehensionnull|Prosody|Finding|false|false||prosodynull|error|Modifier|false|false||errorsnull|Able (qualifier value)|Finding|false|false||Ablenull|Ability|Subject|false|false||Ablenull|MDF Attribute Type - Name|Finding|false|false||name
null|Person Name|Finding|false|false||name
null|Name|Finding|false|false||namenull|Name (property) (qualifier value)|Modifier|false|false||namenull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Low frequency (qualifier value)|Time|false|false||low frequencynull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Frequency|Finding|false|false||frequency
null|How Often|Finding|false|false||frequencynull|With frequency|Time|false|false||frequency
null|Frequencies (time pattern)|Time|false|false||frequencynull|Kind of quantity - Frequency|LabModifier|false|false||frequency
null|Statistical Frequency|LabModifier|false|false||frequency
null|Spatial Frequency|LabModifier|false|false||frequencynull|Physical object|Entity|false|false||objectsnull|Able (qualifier value)|Finding|false|false||Ablenull|Ability|Subject|false|false||Ablenull|Has difficulty doing (qualifier value)|Finding|false|false||difficultynull|Dysarthria|Disorder|true|false||dysarthrianull|Able (qualifier value)|Finding|false|false||Ablenull|Ability|Subject|false|false||Ablenull|midline cell component|Anatomy|false|false||midlinenull|Midline (qualifier value)|Modifier|false|false||midlinenull|Evidence of (contextual qualifier)|Finding|false|false||evidence ofnull|Evidence|Finding|false|false||evidencenull|Apraxias|Disorder|true|false||apraxianull|Victim of neglect (finding)|Finding|false|false||neglectnull|Neglect (event)|Event|false|false||neglectnull|Neoplasm of uncertain or unknown behavior of cranial nerves|Disorder|false|false||Cranial Nerves
null|Benign neoplasm of cranial nerves|Disorder|false|false||Cranial Nervesnull|Cranial Nerves|Anatomy|false|false||Cranial Nervesnull|Bone structure of cranium|Anatomy|false|false||Cranialnull|Cranial|Modifier|false|false||Cranialnull|Nerve|Anatomy|false|false||Nervesnull|Pupil equal round and reacting to light|Finding|false|false||PERRLnull|Brisk|Modifier|false|false||brisknull|Nystagmus|Disorder|false|false||nystagmusnull|Saccades|Finding|false|false||saccadesnull|Social confrontation skill|Finding|false|false||confrontationnull|Confrontation visual field test|Procedure|false|false||confrontation
null|Confrontation|Procedure|false|false||confrontationnull|facial sensation|Finding|false|false||Facial sensationnull|Face|Anatomy|false|false||Facialnull|Facial|Modifier|false|false||Facialnull|Observation of Sensation|Finding|false|false||sensation
null|Sensory perception|Finding|false|false||sensationnull|sensory exam|Procedure|false|false||sensationnull|Sensation quality|Modifier|false|false||sensationnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Light touch|Finding|false|false||light touchnull|TNFSF14 protein, human|Drug|false|false||light
null|TNFSF14 protein, human|Drug|false|false||lightnull|Light - subjective measurement|Finding|false|false||light
null|TNFSF14 wt Allele|Finding|false|false||light
null|TNFSF14 gene|Finding|false|false||light
null|Light color|Finding|false|false||lightnull|Phototherapy|Procedure|false|false||lightnull|Light|Phenomenon|false|false||lightnull|Light (qualifier)|Modifier|false|false||lightnull|Touch sensation|Finding|false|false||touch
null|Touch Perception|Finding|false|false||touchnull|Therapeutic Touch|Procedure|false|false||touchnull|Tactile|Modifier|false|false||touchnull|Roman numeral VII|Finding|false|false||VIInull|Lamina VII of gray matter of spinal cord|Anatomy|false|false||VII
null|lobule VII|Anatomy|false|false||VII
null|layer VII (Cajal)|Anatomy|false|false||VIInull|Facial Paresis|Disorder|true|false||facial droopnull|Unilateral facial palsy|Finding|true|false||facial droopnull|Face|Anatomy|false|false||facialnull|Facial|Modifier|false|false||facialnull|Face|Anatomy|false|false||facialnull|Facial|Modifier|false|false||facialnull|Set of muscles|Anatomy|false|false||musculaturenull|Symmetric Relationship|Finding|false|false||symmetric
null|Symmetrical|Finding|false|false||symmetricnull|Roman numeral VIII|Finding|false|false||VIII
null|COX8A gene|Finding|false|false||VIIInull|Lamina VIII of gray matter of spinal cord|Anatomy|false|false||VIII
null|Cerebellar pyramis|Anatomy|false|false||VIIInull|outcomes otolaryngology hearing|Finding|false|false||Hearing
null|Hearing finding|Finding|false|false||Hearing
null|Hearing|Finding|false|false||Hearingnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Upper extremity>Finger|Anatomy|false|false||finger
null|Fingers|Anatomy|false|false||finger
null|Fingers not including thumb|Anatomy|false|false||fingernull|Snap brand of resin|Drug|false|false||snappingnull|Hearing Aids|Device|false|false||hearing aidsnull|outcomes otolaryngology hearing|Finding|false|false||hearing
null|Hearing finding|Finding|false|false||hearing
null|Hearing|Finding|false|false||hearingnull|Acquired Immunodeficiency Syndrome|Disorder|false|false||aidsnull|Palate|Anatomy|false|false||Palatenull|Strength (attribute)|Finding|false|false||strengthnull|Pharmaceutical Strength|LabModifier|false|false||strength
null|Physical Strength|LabModifier|false|false||strengthnull|Benign neoplasm of tongue|Disorder|false|false||Tonguenull|Procedure on tongue|Procedure|false|false||Tonguenull|Tongue|Anatomy|false|false||Tonguenull|midline cell component|Anatomy|false|false||midlinenull|Midline (qualifier value)|Modifier|false|false||midlinenull|Language Ability Proficiency - Good|Finding|false|false||good
null|Language Proficiency - Good|Finding|false|false||goodnull|Specimen Quality - Good|Modifier|false|false||good
null|Good|Modifier|false|false||goodnull|Strength (attribute)|Finding|false|false||Strengthnull|Pharmaceutical Strength|LabModifier|false|false||Strength
null|Physical Strength|LabModifier|false|false||Strengthnull|Full|Modifier|false|false||fullnull|Benign neoplasm of tongue|Disorder|false|false||tonguenull|Procedure on tongue|Procedure|false|false||tonguenull|Tongue|Anatomy|false|false||tonguenull|Cheek structure|Anatomy|false|false||cheeknull|Testing|Finding|false|false||testing
null|Tests (qualifier value)|Finding|false|false||testingnull|motor movement|Finding|false|false||Motornull|Motor Device|Device|false|false||Motornull|Bulk (conceptual)|Drug|false|false||bulk
null|Dietary Fiber|Drug|false|false||bulknull|Pronator drift|Finding|true|false||pronator driftnull|Movement|Finding|false|false||movementsnull|Tremor|Finding|false|false||tremornull|Asterixis|Finding|false|false||asterixisnull|Sensory (qualifier value)|Modifier|false|false||Sensorynull|Deficit|Modifier|false|false||deficitsnull|Light touch|Finding|false|false||light touchnull|TNFSF14 protein, human|Drug|false|false||light
null|TNFSF14 protein, human|Drug|false|false||lightnull|Light - subjective measurement|Finding|false|false||light
null|TNFSF14 wt Allele|Finding|false|false||light
null|TNFSF14 gene|Finding|false|false||light
null|Light color|Finding|false|false||lightnull|Phototherapy|Procedure|false|false||lightnull|Light|Phenomenon|false|false||lightnull|Light (qualifier)|Modifier|false|false||lightnull|Touch Perception|Finding|false|false||touch
null|Touch sensation|Finding|false|false||touchnull|Therapeutic Touch|Procedure|false|false||touchnull|Tactile|Modifier|false|false||touchnull|Body temperature measurement|Procedure|false|false||temperaturenull|Body Temperature|Subject|false|false||temperaturenull|Temperature|LabModifier|false|false||temperaturenull|Decreased vibratory sense|Finding|false|false||Decreased vibratory sensenull|Decreasing|Finding|false|false||Decreased
null|Reduced|Finding|false|false||Decreasednull|Decreased|LabModifier|false|false||Decreasednull|null|Finding|false|false||vibratory sensenull|Sensory perception|Finding|false|false||sensenull|Foot|Anatomy|false|false||feetnull|Foot Unit of Length|LabModifier|false|false||feetnull|Ankle|Anatomy|false|false||anklesnull|Joint position sense|Finding|false|false||Joint position sensenull|Joint problem|Finding|false|false||Jointnull|null|Anatomy|false|false||Joint
null|Joints|Anatomy|false|false||Joint
null|Articular system|Anatomy|false|false||Jointnull|Joint Device|Device|false|false||Jointnull|Position Sense|Finding|false|false||position sensenull|Position of phenotypic abnormality|Modifier|false|false||position
null|Positioning (attribute)|Modifier|false|false||positionnull|Sensory perception|Finding|false|false||sensenull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Hallux structure|Anatomy|false|false||great toesnull|RXFP2 gene|Finding|false|false||greatnull|Greater|LabModifier|false|false||great
null|Large|LabModifier|false|false||greatnull|Lower extremity>Toes|Anatomy|false|false||toes
null|Toes|Anatomy|false|false||toesnull|Extinction, Psychological|Finding|true|false||extinctionnull|DSS brand of docusate sodium|Drug|false|false||DSS
null|DSS brand of docusate sodium|Drug|false|false||DSSnull|DOSAGE-SENSITIVE SEX REVERSAL|Disorder|false|false||DSS
null|Dejerine-Sottas Disease|Disorder|false|false||DSSnull|PMP22 wt Allele|Finding|false|false||DSS
null|NR0B1 gene|Finding|false|false||DSS
null|NR0B1 wt Allele|Finding|false|false||DSS
null|MPZ wt Allele|Finding|false|false||DSSnull|Facial Hemiatrophy|Disorder|false|false||Rombergnull|Absent|Finding|false|false||absentnull|Expression Negative|Lab|false|false||absentnull|Observation of reflex|Finding|false|false||Reflexes
null|Reflex action|Finding|false|false||Reflexesnull|Examination of reflexes|Procedure|false|false||Reflexesnull|imidazole mustard|Drug|false|false||Bic
null|imidazole mustard|Drug|false|false||Bicnull|MIR155HG gene|Finding|false|false||Bic
null|MIR155 gene|Finding|false|false||Bicnull|BIC Regimen|Procedure|false|false||Bicnull|Structure of inferior brachium of corpora quadrigemina|Anatomy|false|false||Bic
null|nucleus of the brachium of the inferior colliculus|Anatomy|false|false||Bicnull|TRI-AAT9-1 gene|Finding|false|false||Tri
null|Temptation and Restraint Inventory|Finding|false|false||Trinull|Fenamole|Drug|false|false||Pat
null|Fenamole|Drug|false|false||Patnull|Paroxysmal atrial tachycardia|Disorder|false|false||Patnull|glutamate-prephenate aminotransferase activity|Finding|false|false||Pat
null|aspartate-prephenate aminotransferase activity|Finding|false|false||Pat
null|protein acetyltransferase activity|Finding|false|false||Patnull|Thermoacoustic Computed Tomography|Procedure|false|false||Patnull|acetylcholine|Drug|false|false||Ach
null|acetylcholine|Drug|false|false||Ach
null|acetylcholine|Drug|false|false||Achnull|Achondroplasia|Disorder|false|false||Achnull|FGFR3 wt Allele|Finding|false|false||Ach
null|FGFR3 gene|Finding|false|false||Ach
null|Ache|Finding|false|false||Achnull|Acoli Language|Entity|false|false||Achnull|Plantar (qualifier value)|Anatomy|false|false||Plantar
null|Sole of Foot|Anatomy|false|false||Plantarnull|Communication Response|Finding|false|false||response
null|Disease Response|Finding|false|false||response
null|Answer (statement)|Finding|false|false||responsenull|Response process|Subject|false|false||responsenull|Flexor (Anatomical coordinate)|Anatomy|false|false||flexornull|Flexor <Diplocrepinae>|Entity|false|false||flexornull|Coordination of Benefits - Coordination|Finding|false|false||Coordination
null|Coordinated|Finding|false|false||Coordination
null|Physiologic Coordination|Finding|false|false||Coordinationnull|Intention tremor|Finding|true|false||intention tremor
null|Action Tremor|Finding|true|false||intention tremornull|null|Finding|false|false||intentionnull|intent|Modifier|false|false||intentionnull|Tremor|Finding|true|false||tremornull|Cerebellar Dysmetria|Finding|true|false||dysmetrianull|fenofibrate|Drug|false|false||FNF
null|fenofibrate|Drug|false|false||FNFnull|Heel|Anatomy|false|false||heelnull|Cerebellar Dysmetria|Finding|true|false||dysmetrianull|Unable|Finding|false|false||Unablenull|Examination of knee joint|Procedure|false|false||kneenull|Knee region structure|Anatomy|false|false||knee
null|Knee|Anatomy|false|false||knee
null|Lower extremity>Knee|Anatomy|false|false||knee
null|Knee joint|Anatomy|false|false||kneenull|Operative procedure on knee|Procedure|false|false||knee surgerynull|Examination of knee joint|Procedure|false|false||kneenull|Knee region structure|Anatomy|false|false||knee
null|Knee|Anatomy|false|false||knee
null|Lower extremity>Knee|Anatomy|false|false||knee
null|Knee joint|Anatomy|false|false||kneenull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Gait|Finding|false|false||Gaitnull|Unable|Finding|false|false||unablenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Walkers|Device|false|false||walkernull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|Data|Finding|false|false||Datanull|Data call receiving device|Device|false|false||Datanull|Data <Amphipyrinae>|Entity|false|false||Datanull|Last|Modifier|false|false||lastnull|C1orf210 gene|Finding|false|false||Tempnull|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Procedure|false|false||Tempnull|Temperature|LabModifier|false|false||Tempnull|delivery (history)|Finding|false|false||delivery
null|Transfer Technique|Finding|false|false||delivery
null|null|Finding|false|false||deliverynull|Obstetric Delivery|Procedure|false|false||deliverynull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Generalnull|General medical service|Procedure|false|false||Generalnull|Generalized|Modifier|false|false||Generalnull|Awake (finding)|Finding|false|false||Awakenull|Awakening (time frame)|Time|false|false||Awakenull|cooperative|Entity|false|false||cooperativenull|Elderly woman|Subject|false|false||elderly womannull|Elderly (population group)|Subject|false|false||elderlynull|Old age|Time|false|false||elderlynull|Woman|Subject|false|false||woman
null|Human, Female adult|Subject|false|false||womannull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|HEENT|Anatomy|false|false||HEENTnull|Scleral icterus|Finding|true|false||scleral icterusnull|Sclera|Anatomy|false|false||scleralnull|Icterus|Finding|true|false||icterusnull|Icterus <Icteridae>|Entity|true|false||icterusnull|null|LabModifier|false|false||icterusnull|Myelofibrosis|Disorder|false|false||MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false||MMMnull|Lesion|Finding|true|false||lesionsnull|Oropharyngeal|Anatomy|false|false||oropharynxnull|Passive joint movement of neck (finding)|Finding|false|false||Neck
null|Neck problem|Finding|false|false||Necknull|dendritic spine neck|Anatomy|false|false||Neck
null|Neck|Anatomy|false|false||Necknull|Supple|Finding|false|false||Supplenull|Nuchal Rigidity|Finding|true|false||nuchal rigiditynull|nuchal|Modifier|false|false||nuchalnull|Muscle Rigidity|Finding|true|false||rigiditynull|plastic property - rigidity|Phenomenon|true|false||rigiditynull|Pulmonary (intended site)|Finding|false|false||Pulmonarynull|Lung|Anatomy|false|false||Pulmonarynull|null|Attribute|false|false||Pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||Pulmonarynull|Work of Breathing|Finding|false|false||work of breathingnull|Work|Event|false|false||worknull|outcomes otolaryngology breathing|Finding|false|false||breathing
null|Inspiration (function)|Finding|false|false||breathing
null|Respiration|Finding|false|false||breathingnull|null|Attribute|false|false||breathingnull|respiratory system process|Phenomenon|false|false||breathingnull|Cardiac attachment|Finding|false|false||Cardiacnull|Heart|Anatomy|false|false||Cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||Cardiacnull|Feels warm|Finding|false|false||warmnull|warming process|Phenomenon|false|false||warmnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Malignant neoplasm of abdomen|Disorder|false|false||Abdomennull|Abdomen problem|Finding|false|false||Abdomennull|Abdomen|Anatomy|false|false||Abdomen
null|Abdominal Cavity|Anatomy|false|false||Abdomennull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|All extremities|Anatomy|false|false||Extremities
null|Limb structure|Anatomy|false|false||Extremitiesnull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||Skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false||Skinnull|Skin Specimen Source Code|Finding|false|false||Skin
null|Skin Specimen|Finding|false|false||Skinnull|Skin, Human|Anatomy|false|false||Skin
null|Skin|Anatomy|false|false||Skinnull|Ecchymosis|Finding|false|false||ecchymosesnull|Shin|Anatomy|false|false||shinnull|More|LabModifier|false|false||morenull|Extensive|Modifier|false|false||extensivenull|Shin|Anatomy|false|false||shinnull|Neurologic (qualifier value)|Modifier|false|false||Neurologicnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Person Info|Finding|false|false||personnull|null|Attribute|false|false||personnull|Persons|Subject|false|false||personnull|Able (qualifier value)|Finding|false|false||Ablenull|Ability|Subject|false|false||Ablenull|Relate - vinyl resin|Drug|false|false||relatenull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Programming Languages|Finding|false|false||Languagenull|null|Attribute|false|false||Languagenull|Languages|Entity|false|false||Languagenull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Comprehension|Finding|false|false||comprehensionnull|Prosody|Finding|false|false||prosodynull|error|Modifier|false|false||errorsnull|Dysarthria|Disorder|true|false||dysarthrianull|Able (qualifier value)|Finding|false|false||Ablenull|Ability|Subject|false|false||Ablenull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|midline cell component|Anatomy|false|false||midlinenull|Midline (qualifier value)|Modifier|false|false||midlinenull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Apraxias|Disorder|false|false||apraxianull|Victim of neglect (finding)|Finding|false|false||neglectnull|Neglect (event)|Event|false|false||neglectnull|Neoplasm of uncertain or unknown behavior of cranial nerves|Disorder|false|false||Cranial Nerves
null|Benign neoplasm of cranial nerves|Disorder|false|false||Cranial Nervesnull|Cranial Nerves|Anatomy|false|false||Cranial Nervesnull|Bone structure of cranium|Anatomy|false|false||Cranialnull|Cranial|Modifier|false|false||Cranialnull|Nerve|Anatomy|false|false||Nervesnull|Pupil equal round and reacting to light|Finding|false|false||PERRLnull|Brisk|Modifier|false|false||brisknull|Nystagmus|Disorder|false|false||nystagmusnull|Saccades|Finding|false|false||saccadesnull|facial sensation|Finding|false|false||Facial sensationnull|Face|Anatomy|false|false||Facialnull|Facial|Modifier|false|false||Facialnull|Observation of Sensation|Finding|false|false||sensation
null|Sensory perception|Finding|false|false||sensationnull|sensory exam|Procedure|false|false||sensationnull|Sensation quality|Modifier|false|false||sensationnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Light touch|Finding|false|false||light touchnull|TNFSF14 protein, human|Drug|false|false||light
null|TNFSF14 protein, human|Drug|false|false||lightnull|Light - subjective measurement|Finding|false|false||light
null|TNFSF14 wt Allele|Finding|false|false||light
null|TNFSF14 gene|Finding|false|false||light
null|Light color|Finding|false|false||lightnull|Phototherapy|Procedure|false|false||lightnull|Light|Phenomenon|false|false||lightnull|Light (qualifier)|Modifier|false|false||lightnull|Touch sensation|Finding|false|false||touch
null|Touch Perception|Finding|false|false||touchnull|Therapeutic Touch|Procedure|false|false||touchnull|Tactile|Modifier|false|false||touchnull|Roman numeral VII|Finding|false|false||VIInull|Lamina VII of gray matter of spinal cord|Anatomy|false|false||VII
null|lobule VII|Anatomy|false|false||VII
null|layer VII (Cajal)|Anatomy|false|false||VIInull|Facial Paresis|Disorder|true|false||facial droopnull|Unilateral facial palsy|Finding|true|false||facial droopnull|Face|Anatomy|false|false||facialnull|Facial|Modifier|false|false||facialnull|Face|Anatomy|false|false||facialnull|Facial|Modifier|false|false||facialnull|Set of muscles|Anatomy|false|false||musculaturenull|Symmetric Relationship|Finding|false|false||symmetric
null|Symmetrical|Finding|false|false||symmetricnull|Roman numeral VIII|Finding|false|false||VIII
null|COX8A gene|Finding|false|false||VIIInull|Lamina VIII of gray matter of spinal cord|Anatomy|false|false||VIII
null|Cerebellar pyramis|Anatomy|false|false||VIIInull|outcomes otolaryngology hearing|Finding|false|false||Hearing
null|Hearing finding|Finding|false|false||Hearing
null|Hearing|Finding|false|false||Hearingnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|conversation|Finding|false|false||conversationnull|Palate|Anatomy|false|false||Palatenull|Strength (attribute)|Finding|false|false||strengthnull|Pharmaceutical Strength|LabModifier|false|false||strength
null|Physical Strength|LabModifier|false|false||strengthnull|Benign neoplasm of tongue|Disorder|false|false||Tonguenull|Procedure on tongue|Procedure|false|false||Tonguenull|Tongue|Anatomy|false|false||Tonguenull|midline cell component|Anatomy|false|false||midlinenull|Midline (qualifier value)|Modifier|false|false||midlinenull|Language Ability Proficiency - Good|Finding|false|false||good
null|Language Proficiency - Good|Finding|false|false||goodnull|Specimen Quality - Good|Modifier|false|false||good
null|Good|Modifier|false|false||goodnull|motor movement|Finding|false|false||Motornull|Motor Device|Device|false|false||Motornull|Bulk (conceptual)|Drug|false|false||bulk
null|Dietary Fiber|Drug|false|false||bulknull|Pronator drift|Finding|true|false||pronator driftnull|Movement|Finding|false|false||movementsnull|Tremor|Finding|false|false||tremornull|Asterixis|Finding|false|false||asterixisnull|Structure of deltoid muscle|Anatomy|false|false||Deltnull|imidazole mustard|Drug|false|false||Bic
null|imidazole mustard|Drug|false|false||Bicnull|MIR155HG gene|Finding|false|false||Bic
null|MIR155 gene|Finding|false|false||Bicnull|BIC Regimen|Procedure|false|false||Bicnull|Structure of inferior brachium of corpora quadrigemina|Anatomy|false|false||Bic
null|nucleus of the brachium of the inferior colliculus|Anatomy|false|false||Bicnull|TRI-AAT9-1 gene|Finding|false|false||Tri
null|Temptation and Restraint Inventory|Finding|false|false||Trinull|LGR5 wt Allele|Finding|false|false||FEx
null|LGR5 gene|Finding|false|false||FExnull|Ham|Drug|false|false||Ham
null|ATF7IP protein, human|Drug|false|false||Ham
null|ATF7IP protein, human|Drug|false|false||Hamnull|Tropical Spastic Paraparesis|Disorder|false|false||Hamnull|altretamine/doxorubicin/melphalan protocol|Procedure|false|false||Hamnull|Gas - SpecimenType|Drug|false|false||Gas
null|Gases|Drug|false|false||Gas
null|Gas Dosage Form|Drug|false|false||Gasnull|Gas - Specimen Source Codes|Finding|false|false||Gas
null|gastrointestinal gas|Finding|false|false||Gas
null|PAGR1 wt Allele|Finding|false|false||Gas
null|GALNS wt Allele|Finding|false|false||Gas
null|GALNS gene|Finding|false|false||Gas
null|GAST wt Allele|Finding|false|false||Gas
null|GAST gene|Finding|false|false||Gas
null|germacrene-A synthase activity|Finding|false|false||Gas
null|PAGR1 gene|Finding|false|false||Gasnull|Examination of knee joint|Procedure|false|false||Kneenull|Knee region structure|Anatomy|false|false||Knee
null|Knee|Anatomy|false|false||Knee
null|Lower extremity>Knee|Anatomy|false|false||Knee
null|Knee joint|Anatomy|false|false||Kneenull|History of surgery|Finding|false|false||prior surgerynull|null|Time|false|false||priornull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Sensory (qualifier value)|Modifier|false|false||Sensorynull|Deficit|Modifier|false|false||deficitsnull|Light touch|Finding|false|false||light touchnull|TNFSF14 protein, human|Drug|false|false||light
null|TNFSF14 protein, human|Drug|false|false||lightnull|Light - subjective measurement|Finding|false|false||light
null|TNFSF14 wt Allele|Finding|false|false||light
null|TNFSF14 gene|Finding|false|false||light
null|Light color|Finding|false|false||lightnull|Phototherapy|Procedure|false|false||lightnull|Light|Phenomenon|false|false||lightnull|Light (qualifier)|Modifier|false|false||lightnull|Touch Perception|Finding|false|false||touch
null|Touch sensation|Finding|false|false||touchnull|Therapeutic Touch|Procedure|false|false||touchnull|Tactile|Modifier|false|false||touchnull|Coordination of Benefits - Coordination|Finding|false|false||Coordination
null|Coordinated|Finding|false|false||Coordination
null|Physiologic Coordination|Finding|false|false||Coordinationnull|Intention tremor|Finding|true|false||intention tremor
null|Action Tremor|Finding|true|false||intention tremornull|null|Finding|false|false||intentionnull|intent|Modifier|false|false||intentionnull|Tremor|Finding|true|false||tremornull|Cerebellar Dysmetria|Finding|true|false||dysmetrianull|fenofibrate|Drug|false|false||FNF
null|fenofibrate|Drug|false|false||FNFnull|Gait|Finding|false|false||Gaitnull|Walkers|Device|false|false||walkernull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Monos|Drug|false|false||Monos
null|Mono-S|Drug|false|false||Monos
null|Monos|Drug|false|false||Monosnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||Eos
null|Familial eosinophilia|Disorder|false|false||Eosnull|PRSS33 gene|Finding|false|false||Eos
null|IKZF4 gene|Finding|false|false||Eosnull|Eos <Loriini>|Entity|false|false||Eosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MB
null|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MBnull|creatine kinase activity|Finding|false|false||CK-MBnull|Serum creatine phosphokinase MB isoenzyme measurement|Procedure|false|false||CK-MB
null|Creatine kinase MB measurement|Procedure|false|false||CK-MBnull|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|High Density Lipoproteins|Drug|false|false||HDL
null|High Density Lipoproteins|Drug|false|false||HDLnull|HSD11B1 wt Allele|Finding|false|false||HDLnull|High density lipoprotein measurement|Procedure|false|false||HDLnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Glycosylated hemoglobin A|Drug|false|false||HbA1c
null|Glycosylated hemoglobin A|Drug|false|false||HbA1cnull|Glucohemoglobin measurement|Procedure|false|false||HbA1cnull|KCNH1 gene|Finding|false|false||eAGnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|thyrotropin|Drug|false|false||TSH
null|thyrotropin|Drug|false|false||TSH
null|thyrotropin|Drug|false|false||TSHnull|Thyroid stimulating hormone measurement|Procedure|false|false||TSHnull|null|Attribute|false|false||TSHnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|AB(S) hearing assessment list|Device|false|false||Abnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Color of urine|Finding|false|false||URINE Colornull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|color additive|Drug|false|false||Color
null|Coloring Excipient|Drug|false|false||Colornull|color - solid dosage form|Modifier|false|false||Color
null|Color|Modifier|false|false||Colornull|Color quantity|LabModifier|false|false||Colornull|Cereal plant straw|Drug|false|false||Strawnull|Straw package type|Device|false|false||Strawnull|Straw Color|Modifier|false|false||Strawnull|Straw (unit of presentation)|LabModifier|false|false||Strawnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Hematuria|Disorder|false|false||URINE Bloodnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Blood and lymphatic system disorders|Disorder|false|false||Bloodnull|peripheral blood|Finding|false|false||Blood
null|Blood|Finding|false|false||Blood
null|In Blood|Finding|false|false||Bloodnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|nitrite ion|Drug|false|false||Nitrite
null|Nitrites|Drug|false|false||Nitrite
null|Nitrites|Drug|false|false||Nitrite
null|Nitrites|Drug|false|false||Nitrite
null|nitrite ion|Drug|false|false||Nitrite
null|nitrite ion|Drug|false|false||Nitritenull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Proteins|Drug|false|false||Protein
null|Proteins|Drug|false|false||Proteinnull|Protein Info|Finding|false|false||Proteinnull|Protein measurement|Procedure|false|false||Proteinnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Ketones|Drug|false|false||Ketonenull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Cancer/Testis Antigen|Drug|false|false||CTAnull|PCYT1A wt Allele|Finding|false|false||CTA
null|CERNA3 gene|Finding|false|false||CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false||CTAnull|Problems with head|Disorder|false|false||headnull|Procedure on head|Procedure|false|false||headnull|Structure of head of caudate nucleus|Anatomy|false|false||head
null|Head|Anatomy|false|false||headnull|Head Device|Device|false|false||headnull|Passive joint movement of neck (finding)|Finding|false|false||neck
null|Neck problem|Finding|false|false||necknull|dendritic spine neck|Anatomy|false|false||neck
null|Neck|Anatomy|false|false||necknull|Opinions|Finding|false|false||opinionnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Segmental|Modifier|false|false||Segmentalnull|Occlusion of left vertebral artery (disorder)|Finding|false|false||left vertebral artery occlusionnull|Structure of left vertebral artery|Anatomy|false|false||left vertebral arterynull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Vertebral artery obstruction (disorder)|Finding|false|false||vertebral artery occlusionnull|Structure of vertebral artery|Anatomy|false|false||vertebral artery
null|Head+Neck>Vertebral artery|Anatomy|false|false||vertebral arterynull|Bone structure of spine|Anatomy|false|false||vertebralnull|Occlusion of artery (disorder)|Finding|false|false||artery occlusionnull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Complete obstruction|Disorder|false|false||occlusionnull|Cardiovascular occlusion|Finding|false|false||occlusion
null|Occluded|Finding|false|false||occlusion
null|Dental Occlusion|Finding|false|false||occlusion
null|Obstruction|Finding|false|false||occlusion
null|null|Finding|false|false||occlusionnull|Indeterminate|Modifier|false|false||indeterminatenull|Chronicity|Time|false|false||chronicitynull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Ischemia|Finding|true|false||ischemianull|Ischemia Procedure|Procedure|true|false||ischemianull|Somewhat|Finding|false|false||Somewhatnull|Small|LabModifier|false|false||smallnull|Diameter (qualifier value)|LabModifier|false|false||calibernull|Attenuation|Event|false|false||attenuatednull|Attenuated by (contextual qualifier)|Modifier|false|false||attenuatednull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|inferiority|Finding|false|false||inferiornull|Inferior|Modifier|false|false||inferiornull|Macromolecular Branch|Drug|false|false||branchnull|Branch of|Modifier|false|false||branchnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Focal|Modifier|false|false||focalnull|Complete obstruction|Disorder|true|false||occlusionnull|Cardiovascular occlusion|Finding|true|false||occlusion
null|Occluded|Finding|true|false||occlusion
null|Dental Occlusion|Finding|true|false||occlusion
null|Obstruction|Finding|true|false||occlusion
null|null|Finding|true|false||occlusionnull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|false|false||acutenull|Intracranial Route of Administration|Finding|false|false||intracranialnull|Intracranial|Anatomy|false|false||intracranialnull|Congenital Abnormality|Disorder|false|false||abnormalitynull|Abnormality|Finding|false|false||abnormalitynull|CAT scan of head|Procedure|false|false||CT headnull|null|Attribute|false|false||CT headnull|Problems with head|Disorder|false|false||headnull|Procedure on head|Procedure|false|false||headnull|Structure of head of caudate nucleus|Anatomy|false|false||head
null|Head|Anatomy|false|false||headnull|Head Device|Device|false|false||headnull|MRI of head|Procedure|false|false||MRI headnull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|Problems with head|Disorder|false|false||headnull|Procedure on head|Procedure|false|false||headnull|Structure of head of caudate nucleus|Anatomy|false|false||head
null|Head|Anatomy|false|false||headnull|Head Device|Device|false|false||headnull|Contrast Media|Drug|false|false||contrastnull|Contrast|Modifier|false|false||contrastnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|false|false||acutenull|Intracranial Route of Administration|Finding|false|false||intracranialnull|Intracranial|Anatomy|false|false||intracranialnull|Congenital Abnormality|Disorder|true|false||abnormalitynull|Abnormality|Finding|true|false||abnormalitynull|LARGE1 wt Allele|Finding|true|false||large
null|LARGE1 gene|Finding|true|false||largenull|Large|LabModifier|false|false||largenull|Territory|Entity|false|false||territory
null|Geographic state|Entity|false|false||territorynull|Infarction|Finding|false|false||infarctionnull|Hemorrhage|Finding|false|false||hemorrhagenull|Scattered|Modifier|false|false||Scatterednull|Focal|Modifier|false|false||foci ofnull|Foci|Finding|false|false||focinull|Focal|Modifier|false|false||focinull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|signal intensity|LabModifier|false|false||signal intensitynull|Signal|Phenomenon|false|false||signalnull|With intensity|Modifier|false|false||intensitynull|Subcortical|Anatomy|false|false||subcorticalnull|Periventricular white matter|Anatomy|false|false||periventricular white matternull|Periventricular|Modifier|false|false||periventricularnull|White matter|Anatomy|false|false||white matternull|White (population group)|Subject|false|false||white
null|Caucasian|Subject|false|false||white
null|Caucasians|Subject|false|false||whitenull|White color|Modifier|false|false||whitenull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Structure of small blood vessel (organ)|Anatomy|false|false||small vesselnull|Small|LabModifier|false|false||smallnull|Vessel Positions|Anatomy|false|false||vessel
null|Blood Vessel|Anatomy|false|false||vesselnull|Vessel (unit of presentation)|LabModifier|false|false||vesselnull|Disease|Disorder|false|false||diseasenull|Transthoracic echocardiography|Procedure|false|false||TTEnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Structure|Modifier|false|false||structuralnull|Source (property) (qualifier value)|Finding|true|false||source
null|Term Source|Finding|true|false||source
null|Source|Finding|true|false||sourcenull|Thromboembolism|Finding|true|false||thromboembolismnull|Rhythm|Finding|false|false||rhythm
null|rhythmic process (biological)|Finding|false|false||rhythmnull|Thrombus formation|Finding|false|false||thrombus formationnull|Thrombus|Finding|false|false||thrombus
null|Blood Clot|Finding|false|false||thrombusnull|Thrombus <Thrombidae>|Entity|false|false||thrombusnull|Formation|Finding|false|false||formationnull|Anabolism|Phenomenon|false|false||formationnull|Formations|Modifier|false|false||formationnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Heart Ventricle|Anatomy|false|false||ventricularnull|Ventricular|Modifier|false|false||ventricularnull|Systole|Finding|false|false||systolicnull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Variability|Finding|false|false||variabilitynull|Cardiac Arrhythmia|Disorder|false|false||arrhythmianull|Mild to moderate|Modifier|false|false||Mild to moderatenull|Mild Severity of Illness Code|Finding|false|false||Mildnull|Mild (qualifier value)|Modifier|false|false||Mild
null|Mild Allergy Severity|Modifier|false|false||Mildnull|Moderate - Severity of Illness Code|Finding|false|false||moderate
null|Moderate|Finding|false|false||moderatenull|Moderate (severity modifier)|Modifier|false|false||moderate
null|Moderate - Allergy Severity|Modifier|false|false||moderate
null|Moderation|Modifier|false|false||moderatenull|mitral|Modifier|false|false||mitralnull|Tricuspid Valve Insufficiency|Disorder|false|false||tricuspid regurgitationnull|Tricuspid|Modifier|false|false||tricuspidnull|Regurgitation|Finding|false|false||regurgitation
null|Regurgitates after swallowing|Finding|false|false||regurgitationnull|Regurgitation - mechanism|Phenomenon|false|false||regurgitationnull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Very|Modifier|false|false||Verynull|Small|LabModifier|false|false||smallnull|Pericardial effusion|Disorder|false|false||pericardial effusionnull|Pericardial effusion body substance|Finding|false|false||pericardial effusionnull|Pericardial (qualifier value)|Anatomy|false|false||pericardial
null|Pericardial sac structure|Anatomy|false|false||pericardialnull|Effusion (substance)|Finding|false|false||effusion
null|null|Finding|false|false||effusion
null|effusion|Finding|false|false||effusionnull|BRIEF Health Literacy Screening Tool|Finding|false|false||Brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||Briefnull|Brief|Time|false|false||Briefnull|Shortened|Modifier|false|false||Briefnull|Hospital course|Finding|false|false||Hospital Coursenull|null|Attribute|false|false||Hospital Coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||Coursenull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Old|Time|false|false||oldnull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|Atrial Fibrillation|Disorder|false|false||AFibnull|Atrial Fibrillation by ECG Finding|Lab|false|false||AFibnull|Eliquis|Drug|false|false||Eliquis
null|Eliquis|Drug|false|false||Eliquisnull|Congestive heart failure|Disorder|false|false||CHFnull|Choroidal fissure|Anatomy|false|false||CHFnull|Hypertensive disease|Disorder|false|false||HTNnull|Sudden onset (contextual qualifier) (qualifier value)|Finding|false|false||sudden onsetnull|Sudden onset (attribute)|Time|false|false||sudden onsetnull|Sudden (qualifier value)|Modifier|false|false||suddennull|Onset of (contextual qualifier)|Modifier|false|false||onsetnull|Age of Onset|LabModifier|false|false||onsetnull|Dysarthria|Disorder|false|false||dysarthrianull|Observation Interpretation - Abnormal|Finding|false|false||abnormal
null|Abnormal|Finding|false|false||abnormalnull|Anorectal Malformations|Disorder|false|false||armnull|AKR1A1 wt Allele|Finding|false|false||arm
null|ARMC9 gene|Finding|false|false||armnull|Protocol Treatment Arm|Procedure|false|false||arm
null|Axillary Reverse Mapping|Procedure|false|false||arm
null|Study Arm|Procedure|false|false||armnull|Upper arm|Anatomy|false|false||arm
null|null|Anatomy|false|false||arm
null|Upper Extremity|Anatomy|false|false||armnull|Movement|Finding|false|false||movementsnull|Poor balance (finding)|Finding|false|false||poor balancenull|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group|Finding|false|false||poor
null|Patient Condition Code - Poor|Finding|false|false||poornull|Poverty|Subject|false|false||poornull|Language Proficiency - Poor|Modifier|false|false||poor
null|Specimen Quality - Poor|Modifier|false|false||poor
null|Poor - grade|Modifier|false|false||poor
null|Poor - qualifier|Modifier|false|false||poornull|Balance (substance)|Drug|false|false||balance
null|Balance (substance)|Drug|false|false||balancenull|Ability to balance|Finding|false|false||balance
null|Equilibrium|Finding|false|false||balancenull|examination of balance|Procedure|false|false||balancenull|balance device|Device|false|false||balancenull|Balanced (qualifier value)|Modifier|false|false||balancenull|Walkers|Device|false|false||walkernull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|NIH stroke scale|Finding|false|false||NIHSSnull|Speech|Finding|false|false||speechnull|Speech assessment|Procedure|false|false||speechnull|Cancer/Testis Antigen|Drug|false|false||CTAnull|PCYT1A wt Allele|Finding|false|false||CTA
null|CERNA3 gene|Finding|false|false||CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false||CTAnull|Head and neck structure|Anatomy|false|false||head and necknull|Problems with head|Disorder|false|false||headnull|Procedure on head|Procedure|false|false||headnull|Structure of head of caudate nucleus|Anatomy|false|false||head
null|Head|Anatomy|false|false||headnull|Head Device|Device|false|false||headnull|Passive joint movement of neck (finding)|Finding|false|false||neck
null|Neck problem|Finding|false|false||necknull|dendritic spine neck|Anatomy|false|false||neck
null|Neck|Anatomy|false|false||necknull|Concern|Finding|false|false||concernnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Macromolecular Branch|Drug|false|false||branchnull|Branch of|Modifier|false|false||branchnull|Attenuation|Event|false|false||attenuationnull|Stenosis|Finding|false|false||stenosisnull|Stenosis <Pimeliinae>|Entity|false|false||stenosisnull|Stenosis Morphology|Modifier|false|false||stenosisnull|Complete obstruction|Disorder|false|false||occlusionnull|Cardiovascular occlusion|Finding|false|false||occlusion
null|Occluded|Finding|false|false||occlusion
null|Dental Occlusion|Finding|false|false||occlusion
null|Obstruction|Finding|false|false||occlusion
null|null|Finding|false|false||occlusionnull|Consideration|Finding|false|false||considerationnull|Thrombectomy|Procedure|false|false||thrombectomynull|NIH stroke scale|Finding|false|false||NIHSSnull|arrival - ActRelationshipType|Finding|false|false||arrivalnull|null|Event|false|false||arrivalnull|Candidate|Finding|false|false||candidatenull|Neurology speciality|Title|false|false||Neurologynull|Stroke service|Entity|false|false||stroke servicenull|Cerebrovascular accident|Disorder|false|false||strokenull|Stroke (heart beat)|Finding|false|false||strokenull|ActInformationPrivacyReason - service|Finding|false|false||servicenull|Software Service|Device|false|false||servicenull|Services|Event|false|false||servicenull|Further|Modifier|false|false||furthernull|Processing type - Evaluation|Finding|false|false||evaluationnull|Evaluation procedure|Procedure|false|false||evaluation
null|Evaluation|Procedure|false|false||evaluationnull|Possible|Finding|false|false||possiblenull|Possible diagnosis|Modifier|false|false||possible
null|Possibly Related to Intervention|Modifier|false|false||possiblenull|Transient Cerebral Ischemia|Disorder|false|false||TIA
null|Transient Ischemic Attack|Disorder|false|false||TIAnull|Tacca leontopetaloides|Entity|false|false||TIAnull|Cerebrovascular accident|Disorder|false|false||strokenull|Stroke (heart beat)|Finding|false|false||strokenull|Further|Modifier|false|false||furthernull|Symptoms aspect|Finding|true|false||symptoms
null|Symptoms|Finding|true|false||symptomsnull|During admission|Time|false|false||during admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|MRI of head|Procedure|false|false||MRI headnull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|Problems with head|Disorder|false|false||headnull|Procedure on head|Procedure|false|false||headnull|Structure of head of caudate nucleus|Anatomy|false|false||head
null|Head|Anatomy|false|false||headnull|Head Device|Device|false|false||headnull|Contrast Media|Drug|false|false||contrastnull|Contrast|Modifier|false|false||contrastnull|Evidence of (contextual qualifier)|Finding|false|false||evidence ofnull|Evidence|Finding|false|false||evidencenull|Cerebrovascular accident|Disorder|true|false||strokenull|Stroke (heart beat)|Finding|true|false||strokenull|Report (document)|Finding|false|false||Reportsnull|Reporting|Procedure|false|false||Reportsnull|Recent|Time|false|false||recentnull|Echocardiography|Procedure|false|false||echocardiogramnull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Cardiologists|Subject|false|false||cardiologistnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|findings aspects|Finding|false|false||findingsnull|null|Attribute|false|false||findingsnull|Concern|Finding|false|false||concernnull|Memory observations|Finding|false|false||memory
null|Memory G-code|Finding|false|false||memory
null|Memory|Finding|false|false||memorynull|Memory Device|Device|false|false||memorynull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|Activity of daily living (function)|Finding|false|false||ADLsnull|Meal (occasion for eating)|Finding|false|false||mealsnull|With meals|Time|false|false||mealsnull|ALF protein, human|Drug|false|false||ALF
null|ALF protein, human|Drug|false|false||ALFnull|GTF2A1L wt Allele|Finding|false|false||ALF
null|GTF2A1L gene|Finding|false|false||ALFnull|month|Time|false|false||monthsnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Changing|Finding|true|false||changenull|Change - procedure|Procedure|true|false||changenull|Delta (difference)|LabModifier|false|false||change
null|Changed status|LabModifier|false|false||changenull|Once daily|Time|false|false||once dailynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Daily|Time|false|false||dailynull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Candidate|Finding|false|false||candidatenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|atorvastatin|Drug|false|false||atorvastatin
null|atorvastatin|Drug|false|false||atorvastatinnull|Hyperlipidemia|Disorder|false|false||hyperlipidemia
null|Hyperlipoproteinemias|Disorder|false|false||hyperlipidemianull|Serum lipids high (finding)|Finding|false|false||hyperlipidemianull|Low-Density Lipoproteins|Drug|false|false||LDL
null|Low-Density Lipoproteins|Drug|false|false||LDLnull|Low density lipoprotein cholesterol measurement|Procedure|false|false||LDLnull|Cardiovascular system|Anatomy|false|false||cardiologynull|cardiology (field)|Title|false|false||cardiologynull|Cardiology service|Entity|false|false||cardiologynull|Frequently|Time|false|false||frequentnull|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false||sinus
null|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false||sinusnull|pathologic fistula|Disorder|false|false||sinusnull|Sinus - general anatomical term|Anatomy|false|false||sinus
null|Nasal sinus|Anatomy|false|false||sinusnull|null|Attribute|false|false||pausesnull|Pauses|Time|false|false||pausesnull|Telemetry|Procedure|false|false||telemetrynull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|atenolol|Drug|false|false||atenolol
null|atenolol|Drug|false|false||atenololnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|digoxin|Drug|false|false||digoxin
null|digoxin|Drug|false|false||digoxinnull|Digoxin measurement|Procedure|false|false||digoxinnull|Close|Finding|false|false||close
null|Closed|Finding|false|false||closenull|Cardiovascular system|Anatomy|false|false||cardiologynull|cardiology (field)|Title|false|false||cardiologynull|Cardiology service|Entity|false|false||cardiologynull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Close|Finding|false|false||close
null|Closed|Finding|false|false||closenull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Living Arrangement - Transient|Finding|false|false||Transient
null|Encounter due to vagabond status|Finding|false|false||Transientnull|Transient Population Group|Subject|false|false||Transientnull|Transitory|Time|false|false||Transientnull|Speech|Finding|false|false||speechnull|Speech assessment|Procedure|false|false||speechnull|Instability|Finding|false|false||instabilitynull|Transient Cerebral Ischemia|Disorder|false|false||TIA
null|Transient Ischemic Attack|Disorder|false|false||TIAnull|Tacca leontopetaloides|Entity|false|false||TIAnull|Consultation|Procedure|false|false||consultnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Home visit (procedure)|Procedure|false|false||home servicesnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Clinical Service|Procedure|false|false||servicesnull|Services|Event|false|false||servicesnull|atorvastatin|Drug|false|false||atorvastatin
null|atorvastatin|Drug|false|false||atorvastatinnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|apixaban|Drug|false|false||apixaban
null|apixaban|Drug|false|false||apixabannull|Therapeutic brand of coal tar|Drug|false|false||therapeutic
null|Therapeutic brand of coal tar|Drug|false|false||therapeuticnull|Therapeutic - Location Service Code|Finding|false|false||therapeutic
null|Therapeutic|Finding|false|false||therapeuticnull|Therapeutic procedure|Procedure|false|false||therapeuticnull|Cerebrovascular accident|Disorder|false|false||strokenull|Stroke (heart beat)|Finding|false|false||strokenull|Neurology speciality|Title|false|false||neurologynull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Stroke risk|Finding|false|false||stroke risknull|Cerebrovascular accident|Disorder|false|false||strokenull|Stroke (heart beat)|Finding|false|false||strokenull|risk factors - observation list|Finding|false|false||risk factors
null|risk factors|Finding|false|false||risk factors
null|History of - risk factor|Finding|false|false||risk factorsnull|null|Attribute|false|false||risk factorsnull|Risk|Finding|false|false||risknull|United States Military enlisted E3 (qualifier value)|Finding|false|false||A1cnull|Hemoglobin A1c measurement|Procedure|false|false||A1cnull|Probable diagnosis|Finding|false|false||Likely
null|Probably|Finding|false|false||Likelynull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Segmental|Modifier|false|false||segmentalnull|Occlusion of left vertebral artery (disorder)|Finding|false|false||left vertebral artery occlusionnull|Structure of left vertebral artery|Anatomy|false|false||left vertebral arterynull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Vertebral artery obstruction (disorder)|Finding|false|false||vertebral artery occlusionnull|Structure of vertebral artery|Anatomy|false|false||vertebral artery
null|Head+Neck>Vertebral artery|Anatomy|false|false||vertebral arterynull|Bone structure of spine|Anatomy|false|false||vertebralnull|Occlusion of artery (disorder)|Finding|false|false||artery occlusionnull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Complete obstruction|Disorder|false|false||occlusionnull|Cardiovascular occlusion|Finding|false|false||occlusion
null|Occluded|Finding|false|false||occlusion
null|Dental Occlusion|Finding|false|false||occlusion
null|Obstruction|Finding|false|false||occlusion
null|null|Finding|false|false||occlusionnull|Somewhat|Finding|false|false||somewhatnull|Small|LabModifier|false|false||smallnull|Diameter (qualifier value)|LabModifier|false|false||calibernull|Attenuation|Event|false|false||attenuatednull|Attenuated by (contextual qualifier)|Modifier|false|false||attenuatednull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|inferiority|Finding|false|false||inferiornull|Inferior|Modifier|false|false||inferiornull|Macromolecular Branch|Drug|false|false||branchnull|Branch of|Modifier|false|false||branchnull|Hyperlipidemia|Disorder|false|false||Hyperlipidemia
null|Hyperlipoproteinemias|Disorder|false|false||Hyperlipidemianull|Serum lipids high (finding)|Finding|false|false||Hyperlipidemianull|Low-Density Lipoproteins|Drug|false|false||LDL
null|Low-Density Lipoproteins|Drug|false|false||LDLnull|Low density lipoprotein cholesterol measurement|Procedure|false|false||LDLnull|Obesity|Disorder|false|false||Obesitynull|BODY MASS INDEX QUANTITATIVE TRAIT LOCUS 20|Finding|false|false||Obesitynull|Concern|Finding|true|false||concernnull|Sleep Apnea Syndromes|Disorder|false|false||sleep apneanull|SLEEP APNEA (device)|Device|false|false||sleep apneanull|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleep
null|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleepnull|Sleep|Finding|false|false||sleepnull|Apnea|Finding|false|false||apneanull|Diagnosis Classification - Diagnosis|Finding|false|false||diagnosis
null|diagnosis aspects|Finding|false|false||diagnosisnull|Diagnosis|Procedure|false|false||diagnosisnull|null|Attribute|false|false||diagnosisnull|Echocardiography|Procedure|false|false||echocardiogramnull|Study Object|Finding|false|false||studynull|Scientific Study|Procedure|false|false||study
null|Study|Procedure|false|false||study
null|Clinical Research|Procedure|false|false||studynull|Room of building - Study|Device|false|false||studynull|acetohydroxamic acid|Drug|false|false||AHA
null|acetohydroxamic acid|Drug|false|false||AHAnull|Factor 8 deficiency, acquired|Disorder|false|false||AHA
null|Autoimmune hemolytic anemia|Disorder|false|false||AHAnull|American Hospital Association|Entity|false|false||AHAnull|Arylsulfatase A, human|Drug|false|false||ASA
null|Arylsulfatase A, human|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASAnull|ARSA gene|Finding|false|false||ASAnull|Core Specimen|Finding|false|false||Corenull|viral nucleocapsid location|Anatomy|false|false||Corenull|Processor Core|Device|false|false||Core
null|Core Device|Device|false|false||Corenull|Core|Modifier|false|false||Corenull|Measures (attribute)|Finding|false|false||Measuresnull|Measures|LabModifier|false|false||Measuresnull|Ischemic stroke|Disorder|false|false||Ischemic Strokenull|Ischemic|Finding|false|false||Ischemicnull|Cerebrovascular accident|Disorder|false|false||Strokenull|Stroke (heart beat)|Finding|false|false||Strokenull|Living Arrangement - Transient|Finding|false|false||Transient
null|Encounter due to vagabond status|Finding|false|false||Transientnull|Transient Population Group|Subject|false|false||Transientnull|Transitory|Time|false|false||Transientnull|Ischemic|Finding|false|false||Ischemicnull|Attack (finding)|Finding|false|false||Attack
null|Attack behavior|Finding|false|false||Attacknull|Attack device|Device|false|false||Attacknull|Screening for dysphagia|Procedure|false|false||Dysphagia screeningnull|Deglutition Disorders|Disorder|false|false||Dysphagianull|Screening - procedure intent|Finding|false|false||screening
null|Special screening finding|Finding|false|false||screening
null|Aspects of disease screening|Finding|false|false||screeningnull|research subject screening|Procedure|false|false||screening
null|Disease Screening|Procedure|false|false||screening
null|Screening|Procedure|false|false||screening
null|Screening for cancer|Procedure|false|false||screening
null|Screening procedure|Procedure|false|false||screeningnull|Intake|Finding|false|false||intakenull|Measurement of fluid intake|Procedure|false|false||intake
null|Intake (treatment)|Procedure|false|false||intakenull|Yes - Expanded yes/no indicator|Finding|false|false||Yes
null|Yes (qualifier value)|Finding|false|false||Yes
null|Yes - Identity May Be Divulged|Finding|false|false||Yes
null|Yes (indicator)|Finding|false|false||Yes
null|Yes|Finding|false|false||Yes
null|Yes - Yes/no indicator|Finding|false|false||Yes
null|Yes - Event Expected|Finding|false|false||Yes
null|Yes - Assignment of Benefits|Finding|false|false||Yes
null|YES1 wt Allele|Finding|false|false||Yes
null|YES1 gene|Finding|false|false||Yes
null|Yes - Release Information|Finding|false|false||Yes
null|YES Portal|Finding|false|false||Yes
null|Yes - Notify Clergy Code|Finding|false|false||Yesnull|Yes - Event Seriousness|Modifier|false|false||Yesnull|DVT prophylaxis|Procedure|false|false||DVT Prophylaxisnull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|Prophylactic treatment|Procedure|false|false||Prophylaxisnull|prevention & control|Modifier|false|false||Prophylaxisnull|Yes - Expanded yes/no indicator|Finding|false|false||Yes
null|Yes (qualifier value)|Finding|false|false||Yes
null|Yes - Identity May Be Divulged|Finding|false|false||Yes
null|Yes (indicator)|Finding|false|false||Yes
null|Yes|Finding|false|false||Yes
null|Yes - Yes/no indicator|Finding|false|false||Yes
null|Yes - Event Expected|Finding|false|false||Yes
null|Yes - Assignment of Benefits|Finding|false|false||Yes
null|YES1 wt Allele|Finding|false|false||Yes
null|YES1 gene|Finding|false|false||Yes
null|Yes - Release Information|Finding|false|false||Yes
null|YES Portal|Finding|false|false||Yes
null|Yes - Notify Clergy Code|Finding|false|false||Yesnull|Yes - Event Seriousness|Modifier|false|false||Yesnull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|Endoglin, human|Drug|false|false||end
null|Endoglin, human|Drug|false|false||endnull|end - ActRelationshipCheckpoint|Finding|false|false||end
null|ENG gene|Finding|false|false||end
null|ENG wt Allele|Finding|false|false||endnull|Stop (qualifier value)|Time|false|false||endnull|End|Modifier|false|false||endnull|Day hospital|Device|false|false||hospital daynull|Day hospital|Entity|false|false||hospital daynull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Day 2|Finding|false|false||day 2null|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Yes - Expanded yes/no indicator|Finding|false|false||Yes
null|Yes (qualifier value)|Finding|false|false||Yes
null|Yes - Identity May Be Divulged|Finding|false|false||Yes
null|Yes (indicator)|Finding|false|false||Yes
null|Yes|Finding|false|false||Yes
null|Yes - Yes/no indicator|Finding|false|false||Yes
null|Yes - Event Expected|Finding|false|false||Yes
null|Yes - Assignment of Benefits|Finding|false|false||Yes
null|YES1 wt Allele|Finding|false|false||Yes
null|YES1 gene|Finding|false|false||Yes
null|Yes - Release Information|Finding|false|false||Yes
null|YES Portal|Finding|false|false||Yes
null|Yes - Notify Clergy Code|Finding|false|false||Yesnull|Yes - Event Seriousness|Modifier|false|false||Yesnull|Low-Density Lipoproteins|Drug|false|false||LDL
null|Low-Density Lipoproteins|Drug|false|false||LDLnull|Low density lipoprotein cholesterol measurement|Procedure|false|false||LDLnull|Yes - Expanded yes/no indicator|Finding|false|false||Yes
null|Yes (qualifier value)|Finding|false|false||Yes
null|Yes - Identity May Be Divulged|Finding|false|false||Yes
null|Yes (indicator)|Finding|false|false||Yes
null|Yes|Finding|false|false||Yes
null|Yes - Yes/no indicator|Finding|false|false||Yes
null|Yes - Event Expected|Finding|false|false||Yes
null|Yes - Assignment of Benefits|Finding|false|false||Yes
null|YES1 wt Allele|Finding|false|false||Yes
null|YES1 gene|Finding|false|false||Yes
null|Yes - Release Information|Finding|false|false||Yes
null|YES Portal|Finding|false|false||Yes
null|Yes - Notify Clergy Code|Finding|false|false||Yesnull|Yes - Event Seriousness|Modifier|false|false||Yesnull|Low-Density Lipoproteins|Drug|false|false||LDL
null|Low-Density Lipoproteins|Drug|false|false||LDLnull|Low density lipoprotein cholesterol measurement|Procedure|false|false||LDLnull|Administration of prophylactic statin|Procedure|false|false||statin therapynull|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Drug|false|false||statin
null|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Drug|false|false||statinnull|EEF1A2 gene|Finding|false|false||statinnull|3-hydroxy-3-methylglutaryl-coenzyme A reductase inhibitor (disposition)|Modifier|false|false||statinnull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|simvastatin|Drug|false|false||simvastatin
null|simvastatin|Drug|false|false||simvastatinnull|simvastatin|Drug|false|false||simvastatin
null|simvastatin|Drug|false|false||simvastatinnull|atorvastatin|Drug|false|false||atorvastatin
null|atorvastatin|Drug|false|false||atorvastatinnull|rosuvastatin|Drug|false|false||rosuvastatin
null|rosuvastatin|Drug|false|false||rosuvastatinnull|Low-Density Lipoproteins|Drug|false|false||LDL
null|Low-Density Lipoproteins|Drug|false|false||LDLnull|Low density lipoprotein cholesterol measurement|Procedure|false|false||LDLnull|Yes - Expanded yes/no indicator|Finding|false|false||Yes
null|Yes (qualifier value)|Finding|false|false||Yes
null|Yes - Identity May Be Divulged|Finding|false|false||Yes
null|Yes (indicator)|Finding|false|false||Yes
null|Yes|Finding|false|false||Yes
null|Yes - Yes/no indicator|Finding|false|false||Yes
null|Yes - Event Expected|Finding|false|false||Yes
null|Yes - Assignment of Benefits|Finding|false|false||Yes
null|YES1 wt Allele|Finding|false|false||Yes
null|YES1 gene|Finding|false|false||Yes
null|Yes - Release Information|Finding|false|false||Yes
null|YES Portal|Finding|false|false||Yes
null|Yes - Notify Clergy Code|Finding|false|false||Yesnull|Yes - Event Seriousness|Modifier|false|false||Yesnull|Low-Density Lipoproteins|Drug|false|false||LDL
null|Low-Density Lipoproteins|Drug|false|false||LDLnull|Low density lipoprotein cholesterol measurement|Procedure|false|false||LDLnull|Low-Density Lipoproteins|Drug|false|false||LDL
null|Low-Density Lipoproteins|Drug|false|false||LDLnull|Low density lipoprotein cholesterol measurement|Procedure|false|false||LDLnull|Indication of (contextual qualifier)|Finding|false|false||reasonnull|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Drug|false|false||Statin
null|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Drug|false|false||Statinnull|EEF1A2 gene|Finding|false|false||Statinnull|3-hydroxy-3-methylglutaryl-coenzyme A reductase inhibitor (disposition)|Modifier|false|false||Statinnull|Drug Allergy|Finding|false|false||medication allergynull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Allergy - Charge Type Reason|Finding|false|false||allergy
null|Allergic disposition|Finding|false|false||allergy
null|Hypersensitivity|Finding|false|false||allergy
null|Response to antigens|Finding|false|false||allergy
null|History of allergies|Finding|false|false||allergy
null|Allergic Reaction|Finding|false|false||allergynull|Allergy Specialty|Title|false|false||allergynull|Indication of (contextual qualifier)|Finding|false|false||reasonsnull|null|Attribute|false|false||physiciannull|Physicians|Subject|false|false||physiciannull|Advanced phase|Modifier|false|false||advancednull|HL7PublishingSubSection - practice|Finding|false|false||practice
null|Experience (Practice)|Finding|false|false||practicenull|Nurses|Subject|false|false||nursenull|null|Attribute|false|false||physiciannull|Physicians|Subject|false|false||physiciannull|null|Attribute|false|false||physiciannull|Physicians|Subject|false|false||physiciannull|ANPEP wt Allele|Finding|false|false||APNnull|Advanced Practice Nurse|Subject|false|false||APNnull|Primary Observer's Qualification - Pharmacist|Finding|false|false||pharmacistnull|Pharmacist|Subject|false|false||pharmacistnull|Low-Density Lipoproteins|Drug|false|false||LDL
null|Low-Density Lipoproteins|Drug|false|false||LDLnull|Low density lipoprotein cholesterol measurement|Procedure|false|false||LDLnull|Less Than|LabModifier|false|false||less thannull|Smaller|Modifier|false|false||lessnull|Less Than|LabModifier|false|false||lessnull|mg/dL|LabModifier|false|false||mg/dLnull|Per Deciliter|LabModifier|false|false||/dLnull|Cessation of smoking|Finding|false|false||Smoking cessationnull|Smoking cessation therapy|Procedure|false|false||Smoking cessationnull|Location characteristic ID - Smoking|Finding|false|false||Smoking
null|Smoking|Finding|false|false||Smoking
null|Tobacco smoking behavior|Finding|false|false||Smokingnull|Cessation|Event|false|false||cessationnull|Encounter due to counseling|Finding|false|false||counseling
null|duration of counseling|Finding|false|false||counselingnull|Counseling|Procedure|false|false||counseling
null|Counselling service|Procedure|false|false||counselingnull|Yes - Expanded yes/no indicator|Finding|false|false||Yes
null|Yes (qualifier value)|Finding|false|false||Yes
null|Yes - Identity May Be Divulged|Finding|false|false||Yes
null|Yes (indicator)|Finding|false|false||Yes
null|Yes|Finding|false|false||Yes
null|Yes - Yes/no indicator|Finding|false|false||Yes
null|Yes - Event Expected|Finding|false|false||Yes
null|Yes - Assignment of Benefits|Finding|false|false||Yes
null|YES1 wt Allele|Finding|false|false||Yes
null|YES1 gene|Finding|false|false||Yes
null|Yes - Release Information|Finding|false|false||Yes
null|YES Portal|Finding|false|false||Yes
null|Yes - Notify Clergy Code|Finding|false|false||Yesnull|Yes - Event Seriousness|Modifier|false|false||Yesnull|Indication of (contextual qualifier)|Finding|true|false||reasonnull|Unable|Finding|false|false||unablenull|Education about stroke|Procedure|false|false||Stroke educationnull|Cerebrovascular accident|Disorder|false|false||Strokenull|Stroke (heart beat)|Finding|false|false||Strokenull|Details of education|Finding|false|false||education
null|Educational aspects|Finding|false|false||education
null|Educational Status|Finding|false|false||educationnull|Education (procedure)|Procedure|false|false||education
null|Knowledge acquisition|Procedure|false|false||educationnull|Specialty Type - Education|Title|false|false||educationnull|Personal Attribute|Subject|false|false||personalnull|risk factors - observation list|Finding|false|false||risk factors
null|risk factors|Finding|false|false||risk factors
null|History of - risk factor|Finding|false|false||risk factorsnull|null|Attribute|false|false||risk factorsnull|Risk|Finding|false|false||risknull|activate biological process|Finding|false|false||activate
null|activate - Data Operation|Finding|false|false||activatenull|activation [action]|Event|false|false||activatenull|Ethyl Methanesulfonate|Drug|false|false||EMS
null|Ethyl Methanesulfonate|Drug|false|false||EMS
null|Ethyl Methanesulfonate|Drug|false|false||EMSnull|EMSLR gene|Finding|false|false||EMSnull|Emergency Medical Services|Procedure|false|false||EMSnull|Cerebrovascular accident|Disorder|false|false||strokenull|Stroke (heart beat)|Finding|false|false||strokenull|Cerebrovascular accident|Disorder|false|false||strokenull|Stroke (heart beat)|Finding|false|false||strokenull|warning signs|Event|false|false||warning signsnull|Warning - AcknowledgementDetailType|Finding|false|false||warning
null|Cautionary Warning|Finding|false|false||warning
null|System Alert|Finding|false|false||warning
null|Warning - Error severity|Finding|false|false||warning
null|Warning - EquipmentAlertLevel|Finding|false|false||warningnull|Warning - Alert level|Modifier|false|false||warningnull|Signs and Symptoms|Finding|false|false||signs and symptomsnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Patient need for (contextual qualifier)|Finding|false|false||need fornull|Patient need for (contextual qualifier)|Finding|false|false||neednull|Needs|Modifier|false|false||neednull|follow-up|Procedure|false|false||followupnull|Yes - Expanded yes/no indicator|Finding|false|false||Yes
null|Yes (qualifier value)|Finding|false|false||Yes
null|Yes - Identity May Be Divulged|Finding|false|false||Yes
null|Yes (indicator)|Finding|false|false||Yes
null|Yes|Finding|false|false||Yes
null|Yes - Yes/no indicator|Finding|false|false||Yes
null|Yes - Event Expected|Finding|false|false||Yes
null|Yes - Assignment of Benefits|Finding|false|false||Yes
null|YES1 wt Allele|Finding|false|false||Yes
null|YES1 gene|Finding|false|false||Yes
null|Yes - Release Information|Finding|false|false||Yes
null|YES Portal|Finding|false|false||Yes
null|Yes - Notify Clergy Code|Finding|false|false||Yesnull|Yes - Event Seriousness|Modifier|false|false||Yesnull|Assessment for rehabilitation|Procedure|false|false||Assessment for rehabilitationnull|Knowledge acquisition using a method of assessment|Finding|false|false||Assessmentnull|assessment of cognitive functions|Procedure|false|false||Assessment
null|Physical Examination|Procedure|false|false||Assessment
null|Nutrition Assessment|Procedure|false|false||Assessment
null|null|Procedure|false|false||Assessment
null|null|Procedure|false|false||Assessment
null|null|Procedure|false|false||Assessment
null|null|Procedure|false|false||Assessment
null|Personal care assessment|Procedure|false|false||Assessment
null|null|Procedure|false|false||Assessment
null|null|Procedure|false|false||Assessment
null|null|Procedure|false|false||Assessment
null|Evaluation procedure|Procedure|false|false||Assessment
null|Evaluation|Procedure|false|false||Assessment
null|null|Procedure|false|false||Assessment
null|null|Procedure|false|false||Assessment
null|null|Procedure|false|false||Assessment
null|null|Procedure|false|false||Assessment
null|null|Procedure|false|false||Assessmentnull|Assessed|Event|false|false||Assessmentnull|Encounter due to care involving use of rehabilitation procedures|Finding|false|false||rehabilitation
null|Rehabilitation aspects|Finding|false|false||rehabilitationnull|Rehabilitation therapy|Procedure|false|false||rehabilitationnull|null|Title|false|false||rehabilitationnull|Rehabilitation therapy|Procedure|false|false||rehabnull|Clinical Service|Procedure|false|false||servicesnull|Services|Event|false|false||servicesnull|Yes - Expanded yes/no indicator|Finding|false|false||Yes
null|Yes (qualifier value)|Finding|false|false||Yes
null|Yes - Identity May Be Divulged|Finding|false|false||Yes
null|Yes (indicator)|Finding|false|false||Yes
null|Yes|Finding|false|false||Yes
null|Yes - Yes/no indicator|Finding|false|false||Yes
null|Yes - Event Expected|Finding|false|false||Yes
null|Yes - Assignment of Benefits|Finding|false|false||Yes
null|YES1 wt Allele|Finding|false|false||Yes
null|YES1 gene|Finding|false|false||Yes
null|Yes - Release Information|Finding|false|false||Yes
null|YES Portal|Finding|false|false||Yes
null|Yes - Notify Clergy Code|Finding|false|false||Yesnull|Yes - Event Seriousness|Modifier|false|false||Yesnull|Administration of prophylactic statin|Procedure|false|false||statin therapynull|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Drug|false|false||statin
null|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Drug|false|false||statinnull|EEF1A2 gene|Finding|false|false||statinnull|3-hydroxy-3-methylglutaryl-coenzyme A reductase inhibitor (disposition)|Modifier|false|false||statinnull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|Yes - Expanded yes/no indicator|Finding|false|false||Yes
null|Yes (qualifier value)|Finding|false|false||Yes
null|Yes - Identity May Be Divulged|Finding|false|false||Yes
null|Yes (indicator)|Finding|false|false||Yes
null|Yes|Finding|false|false||Yes
null|Yes - Yes/no indicator|Finding|false|false||Yes
null|Yes - Event Expected|Finding|false|false||Yes
null|Yes - Assignment of Benefits|Finding|false|false||Yes
null|YES1 wt Allele|Finding|false|false||Yes
null|YES1 gene|Finding|false|false||Yes
null|Yes - Release Information|Finding|false|false||Yes
null|YES Portal|Finding|false|false||Yes
null|Yes - Notify Clergy Code|Finding|false|false||Yesnull|Yes - Event Seriousness|Modifier|false|false||Yesnull|Low-Density Lipoproteins|Drug|false|false||LDL
null|Low-Density Lipoproteins|Drug|false|false||LDLnull|Low density lipoprotein cholesterol measurement|Procedure|false|false||LDLnull|Indication of (contextual qualifier)|Finding|false|false||reasonnull|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Drug|false|false||Statin
null|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Drug|false|false||Statinnull|EEF1A2 gene|Finding|false|false||Statinnull|3-hydroxy-3-methylglutaryl-coenzyme A reductase inhibitor (disposition)|Modifier|false|false||Statinnull|Drug Allergy|Finding|false|false||medication allergynull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Allergy - Charge Type Reason|Finding|false|false||allergy
null|Allergic disposition|Finding|false|false||allergy
null|Hypersensitivity|Finding|false|false||allergy
null|Response to antigens|Finding|false|false||allergy
null|History of allergies|Finding|false|false||allergy
null|Allergic Reaction|Finding|false|false||allergynull|Allergy Specialty|Title|false|false||allergynull|Indication of (contextual qualifier)|Finding|false|false||reasonsnull|null|Attribute|false|false||physiciannull|Physicians|Subject|false|false||physiciannull|Advanced phase|Modifier|false|false||advancednull|HL7PublishingSubSection - practice|Finding|false|false||practice
null|Experience (Practice)|Finding|false|false||practicenull|Nurses|Subject|false|false||nursenull|null|Attribute|false|false||physiciannull|Physicians|Subject|false|false||physiciannull|null|Attribute|false|false||physiciannull|Physicians|Subject|false|false||physiciannull|ANPEP wt Allele|Finding|false|false||APNnull|Advanced Practice Nurse|Subject|false|false||APNnull|Primary Observer's Qualification - Pharmacist|Finding|false|false||pharmacistnull|Pharmacist|Subject|false|false||pharmacistnull|Low-Density Lipoproteins|Drug|false|false||LDL
null|Low-Density Lipoproteins|Drug|false|false||LDLnull|Low density lipoprotein cholesterol measurement|Procedure|false|false||LDLnull|Less Than|LabModifier|false|false||less thannull|Smaller|Modifier|false|false||lessnull|Less Than|LabModifier|false|false||lessnull|mg/dL|LabModifier|false|false||mg/dLnull|Per Deciliter|LabModifier|false|false||/dLnull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|Yes - Expanded yes/no indicator|Finding|false|false||Yes
null|Yes (qualifier value)|Finding|false|false||Yes
null|Yes - Identity May Be Divulged|Finding|false|false||Yes
null|Yes (indicator)|Finding|false|false||Yes
null|Yes|Finding|false|false||Yes
null|Yes - Yes/no indicator|Finding|false|false||Yes
null|Yes - Event Expected|Finding|false|false||Yes
null|Yes - Assignment of Benefits|Finding|false|false||Yes
null|YES1 wt Allele|Finding|false|false||Yes
null|YES1 gene|Finding|false|false||Yes
null|Yes - Release Information|Finding|false|false||Yes
null|YES Portal|Finding|false|false||Yes
null|Yes - Notify Clergy Code|Finding|false|false||Yesnull|Yes - Event Seriousness|Modifier|false|false||Yesnull|Type - ParameterizedDataType|Finding|false|false||Type
null|SGCG gene|Finding|false|false||Typenull|null|Modifier|false|false||Typenull|Antiplatelet|Drug|false|false||Antiplateletnull|ANTICOAGULATION (finding)|Finding|false|false||Anticoagulation
null|Anticoagulation function|Finding|false|false||Anticoagulation
null|Decreased Coagulation Activity [PE]|Finding|false|false||Anticoagulationnull|Anticoagulation Therapy|Procedure|false|false||Anticoagulationnull|Oral Dosage Form|Drug|false|false||oralnull|Oral Route of Administration|Finding|false|false||oral
null|Oral (intended site)|Finding|false|false||oralnull|Oral cavity|Anatomy|false|false||oralnull|Oral|Modifier|false|false||oralnull|ANTICOAGULATION (finding)|Finding|false|false||anticoagulation
null|Anticoagulation function|Finding|false|false||anticoagulation
null|Decreased Coagulation Activity [PE]|Finding|false|false||anticoagulationnull|Anticoagulation Therapy|Procedure|false|false||anticoagulationnull|Patients|Subject|false|false||patientsnull|Heart Atrium|Anatomy|false|false||atrialnull|Fibrillation|Disorder|false|false||fibrillationnull|Cardiac Flutter|Finding|false|false||flutternull|Flutter (respiratory device)|Device|false|false||flutternull|Yes - Expanded yes/no indicator|Finding|false|false||Yes
null|Yes (qualifier value)|Finding|false|false||Yes
null|Yes - Identity May Be Divulged|Finding|false|false||Yes
null|Yes (indicator)|Finding|false|false||Yes
null|Yes|Finding|false|false||Yes
null|Yes - Yes/no indicator|Finding|false|false||Yes
null|Yes - Event Expected|Finding|false|false||Yes
null|Yes - Assignment of Benefits|Finding|false|false||Yes
null|YES1 wt Allele|Finding|false|false||Yes
null|YES1 gene|Finding|false|false||Yes
null|Yes - Release Information|Finding|false|false||Yes
null|YES Portal|Finding|false|false||Yes
null|Yes - Notify Clergy Code|Finding|false|false||Yesnull|Yes - Event Seriousness|Modifier|false|false||Yesnull|Cognitive|Finding|false|false||Cognitivenull|Complaint (finding)|Finding|false|false||complaintsnull|TNFAIP1 wt Allele|Finding|false|false||B12
null|NDUFB3 gene|Finding|false|false||B12
null|TNFAIP1 gene|Finding|false|false||B12null|one time|Finding|false|false||one timenull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Dietary Supplementation|Procedure|false|false||supplementationnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Oral Dosage Form|Drug|false|false||oralnull|Oral Route of Administration|Finding|false|false||oral
null|Oral (intended site)|Finding|false|false||oralnull|Oral cavity|Anatomy|false|false||oralnull|Oral|Modifier|false|false||oralnull|TNFAIP1 wt Allele|Finding|false|false||B12
null|NDUFB3 gene|Finding|false|false||B12
null|TNFAIP1 gene|Finding|false|false||B12null|Dietary Supplementation|Procedure|false|false||supplementationnull|treponemal|Finding|false|false||Treponemalnull|Antibody NOS negative|Lab|false|false||antibodies negativenull|antibodies (medication)|Drug|false|false||antibodies
null|antibodies (medication)|Drug|false|false||antibodies
null|Antibodies|Drug|false|false||antibodies
null|Antibodies|Drug|false|false||antibodies
null|Antibodies|Drug|false|false||antibodiesnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|consider|Finding|false|false||considernull|Cognitive|Finding|false|false||cognitivenull|Neurology speciality|Title|false|false||neurologynull|Patient referral|Procedure|false|false||referralnull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Memory observations|Finding|false|false||memory
null|Memory G-code|Finding|false|false||memory
null|Memory|Finding|false|false||memorynull|Memory Device|Device|false|false||memorynull|Has difficulty doing (qualifier value)|Finding|true|false||difficultiesnull|Physical Examination|Procedure|false|false||examination
null|Medical Examination|Procedure|false|false||examinationnull|Examination|Event|false|false||examinationnull|Atrial Fibrillation|Disorder|false|false||Afibnull|Atrial Fibrillation by ECG Finding|Lab|false|false||Afibnull|Frequently|Time|false|false||frequentnull|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false||sinus
null|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false||sinusnull|pathologic fistula|Disorder|false|false||sinusnull|Sinus - general anatomical term|Anatomy|false|false||sinus
null|Nasal sinus|Anatomy|false|false||sinusnull|null|Attribute|false|false||pausesnull|Pauses|Time|false|false||pausesnull|digoxin|Drug|false|false||digoxin
null|digoxin|Drug|false|false||digoxinnull|Digoxin measurement|Procedure|false|false||digoxinnull|Cardiologists|Subject|false|false||cardiologistnull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Appropriate|Modifier|false|false||appropriatenull|Therapeutic brand of coal tar|Drug|false|false||therapeutic
null|Therapeutic brand of coal tar|Drug|false|false||therapeuticnull|Therapeutic - Location Service Code|Finding|false|false||therapeutic
null|Therapeutic|Finding|false|false||therapeuticnull|Therapeutic procedure|Procedure|false|false||therapeuticnull|Eliquis|Drug|false|false||Eliquis
null|Eliquis|Drug|false|false||Eliquisnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|atorvastatin|Drug|false|false||atorvastatin
null|atorvastatin|Drug|false|false||atorvastatinnull|Hypertensive disease|Disorder|false|false||HTNnull|Continuous|Finding|false|false||continuenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Antihypertensive Agents|Drug|false|false||antihypertensivesnull|Troponin|Drug|false|false||troponin
null|Troponin|Drug|false|false||troponinnull|Troponin measurement|Procedure|false|false||troponinnull|physiologic resolution|Finding|false|false||RESOLVED
null|Resolution|Finding|false|false||RESOLVEDnull|Resolved|Modifier|false|false||RESOLVEDnull|Troponin|Drug|false|false||Troponin
null|Troponin|Drug|false|false||Troponinnull|Troponin measurement|Procedure|false|false||Troponinnull|Elevated|Modifier|false|false||elevated
null|High|Modifier|false|false||elevatednull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|On admission|Time|false|false||on admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Raised TSH level|Finding|false|false||elevated TSHnull|thyrotropin|Drug|false|false||TSH
null|thyrotropin|Drug|false|false||TSH
null|thyrotropin|Drug|false|false||TSHnull|Thyroid stimulating hormone measurement|Procedure|false|false||TSHnull|null|Attribute|false|false||TSHnull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Accurate (qualifier value)|Modifier|false|false||accuratenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|atenolol|Drug|false|false||Atenolol
null|atenolol|Drug|false|false||Atenololnull|Daily|Time|false|false||DAILYnull|apixaban|Drug|false|false||Apixaban
null|apixaban|Drug|false|false||Apixabannull|Daily|Time|false|false||DAILYnull|losartan potassium|Drug|false|false||Losartan Potassium
null|losartan potassium|Drug|false|false||Losartan Potassiumnull|losartan|Drug|false|false||Losartan
null|losartan|Drug|false|false||Losartannull|Potassium Drug Class|Drug|false|false||Potassium
null|Dietary Potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassiumnull|Potassium metabolic function|Finding|false|false||Potassiumnull|Potassium measurement|Procedure|false|false||Potassiumnull|Daily|Time|false|false||DAILYnull|digoxin|Drug|false|false||Digoxin
null|digoxin|Drug|false|false||Digoxinnull|Digoxin measurement|Procedure|false|false||Digoxinnull|Daily|Time|false|false||DAILYnull|levofloxacin|Drug|false|false||LevoFLOXacin
null|levofloxacin|Drug|false|false||LevoFLOXacinnull|Every twenty four hours|Time|false|false||Q24Hnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|atorvastatin|Drug|false|false||atorvastatin
null|atorvastatin|Drug|false|false||atorvastatinnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Once daily|Time|false|false||once dailynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Daily|Time|false|false||dailynull|Bedtime (qualifier value)|Time|false|false||bedtime
null|Once a day, at bedtime|Time|false|false||bedtimenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|Cyanocobalamin Drug Class|Drug|false|false||Cyanocobalamin
null|Cyanocobalamin Drug Class|Drug|false|false||Cyanocobalamin
null|vitamin B12|Drug|false|false||Cyanocobalamin
null|vitamin B12|Drug|false|false||Cyanocobalamin
null|vitamin B12|Drug|false|false||Cyanocobalaminnull|microgram|LabModifier|false|false||mcgnull|Daily|Time|false|false||DAILYnull|VITAMIN B12 MEASUREMENT|Procedure|false|false||cyanocobalamin (vitamin B-12)null|Cyanocobalamin Drug Class|Drug|false|false||cyanocobalamin
null|Cyanocobalamin Drug Class|Drug|false|false||cyanocobalamin
null|vitamin B12|Drug|false|false||cyanocobalamin
null|vitamin B12|Drug|false|false||cyanocobalamin
null|vitamin B12|Drug|false|false||cyanocobalaminnull|vitamin B12|Drug|false|false||vitamin B-12
null|cobalamins|Drug|false|false||vitamin B-12
null|cobalamins|Drug|false|false||vitamin B-12
null|vitamin B12|Drug|false|false||vitamin B-12
null|vitamin B12|Drug|false|false||vitamin B-12null|VITAMIN B12 MEASUREMENT|Procedure|false|false||vitamin B-12null|vitamin B complex|Drug|false|false||vitamin B
null|vitamin B complex|Drug|false|false||vitamin B
null|vitamin B complex|Drug|false|false||vitamin B
null|B Vitamin Family|Drug|false|false||vitamin B
null|B Vitamin Family|Drug|false|false||vitamin B
null|VITAMIN B|Drug|false|false||vitamin B
null|VITAMIN B|Drug|false|false||vitamin Bnull|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitaminnull|microgram|LabModifier|false|false||mcgnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Once daily|Time|false|false||once dailynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Daily|Time|false|false||dailynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|apixaban|Drug|false|false||Apixaban
null|apixaban|Drug|false|false||Apixabannull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|atenolol|Drug|false|false||Atenolol
null|atenolol|Drug|false|false||Atenololnull|Daily|Time|false|false||DAILYnull|levofloxacin|Drug|false|false||LevoFLOXacin
null|levofloxacin|Drug|false|false||LevoFLOXacinnull|Every twenty four hours|Time|false|false||Q24Hnull|losartan potassium|Drug|false|false||Losartan Potassium
null|losartan potassium|Drug|false|false||Losartan Potassiumnull|losartan|Drug|false|false||Losartan
null|losartan|Drug|false|false||Losartannull|Potassium Drug Class|Drug|false|false||Potassium
null|Dietary Potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassiumnull|Potassium metabolic function|Finding|false|false||Potassiumnull|Potassium measurement|Procedure|false|false||Potassiumnull|Daily|Time|false|false||DAILYnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Encounter due to vagabond status|Finding|false|false||transient
null|Living Arrangement - Transient|Finding|false|false||transientnull|Transient Population Group|Subject|false|false||transientnull|Transitory|Time|false|false||transientnull|Dysarthria|Disorder|false|false||dysarthrianull|Secondary to|Modifier|false|false||secondary tonull|Neoplasm Metastasis|Disorder|true|false||secondarynull|metastatic qualifier|Finding|true|false||secondarynull|Secondary to|Modifier|false|false||secondarynull|second (number)|LabModifier|false|false||secondarynull|Transient Cerebral Ischemia|Disorder|false|false||TIA
null|Transient Ischemic Attack|Disorder|false|false||TIAnull|Tacca leontopetaloides|Entity|false|false||TIAnull|Cerebrovascular accident|Disorder|false|false||strokenull|Stroke (heart beat)|Finding|false|false||strokenull|Mild Severity of Illness Code|Finding|false|false||Mildnull|Mild (qualifier value)|Modifier|false|false||Mild
null|Mild Allergy Severity|Modifier|false|false||Mildnull|Vitamin B 12 Deficiency|Disorder|false|false||Vitamin B12 deficiencynull|Decreased circulating vitamin B12 concentration|Finding|false|false||Vitamin B12 deficiencynull|Vitamin B12 [EPC]|Drug|false|false||Vitamin B12
null|cobalamins|Drug|false|false||Vitamin B12
null|cobalamins|Drug|false|false||Vitamin B12
null|vitamin B12|Drug|false|false||Vitamin B12
null|vitamin B12|Drug|false|false||Vitamin B12
null|vitamin B12|Drug|false|false||Vitamin B12null|VITAMIN B12 MEASUREMENT|Procedure|false|false||Vitamin B12null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|TNFAIP1 wt Allele|Finding|false|false||B12
null|NDUFB3 gene|Finding|false|false||B12
null|TNFAIP1 gene|Finding|false|false||B12null|Malnutrition|Disorder|false|false||deficiencynull|Deficiency|Finding|false|false||deficiencynull|deficiency aspects|Modifier|false|false||deficiencynull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Disease|Disorder|false|false||Conditionnull|Logical Condition|Finding|false|false||Conditionnull|null|Attribute|false|false||Conditionnull|Condition|Modifier|false|false||Conditionnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Helping Behavior|Finding|false|false||assistancenull|Assisted (qualifier value)|Modifier|false|false||assistancenull|AICDA protein, human|Drug|false|false||aid
null|AICDA protein, human|Drug|false|false||aidnull|AICDA wt Allele|Finding|false|false||aid
null|AICDA gene|Finding|false|false||aidnull|AID - Artificial insemination by donor|Procedure|false|false||aid
null|dacarbazine/doxorubicin/ifosfamide protocol|Procedure|false|false||aidnull|Aid (attribute)|Modifier|false|false||aid
null|Assisted (qualifier value)|Modifier|false|false||aidnull|Walkers|Device|false|false||walkernull|CANE, INCLUDES CANES OF ALL MATERIALS, ADJUSTABLE OR FIXED, WITH TIP|Device|false|false||canenull|Cane - plant part|Entity|false|false||canenull|Discharge instructions|Finding|false|false||Discharge Instructionsnull|hospital discharge instructions (treatment)|Procedure|false|false||Discharge Instructionsnull|null|Attribute|false|false||Discharge Instructionsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|FBXW7-AS1 gene|Finding|false|false||Dearnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Speech|Finding|false|false||speechnull|Speech assessment|Procedure|false|false||speechnull|Concern|Finding|false|false||concernnull|Acute Ischemic Stroke|Disorder|false|false||ACUTE ISCHEMIC STROKEnull|Admission Level of Care Code - Acute|Finding|false|false||ACUTE
null|Acute - Triage Code|Finding|false|false||ACUTEnull|acute|Time|false|false||ACUTEnull|Ischemic stroke|Disorder|false|false||ISCHEMIC STROKEnull|Ischemic|Finding|false|false||ISCHEMICnull|Cerebrovascular accident|Disorder|false|false||STROKEnull|Stroke (heart beat)|Finding|false|false||STROKEnull|Disease|Disorder|false|false||conditionnull|Logical Condition|Finding|false|false||conditionnull|null|Attribute|false|false||conditionnull|Condition|Modifier|false|false||conditionnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Vessel Positions|Anatomy|false|false||vessel
null|Blood Vessel|Anatomy|false|false||vesselnull|Vessel (unit of presentation)|LabModifier|false|false||vesselnull|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygennull|Oxygen Therapy Care|Procedure|false|false||oxygennull|Oxygen Equipment Location|Modifier|false|false||oxygennull|Nutrients|Drug|false|false||nutrientsnull|Brain Diseases|Disorder|false|false||brainnull|Head>Brain|Anatomy|false|false||brain
null|Brain|Anatomy|false|false||brainnull|clotrimazole|Drug|false|false||clot
null|clotrimazole|Drug|false|false||clotnull|Blood Clot|Finding|false|false||clotnull|Brain Diseases|Disorder|false|false||brainnull|Head>Brain|Anatomy|false|false||brain
null|Brain|Anatomy|false|false||brainnull|part of|Modifier|false|false||part ofnull|Role Class - part|Finding|false|false||partnull|Part|Modifier|false|false||partnull|Part Dosing Unit|LabModifier|false|false||partnull|Document Body|Finding|false|false||bodynull|Structure of body of caudate nucleus|Anatomy|false|false||body
null|Human body structure|Anatomy|false|false||body
null|Body structure|Anatomy|false|false||body
null|Adult human body|Anatomy|false|false||body
null|Whole body|Anatomy|false|false||bodynull|Human body|Subject|false|false||bodynull|Part|Modifier|false|false||partsnull|Document Body|Finding|false|false||bodynull|Structure of body of caudate nucleus|Anatomy|false|false||body
null|Human body structure|Anatomy|false|false||body
null|Body structure|Anatomy|false|false||body
null|Adult human body|Anatomy|false|false||body
null|Whole body|Anatomy|false|false||bodynull|Human body|Subject|false|false||bodynull|Tissue damage|Disorder|false|false||damagenull|Damage|Finding|false|false||damage
null|MAGEE1 gene|Finding|false|false||damagenull|Brain Diseases|Disorder|false|false||brainnull|Head>Brain|Anatomy|false|false||brain
null|Brain|Anatomy|false|false||brainnull|Vascular blood supply|Finding|false|false||blood supply
null|Arterial blood supply|Finding|false|false||blood supplynull|Blood supply aspects|Modifier|false|false||blood supplynull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|In Blood|Finding|false|false||blood
null|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||bloodnull|Supply (process)|Finding|false|false||supply
null|Supply (system)|Finding|false|false||supply
null|supply aspects|Finding|false|false||supplynull|Healthcare supplies|Device|false|false||supplynull|Providing (action)|Event|false|false||supplynull|supply & distribution|LabModifier|false|false||supply
null|Economic supply|LabModifier|false|false||supplynull|Variety (taxon)|Finding|false|false||variety
null|Assortment|Finding|false|false||varietynull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|Brain Diseases|Disorder|false|false||brainnull|Head>Brain|Anatomy|false|false||brain
null|Brain|Anatomy|false|false||brainnull|Evidence of (contextual qualifier)|Finding|false|false||evidence ofnull|Evidence|Finding|false|false||evidencenull|Cerebrovascular accident|Disorder|false|false||strokenull|Stroke (heart beat)|Finding|false|false||strokenull|Transient Cerebral Ischemia|Disorder|false|false||TIA
null|Transient Ischemic Attack|Disorder|false|false||TIAnull|Tacca leontopetaloides|Entity|false|false||TIAnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Relate - vinyl resin|Drug|false|false||relatednull|Role Link Type - related|Finding|false|false||related
null|Related (finding)|Finding|false|false||relatednull|Definitely Related to Intervention|Modifier|false|false||related
null|Relationships|Modifier|false|false||relatednull|Blood pressure finding|Finding|false|false||blood pressure
null|Systemic arterial pressure|Finding|false|false||blood pressure
null|Blood Pressure|Finding|false|false||blood pressurenull|Blood pressure determination|Procedure|false|false||blood pressurenull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|dehydration (Na, H2O)|Disorder|false|false||dehydration
null|Dehydration|Disorder|false|false||dehydrationnull|Dehydration procedure|Procedure|false|false||dehydrationnull|history of alcohol use|Finding|false|false||alcohol use
null|Alcohol consumption|Finding|false|false||alcohol usenull|Alcohols|Drug|false|false||alcohol
null|Alcohols|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcoholnull|Alcohol - Recreational Drug Use Code|Finding|false|false||alcoholnull|Use - dosing instruction imperative|Finding|false|false||use
null|utilization qualifier|Finding|false|false||use
null|Usage|Finding|false|false||usenull|combination - answer to question|Finding|false|false||combinationnull|combination of objects|Entity|false|false||combinationnull|Combined|Modifier|false|false||combinationnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|apixaban|Drug|false|false||apixaban
null|apixaban|Drug|false|false||apixabannull|Twice a day|Time|false|false||twice dailynull|Daily|Time|false|false||dailynull|Vitamin B12 [EPC]|Drug|false|false||Vitamin B12
null|cobalamins|Drug|false|false||Vitamin B12
null|cobalamins|Drug|false|false||Vitamin B12
null|vitamin B12|Drug|false|false||Vitamin B12
null|vitamin B12|Drug|false|false||Vitamin B12
null|vitamin B12|Drug|false|false||Vitamin B12null|VITAMIN B12 MEASUREMENT|Procedure|false|false||Vitamin B12null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|TNFAIP1 wt Allele|Finding|false|false||B12
null|NDUFB3 gene|Finding|false|false||B12
null|TNFAIP1 gene|Finding|false|false||B12null|Daily|Time|false|false||dailynull|Dietary Supplements|Drug|false|false||supplementnull|Supplement - Diet Code Specification Type|Finding|false|false||supplement
null|Supplement|Finding|false|false||supplement
null|Supplement (document)|Finding|false|false||supplementnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Primary Care Physicians|Subject|false|false||primary care physician
null|Primary care provider|Subject|false|false||primary care physiciannull|Location Service Code - Primary Care|Finding|false|false||primary carenull|Primary Health Care|Procedure|false|false||primary carenull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|null|Attribute|false|false||physiciannull|Physicians|Subject|false|false||physiciannull|Cardiologists|Subject|false|false||cardiologistnull|Infrequent|Time|false|false||occasionalnull|null|Attribute|false|false||pausesnull|Pauses|Time|false|false||pausesnull|Cardiac monitoring|Procedure|false|false||cardiac monitoringnull|Cardiac attachment|Finding|false|false||cardiacnull|Heart|Anatomy|false|false||cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||cardiacnull|Preventive monitoring|Procedure|false|false||monitoringnull|null|Event|false|false||monitoringnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Consent Non-Disclosure Reason - Emergency|Finding|false|false||emergency
null|Admission Type - Emergency|Finding|false|false||emergency
null|Referral category - Emergency|Finding|false|false||emergency
null|Emergencies [Disease/Finding]|Finding|false|false||emergency
null|Consent Bypass Reason - Emergency|Finding|false|false||emergency
null|Level of Care - Emergency|Finding|false|false||emergency
null|Certification patient type - Emergency|Finding|false|false||emergency
null|Encounter Admission Source - emergency|Finding|false|false||emergency
null|Patient Class - Emergency|Finding|false|false||emergency
null|Visit Priority Code - Emergency|Finding|false|false||emergencynull|emergency encounter|Procedure|false|false||emergencynull|Specialty Type - Emergency|Title|false|false||emergencynull|Emergency Situation|Phenomenon|false|false||emergencynull|Bale out|Time|false|false||emergencynull|Medical referral type|Finding|false|false||medical
null|Medical|Finding|false|false||medical
null|Medical school type|Finding|false|false||medicalnull|Medical service|Procedure|false|false||medicalnull|Attention - G-code|Finding|false|false||attention
null|Attention|Finding|false|false||attentionnull|Consent Non-Disclosure Reason - Emergency|Finding|false|false||Emergency
null|Admission Type - Emergency|Finding|false|false||Emergency
null|Referral category - Emergency|Finding|false|false||Emergency
null|Emergencies [Disease/Finding]|Finding|false|false||Emergency
null|Consent Bypass Reason - Emergency|Finding|false|false||Emergency
null|Level of Care - Emergency|Finding|false|false||Emergency
null|Certification patient type - Emergency|Finding|false|false||Emergency
null|Encounter Admission Source - emergency|Finding|false|false||Emergency
null|Patient Class - Emergency|Finding|false|false||Emergency
null|Visit Priority Code - Emergency|Finding|false|false||Emergencynull|emergency encounter|Procedure|false|false||Emergencynull|Specialty Type - Emergency|Title|false|false||Emergencynull|Emergency Situation|Phenomenon|false|false||Emergencynull|Bale out|Time|false|false||Emergencynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Clinical Service|Procedure|false|false||Servicesnull|Services|Event|false|false||Servicesnull|Paid Hours|LabModifier|false|false||pay
null|Wages|LabModifier|false|false||paynull|Attention - G-code|Finding|false|false||attention
null|Attention|Finding|false|false||attentionnull|Sudden onset (contextual qualifier) (qualifier value)|Finding|false|false||sudden onsetnull|Sudden onset (attribute)|Time|false|false||sudden onsetnull|Sudden (qualifier value)|Modifier|false|false||suddennull|Onset of (contextual qualifier)|Modifier|false|false||onsetnull|Age of Onset|LabModifier|false|false||onsetnull|Persistence|Finding|false|false||persistencenull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Sudden (qualifier value)|Modifier|false|false||Suddennull|Target Awareness - partial|Finding|false|false||partialnull|Partial|LabModifier|false|false||partialnull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|Low Vision|Disorder|false|false||loss of vision
null|Blindness|Disorder|false|false||loss of visionnull|Unspecified visual loss|Finding|false|false||loss of vision
null|Abnormal vision|Finding|false|false||loss of visionnull|Loss (adaptation)|Finding|false|false||lossnull|Loss (quantitative)|LabModifier|false|false||lossnull|Vision|Finding|false|false||visionnull|null|Attribute|false|false||visionnull|Specialized Stand Alone Plan - Vision|Entity|false|false||visionnull|Sudden (qualifier value)|Modifier|false|false||Suddennull|Loss (adaptation)|Finding|false|false||lossnull|Loss (quantitative)|LabModifier|false|false||lossnull|Ability Question|Finding|false|false||ability tonull|Oral Intake Ability|Finding|false|false||abilitynull|Ability|Subject|false|false||abilitynull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Sudden (qualifier value)|Modifier|false|false||Suddennull|Loss (adaptation)|Finding|false|false||lossnull|Loss (quantitative)|LabModifier|false|false||lossnull|Ability Question|Finding|false|false||ability tonull|Oral Intake Ability|Finding|false|false||abilitynull|Ability|Subject|false|false||abilitynull|Sudden (qualifier value)|Modifier|false|false||Suddennull|Weakness|Finding|false|false||weakness
null|Asthenia|Finding|false|false||weaknessnull|Unilateral|Modifier|false|false||one sidenull|Side|Modifier|false|false||sidenull|Document Body|Finding|false|false||bodynull|Structure of body of caudate nucleus|Anatomy|false|false||body
null|Human body structure|Anatomy|false|false||body
null|Body structure|Anatomy|false|false||body
null|Adult human body|Anatomy|false|false||body
null|Whole body|Anatomy|false|false||bodynull|Human body|Subject|false|false||bodynull|Sudden (qualifier value)|Modifier|false|false||Suddennull|Unilateral|Modifier|false|false||one sidenull|Side|Modifier|false|false||sidenull|FANCONI ANEMIA, COMPLEMENTATION GROUP E|Disorder|false|false||facenull|FANCE wt Allele|Finding|false|false||face
null|FANCE gene|Finding|false|false||face
null|ELOVL6 gene|Finding|false|false||facenull|Head>Face|Anatomy|false|false||face
null|Face|Anatomy|false|false||facenull|Face (spatial concept)|Modifier|false|false||facenull|Sudden (qualifier value)|Modifier|false|false||Suddennull|Numbness|Finding|false|false||loss of sensationnull|Loss (adaptation)|Finding|false|false||lossnull|Loss (quantitative)|LabModifier|false|false||lossnull|Observation of Sensation|Finding|false|false||sensation
null|Sensory perception|Finding|false|false||sensationnull|sensory exam|Procedure|false|false||sensationnull|Sensation quality|Modifier|false|false||sensationnull|Unilateral|Modifier|false|false||one sidenull|Side|Modifier|false|false||sidenull|Document Body|Finding|false|false||bodynull|Structure of body of caudate nucleus|Anatomy|false|false||body
null|Human body structure|Anatomy|false|false||body
null|Body structure|Anatomy|false|false||body
null|Adult human body|Anatomy|false|false||body
null|Whole body|Anatomy|false|false||bodynull|Human body|Subject|false|false||bodynull|Neurology Team|Title|false|false||Neurology Teamnull|Neurology speciality|Title|false|false||Neurologynull|Team|Subject|false|false||Teamnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions