 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|26,30
No|31,33
:|33,34
_|37,38
_|38,39
_|39,40
<EOL>|40,41
<EOL>|42,43
Admission|43,52
Date|53,57
:|57,58
_|60,61
_|61,62
_|62,63
Discharge|77,86
Date|87,91
:|91,92
_|95,96
_|96,97
_|97,98
<EOL>|98,99
<EOL>|100,101
Date|101,105
of|106,108
Birth|109,114
:|114,115
_|117,118
_|118,119
_|119,120
Sex|133,136
:|136,137
F|140,141
<EOL>|141,142
<EOL>|143,144
Service|144,151
:|151,152
NEUROSURGERY|153,165
<EOL>|165,166
<EOL>|167,168
Allergies|168,177
:|177,178
<EOL>|179,180
Penicillins|180,191
<EOL>|191,192
<EOL>|193,194
Attending|194,203
:|203,204
_|205,206
_|206,207
_|207,208
<EOL>|208,209
<EOL>|210,211
Chief|211,216
Complaint|217,226
:|226,227
<EOL>|227,228
Left|228,232
hand|233,237
and|238,241
face|242,246
numbness|247,255
,|255,256
left|257,261
hand|262,266
weakness|267,275
and|276,279
clumsiness|280,290
,|290,291
<EOL>|292,293
fever|293,298
,|298,299
and|300,303
headache|304,312
.|312,313
<EOL>|313,314
<EOL>|315,316
Major|316,321
Surgical|322,330
or|331,333
Invasive|334,342
Procedure|343,352
:|352,353
<EOL>|353,354
Right|354,359
parietal|360,368
craniotomy|369,379
for|380,383
abscess|384,391
incision|392,400
and|401,404
drainage|405,413
.|413,414
<EOL>|414,415
<EOL>|416,417
History|417,424
of|425,427
Present|428,435
Illness|436,443
:|443,444
<EOL>|444,445
Mrs.|445,449
_|450,451
_|451,452
_|452,453
is|454,456
a|457,458
_|459,460
_|460,461
_|461,462
y|463,464
/|464,465
o|465,466
F|467,468
from|469,473
_|474,475
_|475,476
_|476,477
with|478,482
history|483,490
of|491,493
MS|494,496
<EOL>|497,498
presents|498,506
with|507,511
headaches|512,521
and|522,525
left|526,530
hand|531,535
clumsiness|536,546
.|546,547
Patient|548,555
states|556,562
<EOL>|563,564
that|564,568
her|569,572
headaches|573,582
first|583,588
presented|589,598
on|599,601
_|602,603
_|603,604
_|604,605
of|606,608
this|609,613
week|614,618
in|619,621
<EOL>|622,623
which|623,628
she|629,632
did|633,636
not|637,640
think|641,646
much|647,651
of|652,654
,|654,655
but|656,659
on|660,662
_|663,664
_|664,665
_|665,666
,|666,667
developed|668,677
left|678,682
<EOL>|683,684
hand|684,688
clumsiness|689,699
.|699,700
She|701,704
states|705,711
that|712,716
she|717,720
had|721,724
difficulty|725,735
with|736,740
<EOL>|741,742
grasping|742,750
objects|751,758
and|759,762
using|763,768
her|769,772
fingers|773,780
.|780,781
She|782,785
also|786,790
reported|791,799
some|800,804
<EOL>|805,806
numbness|806,814
in|815,817
the|818,821
hand|822,826
.|826,827
Today|828,833
,|833,834
she|835,838
presented|839,848
to|849,851
the|852,855
ED|856,858
because|859,866
she|867,870
<EOL>|871,872
was|872,875
found|876,881
to|882,884
have|885,889
a|890,891
temperature|892,903
of|904,906
101.7|907,912
in|913,915
which|916,921
she|922,925
took|926,930
<EOL>|931,932
Tylenol|932,939
and|940,943
was|944,947
normothermic|948,960
after|961,966
.|966,967
Once|968,972
in|973,975
the|976,979
ED|980,982
,|982,983
patient|984,991
was|992,995
<EOL>|996,997
seen|997,1001
by|1002,1004
neurology|1005,1014
who|1015,1018
recommended|1019,1030
an|1031,1033
MRI|1034,1037
head|1038,1042
.|1042,1043
MRI|1044,1047
head|1048,1052
revealed|1053,1061
<EOL>|1062,1063
a|1063,1064
R|1065,1066
parietal|1067,1075
lesion|1076,1082
concerning|1083,1093
for|1094,1097
MS|1098,1100
,|1100,1101
metastatic|1102,1112
disease|1113,1120
,|1120,1121
or|1122,1124
<EOL>|1125,1126
abscess|1126,1133
.|1133,1134
Neurosurgery|1135,1147
was|1148,1151
consulted|1152,1161
for|1162,1165
further|1166,1173
evaluation|1174,1184
.|1184,1185
<EOL>|1185,1186
<EOL>|1186,1187
She|1187,1190
reports|1191,1198
a|1199,1200
mild|1201,1205
headache|1206,1214
,|1214,1215
numbness|1216,1224
on|1225,1227
the|1228,1231
left|1232,1236
side|1237,1241
of|1242,1244
face|1245,1249
<EOL>|1250,1251
and|1251,1254
difficulty|1255,1265
using|1266,1271
her|1272,1275
left|1276,1280
hand|1281,1285
.|1285,1286
She|1287,1290
denies|1291,1297
any|1298,1301
recent|1302,1308
travel|1309,1315
<EOL>|1316,1317
outside|1317,1324
of|1325,1327
_|1328,1329
_|1329,1330
_|1330,1331
and|1332,1335
the|1336,1339
_|1340,1341
_|1341,1342
_|1342,1343
.|1343,1344
or|1345,1347
ingesting|1348,1357
any|1358,1361
raw|1362,1365
or|1366,1368
uncooked|1369,1377
<EOL>|1378,1379
meats|1379,1384
.|1384,1385
She|1386,1389
also|1390,1394
denies|1395,1401
any|1402,1405
changes|1406,1413
in|1414,1416
vision|1417,1423
,|1423,1424
dysarthria|1425,1435
,|1435,1436
<EOL>|1437,1438
weakness|1438,1446
,|1446,1447
nausea|1448,1454
,|1454,1455
vomitting|1456,1465
,|1465,1466
diarrhea|1467,1475
,|1475,1476
cough|1477,1482
,|1482,1483
or|1484,1486
chills|1487,1493
.|1493,1494
<EOL>|1494,1495
<EOL>|1495,1496
<EOL>|1497,1498
Past|1498,1502
Medical|1503,1510
History|1511,1518
:|1518,1519
<EOL>|1519,1520
Multiple|1520,1528
sclerosis|1529,1538
<EOL>|1538,1539
<EOL>|1540,1541
Social|1541,1547
History|1548,1555
:|1555,1556
<EOL>|1556,1557
_|1557,1558
_|1558,1559
_|1559,1560
<EOL>|1560,1561
Family|1561,1567
History|1568,1575
:|1575,1576
<EOL>|1576,1577
Mother|1577,1583
with|1584,1588
pancreatic|1589,1599
cancer|1600,1606
,|1606,1607
brother|1608,1615
-|1615,1616
lung|1616,1620
cancer|1621,1627
,|1627,1628
two|1629,1632
sisters|1633,1640
<EOL>|1641,1642
with|1642,1646
brain|1647,1652
cancer|1653,1659
.|1659,1660
<EOL>|1660,1661
<EOL>|1661,1662
<EOL>|1663,1664
Physical|1664,1672
Exam|1673,1677
:|1677,1678
<EOL>|1678,1679
PHYSICAL|1679,1687
EXAM|1688,1692
ON|1693,1695
ADMISSION|1696,1705
:|1705,1706
<EOL>|1706,1707
O|1707,1708
:|1708,1709
T|1710,1711
:|1711,1712
99|1712,1714
BP|1716,1718
:|1718,1719
160|1719,1722
/|1722,1723
102|1723,1726
HR|1728,1730
:|1730,1731
81|1732,1734
R|1738,1739
:|1739,1740
16|1741,1743
O2Sats|1747,1753
:|1753,1754
97|1755,1757
%|1757,1758
RA|1759,1761
<EOL>|1761,1762
Gen|1762,1765
:|1765,1766
WD|1767,1769
/|1769,1770
WN|1770,1772
,|1772,1773
comfortable|1774,1785
,|1785,1786
NAD|1787,1790
.|1790,1791
<EOL>|1791,1792
HEENT|1792,1797
:|1797,1798
atraumatic|1799,1809
,|1809,1810
normocephalic|1811,1824
<EOL>|1824,1825
Pupils|1825,1831
:|1831,1832
4|1833,1834
-|1834,1835
3mm|1835,1838
bilaterally|1839,1850
EOMs|1859,1863
:|1863,1864
intact|1865,1871
<EOL>|1871,1872
<EOL>|1872,1873
Neuro|1873,1878
:|1878,1879
<EOL>|1879,1880
Mental|1880,1886
status|1887,1893
:|1893,1894
Awake|1895,1900
and|1901,1904
alert|1905,1910
,|1910,1911
cooperative|1912,1923
with|1924,1928
exam|1929,1933
,|1933,1934
normal|1935,1941
<EOL>|1941,1942
affect|1942,1948
.|1948,1949
<EOL>|1949,1950
Orientation|1950,1961
:|1961,1962
Oriented|1963,1971
to|1972,1974
person|1975,1981
,|1981,1982
place|1983,1988
,|1988,1989
and|1990,1993
date|1994,1998
.|1998,1999
<EOL>|1999,2000
Recall|2000,2006
:|2006,2007
_|2008,2009
_|2009,2010
_|2010,2011
objects|2012,2019
at|2020,2022
5|2023,2024
minutes|2025,2032
.|2032,2033
<EOL>|2033,2034
Language|2034,2042
:|2042,2043
Speech|2044,2050
fluent|2051,2057
with|2058,2062
good|2063,2067
comprehension|2068,2081
and|2082,2085
repetition|2086,2096
.|2096,2097
<EOL>|2097,2098
Naming|2098,2104
intact|2105,2111
.|2111,2112
No|2113,2115
dysarthria|2116,2126
or|2127,2129
paraphasic|2130,2140
errors|2141,2147
.|2147,2148
<EOL>|2148,2149
<EOL>|2149,2150
Cranial|2150,2157
Nerves|2158,2164
:|2164,2165
<EOL>|2165,2166
I|2166,2167
:|2167,2168
Not|2169,2172
tested|2173,2179
<EOL>|2179,2180
II|2180,2182
:|2182,2183
Pupils|2184,2190
equally|2191,2198
round|2199,2204
and|2205,2208
reactive|2209,2217
to|2218,2220
light|2221,2226
,|2226,2227
4|2228,2229
to|2230,2232
3|2233,2234
<EOL>|2234,2235
mm|2235,2237
bilaterally|2238,2249
.|2249,2250
Visual|2251,2257
fields|2258,2264
are|2265,2268
full|2269,2273
to|2274,2276
confrontation|2277,2290
.|2290,2291
<EOL>|2291,2292
III|2292,2295
,|2295,2296
IV|2297,2299
,|2299,2300
VI|2301,2303
:|2303,2304
Extraocular|2305,2316
movements|2317,2326
intact|2327,2333
bilaterally|2334,2345
without|2346,2353
<EOL>|2353,2354
nystagmus|2354,2363
.|2363,2364
<EOL>|2364,2365
V|2365,2366
,|2366,2367
VII|2368,2371
:|2371,2372
Facial|2373,2379
strength|2380,2388
and|2389,2392
sensation|2393,2402
intact|2403,2409
and|2410,2413
symmetric|2414,2423
.|2423,2424
<EOL>|2424,2425
VIII|2425,2429
:|2429,2430
Hearing|2431,2438
intact|2439,2445
to|2446,2448
voice|2449,2454
.|2454,2455
<EOL>|2455,2456
IX|2456,2458
,|2458,2459
X|2460,2461
:|2461,2462
Palatal|2463,2470
elevation|2471,2480
symmetrical|2481,2492
.|2492,2493
<EOL>|2493,2494
XI|2494,2496
:|2496,2497
Sternocleidomastoid|2498,2517
and|2518,2521
trapezius|2522,2531
normal|2532,2538
bilaterally|2539,2550
.|2550,2551
<EOL>|2551,2552
XII|2552,2555
:|2555,2556
Tongue|2557,2563
midline|2564,2571
without|2572,2579
fasciculations|2580,2594
.|2594,2595
<EOL>|2595,2596
<EOL>|2596,2597
Motor|2597,2602
:|2602,2603
Normal|2604,2610
bulk|2611,2615
and|2616,2619
tone|2620,2624
bilaterally|2625,2636
.|2636,2637
No|2638,2640
abnormal|2641,2649
movements|2650,2659
,|2659,2660
<EOL>|2660,2661
tremors|2661,2668
.|2668,2669
Strength|2670,2678
L|2679,2680
FI|2681,2683
_|2684,2685
_|2685,2686
_|2686,2687
,|2687,2688
otherwise|2689,2698
full|2699,2703
power|2704,2709
_|2710,2711
_|2711,2712
_|2712,2713
<EOL>|2714,2715
throughout|2715,2725
.|2725,2726
<EOL>|2726,2727
No|2727,2729
pronator|2730,2738
drift|2739,2744
<EOL>|2744,2745
<EOL>|2745,2746
Sensation|2746,2755
:|2755,2756
Intact|2757,2763
to|2764,2766
light|2767,2772
touch|2773,2778
<EOL>|2778,2779
<EOL>|2779,2780
PHYSICAL|2780,2788
EXAM|2789,2793
ON|2794,2796
DISCHARGE|2797,2806
:|2806,2807
<EOL>|2807,2808
<EOL>|2808,2809
T|2809,2810
:|2810,2811
98.1|2811,2815
BP|2817,2819
:|2819,2820
133|2820,2823
/|2823,2824
95|2824,2826
HR|2828,2830
:|2830,2831
95|2832,2834
RR|2835,2837
:|2837,2838
18|2839,2841
O2Sats|2842,2848
:|2848,2849
98|2850,2852
%|2852,2853
RA|2854,2856
<EOL>|2856,2857
Gen|2857,2860
:|2860,2861
WD|2862,2864
/|2864,2865
WN|2865,2867
,|2867,2868
comfortable|2869,2880
,|2880,2881
NAD|2882,2885
.|2885,2886
<EOL>|2886,2887
HEENT|2887,2892
:|2892,2893
atraumatic|2894,2904
,|2904,2905
normocephalic|2906,2919
,|2919,2920
with|2921,2925
right|2926,2931
craniotomy|2932,2942
<EOL>|2943,2944
incision|2944,2952
.|2952,2953
<EOL>|2953,2954
Pupils|2954,2960
:|2960,2961
4|2962,2963
-|2963,2964
3mm|2964,2967
bilaterally|2968,2979
,|2979,2980
EOMs|2981,2985
:|2985,2986
intact|2987,2993
<EOL>|2993,2994
<EOL>|2994,2995
Neuro|2995,3000
:|3000,3001
<EOL>|3001,3002
Mental|3002,3008
status|3009,3015
:|3015,3016
Awake|3017,3022
and|3023,3026
alert|3027,3032
,|3032,3033
cooperative|3034,3045
with|3046,3050
exam|3051,3055
,|3055,3056
normal|3057,3063
<EOL>|3063,3064
affect|3064,3070
.|3070,3071
<EOL>|3071,3072
Orientation|3072,3083
:|3083,3084
Oriented|3085,3093
to|3094,3096
person|3097,3103
,|3103,3104
place|3105,3110
,|3110,3111
and|3112,3115
date|3116,3120
.|3120,3121
<EOL>|3121,3122
Recall|3122,3128
:|3128,3129
_|3130,3131
_|3131,3132
_|3132,3133
objects|3134,3141
at|3142,3144
5|3145,3146
minutes|3147,3154
.|3154,3155
<EOL>|3155,3156
Language|3156,3164
:|3164,3165
Speech|3166,3172
fluent|3173,3179
with|3180,3184
good|3185,3189
comprehension|3190,3203
and|3204,3207
repetition|3208,3218
.|3218,3219
<EOL>|3219,3220
Naming|3220,3226
intact|3227,3233
.|3233,3234
No|3235,3237
dysarthria|3238,3248
or|3249,3251
paraphasic|3252,3262
errors|3263,3269
.|3269,3270
<EOL>|3270,3271
<EOL>|3271,3272
Cranial|3272,3279
Nerves|3280,3286
:|3286,3287
<EOL>|3287,3288
I|3288,3289
:|3289,3290
Not|3291,3294
tested|3295,3301
<EOL>|3301,3302
II|3302,3304
:|3304,3305
Pupils|3306,3312
equally|3313,3320
round|3321,3326
and|3327,3330
reactive|3331,3339
to|3340,3342
light|3343,3348
,|3348,3349
4|3350,3351
to|3352,3354
3|3355,3356
mm|3357,3359
<EOL>|3360,3361
bilaterally|3361,3372
.|3372,3373
Visual|3374,3380
fields|3381,3387
are|3388,3391
full|3392,3396
to|3397,3399
confrontation|3400,3413
.|3413,3414
<EOL>|3414,3415
III|3415,3418
,|3418,3419
IV|3420,3422
,|3422,3423
VI|3424,3426
:|3426,3427
Extraocular|3428,3439
movements|3440,3449
intact|3450,3456
bilaterally|3457,3468
without|3469,3476
<EOL>|3476,3477
nystagmus|3477,3486
.|3486,3487
<EOL>|3487,3488
V|3488,3489
,|3489,3490
VII|3491,3494
:|3494,3495
Facial|3496,3502
strength|3503,3511
and|3512,3515
sensation|3516,3525
intact|3526,3532
and|3533,3536
symmetric|3537,3546
.|3546,3547
<EOL>|3547,3548
VIII|3548,3552
:|3552,3553
Hearing|3554,3561
intact|3562,3568
to|3569,3571
voice|3572,3577
.|3577,3578
<EOL>|3578,3579
IX|3579,3581
,|3581,3582
X|3583,3584
:|3584,3585
Palatal|3586,3593
elevation|3594,3603
symmetrical|3604,3615
.|3615,3616
<EOL>|3616,3617
XI|3617,3619
:|3619,3620
Sternocleidomastoid|3621,3640
and|3641,3644
trapezius|3645,3654
normal|3655,3661
bilaterally|3662,3673
.|3673,3674
<EOL>|3674,3675
XII|3675,3678
:|3678,3679
Tongue|3680,3686
midline|3687,3694
without|3695,3702
fasciculations|3703,3717
.|3717,3718
<EOL>|3718,3719
<EOL>|3719,3720
Motor|3720,3725
:|3725,3726
Normal|3727,3733
bulk|3734,3738
and|3739,3742
tone|3743,3747
bilaterally|3748,3759
.|3759,3760
No|3761,3763
abnormal|3764,3772
<EOL>|3773,3774
movements|3774,3783
,|3783,3784
tremors|3784,3791
.|3791,3792
Strength|3793,3801
L|3802,3803
FI|3804,3806
_|3807,3808
_|3808,3809
_|3809,3810
,|3810,3811
otherwise|3812,3821
full|3822,3826
power|3827,3832
_|3833,3834
_|3834,3835
_|3835,3836
<EOL>|3837,3838
throughout|3838,3848
.|3848,3849
<EOL>|3849,3850
No|3850,3852
pronator|3853,3861
drift|3862,3867
<EOL>|3867,3868
<EOL>|3868,3869
Sensation|3869,3878
:|3878,3879
Intact|3880,3886
to|3887,3889
light|3890,3895
touch|3896,3901
<EOL>|3901,3902
<EOL>|3902,3903
<EOL>|3904,3905
Pertinent|3905,3914
Results|3915,3922
:|3922,3923
<EOL>|3923,3924
_|3924,3925
_|3925,3926
_|3926,3927
MRI|3928,3931
HEAD|3932,3936
W|3937,3938
/|3938,3939
WO|3939,3941
CONTRAST|3942,3950
<EOL>|3951,3952
IMPRESSION|3952,3962
:|3962,3963
<EOL>|3964,3965
<EOL>|3967,3968
1.|3968,3970
Ring|3972,3976
-|3976,3977
enhancing|3977,3986
lesion|3987,3993
identified|3994,4004
in|4005,4007
the|4008,4011
area|4012,4016
of|4017,4019
the|4020,4023
right|4024,4029
<EOL>|4030,4031
precentral|4031,4041
<EOL>|4042,4043
sulcus|4043,4049
frontal|4050,4057
lobe|4058,4062
,|4062,4063
with|4064,4068
associated|4069,4079
vasogenic|4080,4089
edema|4090,4095
,|4095,4096
restricted|4097,4107
<EOL>|4108,4109
diffusion|4109,4118
,|4118,4119
possibly|4120,4128
consistent|4129,4139
with|4140,4144
an|4145,4147
abscess|4148,4155
,|4155,4156
other|4157,4162
entities|4163,4171
<EOL>|4172,4173
can|4173,4176
not|4176,4179
be|4180,4182
completely|4183,4193
ruled|4194,4199
out|4200,4203
such|4204,4208
as|4209,4211
metastases|4212,4222
or|4223,4225
primary|4226,4233
<EOL>|4234,4235
brain|4235,4240
neoplasm|4241,4249
.|4249,4250
<EOL>|4251,4252
<EOL>|4254,4255
2.|4255,4257
Multiple|4259,4267
FLAIR|4268,4273
and|4274,4277
T2|4278,4280
hyperintense|4281,4293
lesions|4294,4301
in|4302,4304
the|4305,4308
<EOL>|4309,4310
subcortical|4310,4321
white|4322,4327
matter|4328,4334
along|4335,4340
the|4341,4344
callososeptal|4345,4358
region|4359,4365
,|4365,4366
<EOL>|4367,4368
consistent|4368,4378
with|4379,4383
known|4384,4389
multiple|4390,4398
sclerosis|4399,4408
disease|4409,4416
.|4416,4417
<EOL>|4418,4419
<EOL>|4419,4420
_|4420,4421
_|4421,4422
_|4422,4423
MRI|4424,4427
HEAD|4428,4432
W|4433,4434
/|4434,4435
CONTRAST|4436,4444
<EOL>|4445,4446
IMPRESSION|4446,4456
:|4456,4457
Unchanged|4459,4468
ring|4469,4473
-|4473,4474
enhancing|4474,4483
lesion|4484,4490
identified|4491,4501
in|4502,4504
the|4505,4508
<EOL>|4509,4510
area|4510,4514
of|4515,4517
the|4518,4521
<EOL>|4522,4523
right|4523,4528
precentral|4529,4539
sulcus|4540,4546
of|4547,4549
the|4550,4553
frontal|4554,4561
lobe|4562,4566
,|4566,4567
with|4568,4572
associated|4573,4583
<EOL>|4584,4585
vasogenic|4585,4594
edema|4595,4600
.|4600,4601
The|4603,4606
differential|4607,4619
diagnosis|4620,4629
again|4630,4635
includes|4636,4644
<EOL>|4645,4646
possible|4646,4654
abscess|4655,4662
,|4662,4663
other|4664,4669
entities|4670,4678
,|4678,4679
however|4680,4687
,|4687,4688
can|4689,4692
not|4692,4695
be|4696,4698
completely|4699,4709
<EOL>|4710,4711
excluded|4711,4719
.|4719,4720
<EOL>|4721,4722
<EOL>|4722,4723
_|4723,4724
_|4724,4725
_|4725,4726
NON|4727,4730
CONTRAST|4731,4739
HEAD|4740,4744
CT|4745,4747
<EOL>|4748,4749
IMPRESSION|4749,4759
:|4759,4760
<EOL>|4761,4762
<EOL>|4764,4765
1.|4765,4767
Status|4769,4775
post|4776,4780
right|4781,4786
parietal|4787,4795
craniotomy|4796,4806
with|4807,4811
mixed|4812,4817
density|4818,4825
<EOL>|4826,4827
lesion|4827,4833
in|4834,4836
the|4837,4840
<EOL>|4841,4842
right|4842,4847
precentral|4848,4858
sulcus|4859,4865
and|4866,4869
surrounding|4870,4881
edema|4882,4887
not|4888,4891
significantly|4892,4905
<EOL>|4906,4907
changed|4907,4914
from|4915,4919
prior|4920,4925
MR|4926,4928
of|4929,4931
_|4932,4933
_|4933,4934
_|4934,4935
allowing|4936,4944
for|4945,4948
<EOL>|4949,4950
difference|4950,4960
in|4961,4963
technique|4964,4973
.|4973,4974
<EOL>|4976,4977
<EOL>|4979,4980
2|4980,4981
.|4981,4982
No|4984,4986
acute|4987,4992
intracranial|4993,5005
hemorrhage|5006,5016
or|5017,5019
major|5020,5025
vascular|5026,5034
<EOL>|5035,5036
territorial|5036,5047
infarct|5048,5055
.|5055,5056
<EOL>|5058,5059
<EOL>|5061,5062
3.|5062,5064
Bifrontal|5066,5075
subcortical|5076,5087
white|5088,5093
matter|5094,5100
hypodensities|5101,5114
compatible|5115,5125
<EOL>|5126,5127
with|5127,5131
<EOL>|5132,5133
underlying|5133,5143
multiple|5144,5152
sclerosis|5153,5162
.|5162,5163
<EOL>|5165,5166
<EOL>|5166,5167
_|5167,5168
_|5168,5169
_|5169,5170
2|5171,5172
:|5172,5173
37|5173,5175
am|5176,5178
CSF|5179,5182
;|5182,5183
SPINAL|5183,5189
FLUID|5190,5195
TUBE|5201,5205
#|5206,5207
1|5207,5208
.|5208,5209
<EOL>|5210,5211
<EOL>|5211,5212
GRAM|5215,5219
STAIN|5220,5225
(|5226,5227
Final|5227,5232
_|5233,5234
_|5234,5235
_|5235,5236
:|5236,5237
<EOL>|5238,5239
NO|5245,5247
POLYMORPHONUCLEAR|5248,5265
LEUKOCYTES|5266,5276
SEEN|5277,5281
.|5281,5282
<EOL>|5283,5284
NO|5290,5292
MICROORGANISMS|5293,5307
SEEN|5308,5312
.|5312,5313
<EOL>|5314,5315
This|5321,5325
is|5326,5328
a|5329,5330
concentrated|5331,5343
smear|5344,5349
made|5350,5354
by|5355,5357
cytospin|5358,5366
method|5367,5373
,|5373,5374
<EOL>|5375,5376
please|5376,5382
refer|5383,5388
to|5389,5391
<EOL>|5391,5392
hematology|5398,5408
for|5409,5412
a|5413,5414
quantitative|5415,5427
white|5428,5433
blood|5434,5439
cell|5440,5444
count|5445,5450
.|5450,5451
.|5451,5452
<EOL>|5453,5454
<EOL>|5454,5455
FLUID|5458,5463
CULTURE|5464,5471
(|5472,5473
Preliminary|5473,5484
)|5484,5485
:|5485,5486
NO|5490,5492
GROWTH|5493,5499
.|5499,5500
<EOL>|5500,5501
<EOL>|5501,5502
<EOL>|5503,5504
Brief|5504,5509
Hospital|5510,5518
Course|5519,5525
:|5525,5526
<EOL>|5526,5527
Mrs.|5527,5531
_|5532,5533
_|5533,5534
_|5534,5535
presented|5536,5545
to|5546,5548
the|5549,5552
_|5553,5554
_|5554,5555
_|5555,5556
Emergency|5557,5566
Department|5567,5577
on|5578,5580
<EOL>|5581,5582
_|5582,5583
_|5583,5584
_|5584,5585
with|5586,5590
left|5591,5595
-|5595,5596
sided|5596,5601
numbness|5602,5610
of|5611,5613
her|5614,5617
hand|5618,5622
and|5623,5626
face|5627,5631
and|5632,5635
left|5636,5640
<EOL>|5641,5642
hand|5642,5646
clumsiness|5647,5657
.|5657,5658
She|5660,5663
was|5664,5667
evaluated|5668,5677
in|5678,5680
the|5681,5684
ED|5685,5687
and|5688,5691
initially|5692,5701
<EOL>|5702,5703
believed|5703,5711
to|5712,5714
have|5715,5719
an|5720,5722
MS|5723,5725
flare|5726,5731
and|5732,5735
she|5736,5739
was|5740,5743
evaluted|5744,5752
by|5753,5755
Neurology|5756,5765
<EOL>|5766,5767
service|5767,5774
which|5775,5780
resulted|5781,5789
in|5790,5792
the|5793,5796
recommendation|5797,5811
for|5812,5815
an|5816,5818
MRI|5819,5822
brain|5823,5828
.|5828,5829
<EOL>|5831,5832
The|5832,5835
MRI|5836,5839
was|5840,5843
read|5844,5848
to|5849,5851
demonstrate|5852,5863
a|5864,5865
right|5866,5871
parietal|5872,5880
lesion|5881,5887
<EOL>|5888,5889
concerning|5889,5899
for|5900,5903
MS|5904,5906
,|5906,5907
metastatic|5908,5918
disease|5919,5926
or|5927,5929
abscess|5930,5937
.|5937,5938
She|5939,5942
was|5943,5946
<EOL>|5947,5948
admitted|5948,5956
to|5957,5959
Neurosurgery|5960,5972
for|5973,5976
further|5977,5984
evaluation|5985,5995
and|5996,5999
treatment|6000,6009
.|6009,6010
<EOL>|6012,6013
<EOL>|6013,6014
On|6014,6016
_|6017,6018
_|6018,6019
_|6019,6020
,|6020,6021
Mrs.|6022,6026
_|6027,6028
_|6028,6029
_|6029,6030
was|6031,6034
taken|6035,6040
to|6041,6043
the|6044,6047
OR|6048,6050
for|6051,6054
a|6055,6056
right|6057,6062
<EOL>|6063,6064
parietal|6064,6072
craniotomy|6073,6083
with|6084,6088
cordisectomy|6089,6101
,|6101,6102
drainage|6103,6111
and|6112,6115
irrigation|6116,6126
<EOL>|6127,6128
of|6128,6130
brain|6131,6136
abscess|6137,6144
.|6144,6145
She|6146,6149
tolerated|6150,6159
the|6160,6163
procedure|6164,6173
well|6174,6178
.|6178,6179
She|6180,6183
was|6184,6187
<EOL>|6188,6189
taken|6189,6194
to|6195,6197
PACU|6198,6202
to|6203,6205
recover|6206,6213
then|6214,6218
to|6219,6221
the|6222,6225
ICU|6226,6229
.|6229,6230
ID|6231,6233
recommmend|6234,6244
<EOL>|6245,6246
Vancomycin|6246,6256
and|6257,6260
Meropenem|6261,6270
.|6270,6271
Gram|6272,6276
stain|6277,6282
PRELIM|6283,6289
:|6289,6290
gram|6291,6295
negative|6296,6304
rods|6305,6309
<EOL>|6310,6311
and|6311,6314
gram|6315,6319
positive|6320,6328
cocci|6329,6334
in|6335,6337
pairs|6338,6343
and|6344,6347
chains|6348,6354
.|6354,6355
Post|6356,6360
operative|6361,6370
head|6371,6375
<EOL>|6376,6377
CT|6377,6379
showed|6380,6386
post|6387,6391
operative|6392,6401
changes|6402,6409
.|6409,6410
On|6411,6413
post|6414,6418
operative|6419,6428
exam|6429,6433
she|6434,6437
had|6438,6441
<EOL>|6442,6443
left|6443,6447
arm|6448,6451
weakness|6452,6460
.|6460,6461
<EOL>|6462,6463
<EOL>|6463,6464
On|6464,6466
_|6467,6468
_|6468,6469
_|6469,6470
the|6471,6474
patient|6475,6482
continued|6483,6492
on|6493,6495
vancomycin|6496,6506
and|6507,6510
Meropenem|6511,6520
.|6520,6521
<EOL>|6522,6523
WBC|6523,6526
was|6527,6530
elevated|6531,6539
to|6540,6542
19.0|6543,6547
from|6548,6552
15.7|6553,6557
on|6558,6560
_|6561,6562
_|6562,6563
_|6563,6564
.|6564,6565
She|6566,6569
was|6570,6573
<EOL>|6574,6575
transferred|6575,6586
to|6587,6589
the|6590,6593
floor|6594,6599
.|6599,6600
Left|6601,6605
arm|6606,6609
weakness|6610,6618
was|6619,6622
slightly|6623,6631
<EOL>|6632,6633
improved.|6633,6642
the|6643,6646
patient|6647,6654
reported|6655,6663
lethargy|6664,6672
and|6673,6676
left|6677,6681
leg|6682,6685
weakness|6686,6694
.|6694,6695
<EOL>|6696,6697
on|6697,6699
exam|6700,6704
the|6705,6708
patient|6709,6716
was|6717,6720
sleepy|6721,6727
but|6728,6731
awake|6732,6737
.|6737,6738
she|6740,6743
was|6744,6747
oriented|6748,6756
to|6757,6759
<EOL>|6760,6761
person|6761,6767
place|6768,6773
and|6774,6777
time|6778,6782
.|6782,6783
right|6785,6790
sided|6791,6796
strength|6797,6805
was|6806,6809
_|6810,6811
_|6811,6812
_|6812,6813
and|6814,6817
left|6818,6822
<EOL>|6823,6824
upper|6824,6829
extremity|6830,6839
was|6840,6843
_|6844,6845
_|6845,6846
_|6846,6847
and|6848,6851
left|6852,6856
lower|6857,6862
extremity|6863,6872
was|6873,6876
full|6877,6881
except|6882,6888
<EOL>|6889,6890
for|6890,6893
IP|6894,6896
which|6897,6902
was|6903,6906
5|6907,6908
-|6908,6909
.|6909,6910
A|6911,6912
stat|6913,6917
NCHCT|6918,6923
was|6924,6927
performed|6928,6937
which|6938,6943
was|6944,6947
<EOL>|6948,6949
stable|6949,6955
.|6955,6956
<EOL>|6956,6957
<EOL>|6957,6958
On|6958,6960
_|6961,6962
_|6962,6963
_|6963,6964
,|6964,6965
consent|6966,6973
for|6974,6977
picc|6978,6982
line|6983,6987
placement|6988,6997
obtained|6998,7006
,|7006,7007
picc|7008,7012
line|7013,7017
<EOL>|7018,7019
placed|7019,7025
by|7026,7028
IV|7029,7031
nurse|7032,7037
.|7037,7038
She|7039,7042
will|7043,7047
continue|7048,7056
with|7057,7061
vanco|7062,7067
and|7068,7071
meropenum|7072,7081
<EOL>|7082,7083
IV|7083,7085
.|7085,7086
Final|7087,7092
abcess|7093,7099
culture|7100,7107
result|7108,7114
is|7115,7117
still|7118,7123
pending|7124,7131
.|7131,7132
Exam|7133,7137
remains|7138,7145
<EOL>|7146,7147
stable|7147,7153
.|7153,7154
<EOL>|7155,7156
<EOL>|7156,7157
On|7157,7159
_|7160,7161
_|7161,7162
_|7162,7163
_|7164,7165
_|7165,7166
_|7166,7167
evaluated|7168,7177
the|7178,7181
patient|7182,7189
and|7190,7193
found|7194,7199
that|7200,7204
she|7205,7208
continues|7209,7218
<EOL>|7219,7220
to|7220,7222
have|7223,7227
an|7228,7230
unsteady|7231,7239
gait|7240,7244
and|7245,7248
would|7249,7254
not|7255,7258
be|7259,7261
safe|7262,7266
to|7267,7269
go|7270,7272
home|7273,7277
.|7277,7278
They|7280,7284
<EOL>|7285,7286
planned|7286,7293
to|7294,7296
visit|7297,7302
her|7303,7306
again|7307,7312
on|7313,7315
_|7316,7317
_|7317,7318
_|7318,7319
for|7320,7323
re-evaluation|7324,7337
and|7338,7341
to|7342,7344
<EOL>|7345,7346
perform|7346,7353
stair|7354,7359
maneuvers|7360,7369
with|7370,7374
her|7375,7378
.|7378,7379
The|7380,7383
final|7384,7389
results|7390,7397
on|7398,7400
the|7401,7404
<EOL>|7405,7406
abcess|7406,7412
culture|7413,7420
was|7421,7424
streptococcus|7425,7438
Milleri|7439,7446
.|7446,7447
New|7448,7451
ID|7452,7454
recommendations|7455,7470
<EOL>|7471,7472
were|7472,7476
to|7477,7479
discontiniu|7480,7491
Vanco|7492,7497
and|7498,7501
Meropenum|7502,7511
,|7511,7512
she|7513,7516
was|7517,7520
started|7521,7528
on|7529,7531
<EOL>|7532,7533
Ceftriaxone|7533,7544
2|7545,7546
grams|7547,7552
and|7553,7556
and|7557,7560
Flagyl|7561,7567
Tid|7568,7571
.|7571,7572
<EOL>|7573,7574
<EOL>|7574,7575
On|7575,7577
_|7578,7579
_|7579,7580
_|7580,7581
,|7581,7582
patient|7583,7590
was|7591,7594
re-evaluated|7595,7607
by|7608,7610
_|7611,7612
_|7612,7613
_|7613,7614
and|7615,7618
OT|7619,7621
and|7622,7625
cleared|7626,7633
to|7634,7636
be|7637,7639
<EOL>|7640,7641
discharged|7641,7651
home|7652,7656
with|7657,7661
the|7662,7665
assistance|7666,7676
of|7677,7679
a|7680,7681
cane|7682,7686
.|7686,7687
They|7688,7692
also|7693,7697
<EOL>|7698,7699
recommend|7699,7708
services|7709,7717
while|7718,7723
patient|7724,7731
is|7732,7734
at|7735,7737
home|7738,7742
.|7742,7743
She|7744,7747
remained|7748,7756
stable|7757,7763
<EOL>|7764,7765
on|7765,7767
examination|7768,7779
.|7779,7780
<EOL>|7780,7781
<EOL>|7781,7782
On|7782,7784
_|7785,7786
_|7786,7787
_|7787,7788
,|7788,7789
Mrs.|7790,7794
_|7795,7796
_|7796,7797
_|7797,7798
was|7799,7802
seen|7803,7807
and|7808,7811
evaluated|7812,7821
,|7821,7822
she|7823,7826
<EOL>|7827,7828
complained|7828,7838
of|7839,7841
headache|7842,7850
and|7851,7854
a|7855,7856
non-contrast|7857,7869
head|7870,7874
CT|7875,7877
was|7878,7881
ordered|7882,7889
.|7889,7890
<EOL>|7891,7892
This|7892,7896
showed|7897,7903
the|7904,7907
stable|7908,7914
post-operative|7915,7929
changes|7930,7937
.|7937,7938
Home|7940,7944
services|7945,7953
<EOL>|7954,7955
were|7955,7959
established|7960,7971
and|7972,7975
the|7976,7979
patient|7980,7987
was|7988,7991
discharged|7992,8002
.|8002,8003
<EOL>|8003,8004
<EOL>|8004,8005
<EOL>|8006,8007
Medications|8007,8018
on|8019,8021
Admission|8022,8031
:|8031,8032
<EOL>|8032,8033
Ibuprofen|8033,8042
<EOL>|8042,8043
<EOL>|8044,8045
Discharge|8045,8054
Medications|8055,8066
:|8066,8067
<EOL>|8067,8068
1.|8068,8070
Acetaminophen|8071,8084
325|8085,8088
-|8088,8089
650|8089,8092
mg|8093,8095
PO|8096,8098
Q6H|8099,8102
:|8102,8103
PRN|8103,8106
pain|8107,8111
<EOL>|8112,8113
RX|8113,8115
*|8116,8117
acetaminophen|8117,8130
325|8131,8134
mg|8135,8137
_|8138,8139
_|8139,8140
_|8140,8141
tablet|8142,8148
(|8148,8149
s|8149,8150
)|8150,8151
by|8152,8154
mouth|8155,8160
every|8161,8166
six|8167,8170
(|8171,8172
6|8172,8173
)|8173,8174
<EOL>|8175,8176
hours|8176,8181
Disp|8182,8186
#|8187,8188
*|8188,8189
112|8189,8192
Tablet|8193,8199
Refills|8200,8207
:|8207,8208
*|8208,8209
0|8209,8210
<EOL>|8210,8211
2.|8211,8213
CeftriaXONE|8214,8225
2|8226,8227
gm|8228,8230
IV|8231,8233
Q12H|8234,8238
<EOL>|8239,8240
RX|8240,8242
*|8243,8244
ceftriaxone|8244,8255
2|8256,8257
gram|8258,8262
2|8263,8264
gm|8265,8267
IV|8268,8270
every|8271,8276
twelve|8277,8283
(|8284,8285
12|8285,8287
)|8287,8288
hours|8289,8294
Disp|8295,8299
#|8300,8301
*|8301,8302
84|8302,8304
<EOL>|8305,8306
Vial|8306,8310
Refills|8311,8318
:|8318,8319
*|8319,8320
0|8320,8321
<EOL>|8321,8322
3.|8322,8324
Docusate|8325,8333
Sodium|8334,8340
100|8341,8344
mg|8345,8347
PO|8348,8350
BID|8351,8354
<EOL>|8355,8356
RX|8356,8358
*|8359,8360
docusate|8360,8368
sodium|8369,8375
[|8376,8377
Colace|8377,8383
]|8383,8384
100|8385,8388
mg|8389,8391
1|8392,8393
capsule|8394,8401
(|8401,8402
s|8402,8403
)|8403,8404
by|8405,8407
mouth|8408,8413
twice|8414,8419
<EOL>|8420,8421
a|8421,8422
day|8423,8426
Disp|8427,8431
#|8432,8433
*|8433,8434
45|8434,8436
Capsule|8437,8444
Refills|8445,8452
:|8452,8453
*|8453,8454
0|8454,8455
<EOL>|8455,8456
4.|8456,8458
LeVETiracetam|8459,8472
1000|8473,8477
mg|8478,8480
PO|8481,8483
BID|8484,8487
<EOL>|8488,8489
RX|8489,8491
*|8492,8493
levetiracetam|8493,8506
[|8507,8508
Keppra|8508,8514
]|8514,8515
1,000|8516,8521
mg|8522,8524
1|8525,8526
tablet|8527,8533
(|8533,8534
s|8534,8535
)|8535,8536
by|8537,8539
mouth|8540,8545
twice|8546,8551
a|8552,8553
<EOL>|8554,8555
day|8555,8558
Disp|8559,8563
#|8564,8565
*|8565,8566
56|8566,8568
Tablet|8569,8575
Refills|8576,8583
:|8583,8584
*|8584,8585
0|8585,8586
<EOL>|8586,8587
5.|8587,8589
MetRONIDAZOLE|8590,8603
(|8604,8605
FLagyl|8605,8611
)|8611,8612
500|8613,8616
mg|8617,8619
PO|8620,8622
TID|8623,8626
<EOL>|8627,8628
RX|8628,8630
*|8631,8632
metronidazole|8632,8645
[|8646,8647
Flagyl|8647,8653
]|8653,8654
500|8655,8658
mg|8659,8661
1|8662,8663
tablet|8664,8670
(|8670,8671
s|8671,8672
)|8672,8673
by|8674,8676
mouth|8677,8682
three|8683,8688
<EOL>|8689,8690
times|8690,8695
a|8696,8697
day|8698,8701
Disp|8702,8706
#|8707,8708
*|8708,8709
126|8709,8712
Tablet|8713,8719
Refills|8720,8727
:|8727,8728
*|8728,8729
0|8729,8730
<EOL>|8730,8731
6.|8731,8733
OxycoDONE|8734,8743
(|8744,8745
Immediate|8745,8754
Release|8755,8762
)|8762,8763
5|8765,8766
mg|8767,8769
PO|8770,8772
Q6H|8773,8776
:|8776,8777
PRN|8777,8780
pain|8781,8785
<EOL>|8786,8787
RX|8787,8789
*|8790,8791
oxycodone|8791,8800
[|8801,8802
Oxecta|8802,8808
]|8808,8809
5|8810,8811
mg|8812,8814
1|8815,8816
tablet|8817,8823
,|8823,8824
oral|8825,8829
only|8830,8834
(|8834,8835
s|8835,8836
)|8836,8837
by|8838,8840
mouth|8841,8846
<EOL>|8847,8848
every|8848,8853
six|8854,8857
(|8858,8859
6|8859,8860
)|8860,8861
hours|8862,8867
Disp|8868,8872
#|8873,8874
*|8874,8875
168|8875,8878
Tablet|8879,8885
Refills|8886,8893
:|8893,8894
*|8894,8895
0|8895,8896
<EOL>|8896,8897
7.|8897,8899
Heparin|8900,8907
Flush|8908,8913
(|8914,8915
10|8915,8917
units|8918,8923
/|8923,8924
ml|8924,8926
)|8926,8927
2|8928,8929
mL|8930,8932
IV|8933,8935
DAILY|8936,8941
and|8942,8945
PRN|8946,8949
,|8949,8950
line|8951,8955
flush|8956,8961
<EOL>|8962,8963
<EOL>|8963,8964
RX|8964,8966
*|8967,8968
heparin|8968,8975
lock|8976,8980
flush|8981,8986
(|8987,8988
porcine|8988,8995
)|8995,8996
[|8997,8998
heparin|8998,9005
lock|9006,9010
flush|9011,9016
]|9016,9017
10|9018,9020
unit|9021,9025
/|9025,9026
mL|9026,9028
<EOL>|9029,9030
1|9030,9031
ml|9032,9034
IV|9035,9037
every|9038,9043
eight|9044,9049
(|9050,9051
8|9051,9052
)|9052,9053
hours|9054,9059
Disp|9060,9064
#|9065,9066
*|9066,9067
126|9067,9070
Vial|9071,9075
Refills|9076,9083
:|9083,9084
*|9084,9085
0|9085,9086
<EOL>|9086,9087
8.|9087,9089
Sodium|9090,9096
Chloride|9097,9105
0.9|9106,9109
%|9109,9110
Flush|9112,9117
10|9118,9120
mL|9121,9123
IV|9124,9126
Q8H|9127,9130
and|9131,9134
PRN|9135,9138
,|9138,9139
line|9140,9144
flush|9145,9150
<EOL>|9151,9152
Flush|9152,9157
before|9158,9164
and|9165,9168
after|9169,9174
each|9175,9179
infusion|9180,9188
of|9189,9191
antibiotics|9192,9203
.|9203,9204
<EOL>|9205,9206
RX|9206,9208
*|9209,9210
sodium|9210,9216
chloride|9217,9225
0.9|9226,9229
%|9230,9231
[|9232,9233
Normal|9233,9239
Saline|9240,9246
Flush|9247,9252
]|9252,9253
0.9|9254,9257
%|9258,9259
10|9260,9262
ml|9263,9265
IV|9266,9268
<EOL>|9269,9270
q12|9270,9273
Disp|9274,9278
#|9279,9280
*|9280,9281
168|9281,9284
Syringe|9285,9292
Refills|9293,9300
:|9300,9301
*|9301,9302
1|9302,9303
<EOL>|9303,9304
<EOL>|9304,9305
<EOL>|9306,9307
Discharge|9307,9316
Disposition|9317,9328
:|9328,9329
<EOL>|9329,9330
Home|9330,9334
With|9335,9339
Service|9340,9347
<EOL>|9347,9348
<EOL>|9349,9350
Facility|9350,9358
:|9358,9359
<EOL>|9359,9360
_|9360,9361
_|9361,9362
_|9362,9363
<EOL>|9363,9364
<EOL>|9365,9366
Discharge|9366,9375
Diagnosis|9376,9385
:|9385,9386
<EOL>|9386,9387
Brain|9387,9392
abscess|9393,9400
<EOL>|9400,9401
<EOL>|9401,9402
<EOL>|9403,9404
Discharge|9404,9413
Condition|9414,9423
:|9423,9424
<EOL>|9424,9425
Mental|9425,9431
Status|9432,9438
:|9438,9439
Clear|9440,9445
and|9446,9449
coherent|9450,9458
.|9458,9459
<EOL>|9459,9460
Level|9460,9465
of|9466,9468
Consciousness|9469,9482
:|9482,9483
Alert|9484,9489
and|9490,9493
interactive|9494,9505
.|9505,9506
<EOL>|9506,9507
Activity|9507,9515
Status|9516,9522
:|9522,9523
Ambulatory|9524,9534
-|9535,9536
requires|9537,9545
assistance|9546,9556
or|9557,9559
aid|9560,9563
(|9564,9565
walker|9565,9571
<EOL>|9572,9573
or|9573,9575
cane|9576,9580
)|9580,9581
.|9581,9582
<EOL>|9582,9583
<EOL>|9583,9584
<EOL>|9585,9586
Discharge|9586,9595
Instructions|9596,9608
:|9608,9609
<EOL>|9609,9610
|9610,9611
Have|9611,9615
a|9616,9617
friend|9618,9624
/|9624,9625
family|9625,9631
member|9632,9638
check|9639,9644
your|9645,9649
incision|9650,9658
daily|9659,9664
for|9665,9668
<EOL>|9669,9670
signs|9670,9675
of|9676,9678
infection|9679,9688
.|9688,9689
<EOL>|9689,9690
|9690,9691
Take|9691,9695
your|9696,9700
pain|9701,9705
medicine|9706,9714
as|9715,9717
prescribed|9718,9728
.|9728,9729
<EOL>|9729,9730
|9730,9731
Exercise|9731,9739
should|9740,9746
be|9747,9749
limited|9750,9757
to|9758,9760
walking|9761,9768
;|9768,9769
no|9770,9772
lifting|9773,9780
,|9780,9781
straining|9782,9791
,|9791,9792
<EOL>|9793,9794
or|9794,9796
excessive|9797,9806
bending|9807,9814
.|9814,9815
<EOL>|9815,9816
|9816,9817
*|9817,9818
*|9818,9819
Your|9819,9823
wound|9824,9829
was|9830,9833
closed|9834,9840
with|9841,9845
sutures|9846,9853
.|9853,9854
You|9855,9858
may|9859,9862
wash|9863,9867
your|9868,9872
hair|9873,9877
<EOL>|9878,9879
only|9879,9883
after|9884,9889
sutures|9890,9897
and|9898,9901
/|9901,9902
or|9902,9904
staples|9905,9912
have|9913,9917
been|9918,9922
removed|9923,9930
.|9930,9931
<EOL>|9932,9933
|9933,9934
You|9934,9937
may|9938,9941
shower|9942,9948
before|9949,9955
this|9956,9960
time|9961,9965
using|9966,9971
a|9972,9973
shower|9974,9980
cap|9981,9984
to|9985,9987
cover|9988,9993
<EOL>|9994,9995
your|9995,9999
head|10000,10004
.|10004,10005
<EOL>|10005,10006
|10006,10007
Increase|10007,10015
your|10016,10020
intake|10021,10027
of|10028,10030
fluids|10031,10037
and|10038,10041
fiber|10042,10047
,|10047,10048
as|10049,10051
narcotic|10052,10060
pain|10061,10065
<EOL>|10066,10067
medicine|10067,10075
can|10076,10079
cause|10080,10085
constipation|10086,10098
.|10098,10099
We|10100,10102
generally|10103,10112
recommend|10113,10122
taking|10123,10129
<EOL>|10130,10131
an|10131,10133
over|10134,10138
the|10139,10142
counter|10143,10150
stool|10151,10156
softener|10157,10165
,|10165,10166
such|10167,10171
as|10172,10174
Docusate|10175,10183
(|10184,10185
Colace|10185,10191
)|10191,10192
<EOL>|10193,10194
while|10194,10199
taking|10200,10206
narcotic|10207,10215
pain|10216,10220
medication|10221,10231
.|10231,10232
<EOL>|10232,10233
|10233,10234
Unless|10234,10240
directed|10241,10249
by|10250,10252
your|10253,10257
doctor|10258,10264
,|10264,10265
do|10266,10268
not|10269,10272
take|10273,10277
any|10278,10281
<EOL>|10282,10283
anti-inflammatory|10283,10300
medicines|10301,10310
such|10311,10315
as|10316,10318
Motrin|10319,10325
,|10325,10326
Aspirin|10327,10334
,|10334,10335
Advil|10336,10341
,|10341,10342
and|10343,10346
<EOL>|10347,10348
Ibuprofen|10348,10357
etc|10358,10361
.|10361,10362
<EOL>|10363,10364
|10364,10365
You|10365,10368
have|10369,10373
been|10374,10378
discharged|10379,10389
on|10390,10392
Keppra|10393,10399
(|10400,10401
Levetiracetam|10401,10414
)|10414,10415
,|10415,10416
you|10417,10420
will|10421,10425
<EOL>|10426,10427
not|10427,10430
require|10431,10438
blood|10439,10444
work|10445,10449
monitoring|10450,10460
.|10460,10461
<EOL>|10461,10462
|10462,10463
Clearance|10463,10472
to|10473,10475
drive|10476,10481
and|10482,10485
return|10486,10492
to|10493,10495
work|10496,10500
will|10501,10505
be|10506,10508
addressed|10509,10518
at|10519,10521
<EOL>|10522,10523
your|10523,10527
post-operative|10528,10542
office|10543,10549
visit|10550,10555
.|10555,10556
<EOL>|10556,10557
|10557,10558
Make|10558,10562
sure|10563,10567
to|10568,10570
continue|10571,10579
to|10580,10582
use|10583,10586
your|10587,10591
incentive|10592,10601
spirometer|10602,10612
while|10613,10618
<EOL>|10619,10620
at|10620,10622
home|10623,10627
,|10627,10628
unless|10629,10635
you|10636,10639
have|10640,10644
been|10645,10649
instructed|10650,10660
not|10661,10664
to|10665,10667
.|10667,10668
<EOL>|10669,10670
<EOL>|10670,10671
<EOL>|10672,10673
Followup|10673,10681
Instructions|10682,10694
:|10694,10695
<EOL>|10695,10696
_|10696,10697
_|10697,10698
_|10698,10699
<EOL>|10699,10700

