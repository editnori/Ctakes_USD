CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|true|false||Unit
null|Unit device|Device|true|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|true|false||Unit
null|Unit of Measure|LabModifier|true|false||Unit
null|Unit|LabModifier|true|false||Unit
null|Enzyme Unit|LabModifier|true|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|codeine|Drug|false|false||Codeine
null|codeine|Drug|false|false||Codeinenull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|null|Finding|false|false||Dyspnea
null|Dyspnea|Finding|false|false||Dyspneanull|Melena|Finding|false|false||melenanull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Tumor stage|Attribute|false|false||stagenull|Stage|Time|false|false||stage
null|Phase|Time|false|false||stagenull|CELP gene|Finding|false|false||cell
null|CEL gene|Finding|false|false||cellnull|Cells|Anatomy|false|false||cellnull|Cell Device|Device|false|false||cell
null|Cellular Phone|Device|false|false||cellnull|Cell (compartment)|Modifier|false|false||cellnull|Malignant neoplasm of lung|Disorder|false|false||lung cancer
null|Carcinoma of lung|Disorder|false|false||lung cancernull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Chronic Kidney Diseases|Disorder|false|false||CKDnull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|Productive Cough|Finding|false|false||productive coughnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Melena|Finding|false|false||melenanull|Has patient|Finding|false|false||Patient hasnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|day|Time|true|false||daysnull|Melena|Finding|true|false||melenanull|Abdominal Pain|Finding|true|false||abdominal painnull|Abdomen|Anatomy|true|false||abdominalnull|Abdominal (qualifier value)|Modifier|true|false||abdominalnull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|null|Finding|true|false||dyspnea
null|Dyspnea|Finding|true|false||dyspneanull|Patient Outcome - Worsening|Finding|true|false||worseningnull|Worsening (qualifier value)|Modifier|true|false||worseningnull|Cough (guaifenesin)|Drug|true|false||cough
null|Cough (guaifenesin)|Drug|true|false||coughnull|Coughing|Finding|true|false||coughnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Fever|Finding|true|false||feversnull|Chest Pain|Finding|true|false||chest painnull|null|Attribute|true|false||chest painnull|Chest problem|Finding|true|false||chestnull|Chest|Anatomy|true|false||chest
null|Anterior thoracic region|Anatomy|true|false||chestnull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Initial (abbreviation)|Finding|false|false||initialnull|Initially|Time|false|false||initialnull|Firstly|Modifier|false|false||initialnull|Hemopoietic stem cell transplant|Procedure|false|false||hct
null|Hematocrit Measurement|Procedure|false|false||hctnull|Recent|Time|false|false||recentnull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|null|Finding|false|false||transfusionnull|Transfusion (procedure)|Procedure|false|false||transfusion
null|Blood Transfusion|Procedure|false|false||transfusionnull|dependent|Finding|false|false||dependentnull|Dependent - ability|Modifier|false|false||dependent
null|Conditional|Modifier|false|false||dependentnull|Anemia|Disorder|false|false||anemianull|Anemia <Anemiaceae>|Entity|false|false||anemianull|Initially|Time|false|false||initiallynull|Hypoxia|Finding|false|false||hypoxicnull|A1BG gene|Finding|false|false||ABGnull|Analysis of arterial blood gases and pH|Procedure|false|false||ABGnull|lactate|Drug|false|false||lactate
null|lactate|Drug|false|false||lactate
null|Lactates|Drug|false|false||lactatenull|Lactic acid measurement|Procedure|false|false||lactatenull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Nebulizer solution|Drug|false|false||nebsnull|Stress bismuth subsalicylate|Drug|false|false||stress
null|Stress bismuth subsalicylate|Drug|false|false||stressnull|Stress|Finding|false|false||stressnull|W stress|Attribute|false|false||stressnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Steroids|Drug|false|false||steroids
null|Steroids|Drug|false|false||steroidsnull|Levaquin|Drug|false|false||levaquin
null|Levaquin|Drug|false|false||levaquinnull|ceftriaxone|Drug|false|false||ceftriaxone
null|ceftriaxone|Drug|false|false||ceftriaxonenull|Improvement|Finding|false|false||improvementnull|short-acting thyroid stimulator|Drug|false|false||sats
null|short-acting thyroid stimulator|Drug|false|false||satsnull|Middle|Modifier|false|false||midnull|On IV|Finding|false|false||on IVnull|Proton Pump Inhibitors|Drug|false|false||PPInull|Prepulse Inhibition|Finding|false|false||PPInull|guaiac positive|Lab|false|false||guaiac positivenull|guaiac|Drug|false|false||guaiac
null|guaiac|Drug|false|false||guaiacnull|BRAF Gene Rearrangement|Disorder|false|false||positivenull|Rh Positive Blood Group|Finding|false|false||positive
null|Positive Finding|Finding|false|false||positive
null|Positive|Finding|false|false||positivenull|Positive Charge|Modifier|false|false||positivenull|Positive Number|LabModifier|false|false||positivenull|Dark Brown|Modifier|false|false||dark brownnull|Dark color|Modifier|false|false||darknull|Brown color of stool|Finding|false|false||brown stoolnull|Brown Tendon Sheath Syndrome|Disorder|false|false||brownnull|Brown color|Modifier|false|false||brownnull|Feces|Finding|false|false||stoolnull|Stool seat|Device|false|false||stoolnull|Plain chest X-ray|Procedure|false|false||CXRnull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|Pleural Diseases|Disorder|false|false||pleuralnull|Pleura|Anatomy|false|false||pleuralnull|Pleural|Modifier|false|false||pleuralnull|Effusion (substance)|Finding|false|false||effusion
null|null|Finding|false|false||effusion
null|effusion|Finding|false|false||effusionnull|Equivocal|Modifier|false|false||questionablenull|Structure of lower lobe of lung|Anatomy|false|false||lower lobenull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|AKT1S1 wt Allele|Finding|false|false||lobe
null|AKT1S1 gene|Finding|false|false||lobenull|lobe|Anatomy|false|false||lobenull|Collapse (finding)|Finding|false|false||collapse
null|Shock|Finding|false|false||collapse
null|null|Finding|false|false||collapsenull|Collapse (morphologic abnormality)|Phenomenon|false|false||collapsenull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|Sinus Tachycardia|Disorder|false|false||sinus tachnull|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false||sinus
null|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false||sinusnull|pathologic fistula|Disorder|false|false||sinusnull|Sinus - general anatomical term|Anatomy|false|false||sinus
null|Nasal sinus|Anatomy|false|false||sinusnull|Mental Depression|Disorder|false|false||depressionsnull|Transfer - product ownership|Finding|false|false||transfer
null|Transfer Technique|Finding|false|false||transfer
null|ActClass - transfer|Finding|false|false||transfer
null|null|Finding|false|false||transfernull|Transfer (immobility management)|Procedure|false|false||transfernull|Psychological Well Being|Finding|false|false||feeling betternull|Observation Interpretation - better|Finding|false|false||betternull|Better|Modifier|false|false||betternull|outcomes otolaryngology breathing|Finding|false|false||breathing
null|Inspiration (function)|Finding|false|false||breathing
null|Respiration|Finding|false|false||breathingnull|null|Attribute|false|false||breathingnull|respiratory system process|Phenomenon|false|false||breathingnull|Therapeutic procedure|Procedure|false|false||treatmentsnull|Has difficulty doing (qualifier value)|Finding|false|false||difficultynull|ErbB Receptors|Drug|false|false||her family
null|ErbB Receptors|Drug|false|false||her familynull|ErbB Receptors|Finding|false|false||her familynull|Entity Name Part Type - family|Finding|false|false||family
null|Last Name|Finding|false|false||family
null|Living Arrangement - Family|Finding|false|false||family
null|Family (taxonomic)|Finding|false|false||family
null|Family Collection|Finding|false|false||familynull|Family|Subject|false|false||familynull|hearing impairment|Disorder|false|true||difficulty hearingnull|Partial Hearing Loss|Finding|false|true||difficulty hearingnull|Has difficulty doing (qualifier value)|Finding|false|false||difficultynull|outcomes otolaryngology hearing|Finding|false|false||hearing
null|Hearing finding|Finding|false|false||hearing
null|Hearing|Finding|false|false||hearingnull|Amnesia|Disorder|true|false||memory lossnull|Memory Loss|Finding|true|false||memory lossnull|Memory observations|Finding|true|false||memory
null|Memory G-code|Finding|true|false||memory
null|Memory|Finding|true|false||memorynull|Memory Device|Device|true|false||memorynull|Loss (adaptation)|Finding|true|false||lossnull|Loss (quantitative)|LabModifier|true|false||lossnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Intermittent|Time|false|false||intermittentnull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|week|Time|false|false||weeksnull|null|Drug|false|false||codeine syrupnull|codeine|Drug|false|false||codeine
null|codeine|Drug|false|false||codeinenull|Syrup Drug Form|Drug|false|false||syrup
null|Syrup (dietary)|Drug|false|false||syrupnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Menstruation|Finding|false|false||periodnull|Clinical Trial Period|Procedure|false|false||periodnull|per period (qualifier value)|Time|false|false||period
null|Time periods|Time|false|false||periodnull|Transaction counts and value totals - Period|LabModifier|false|false||periodnull|Improvement|Finding|false|false||improvementnull|Cough (guaifenesin)|Drug|true|false||cough
null|Cough (guaifenesin)|Drug|true|false||coughnull|Coughing|Finding|true|false||coughnull|Fever|Finding|true|false||feversnull|Chills|Finding|true|false||chillsnull|Chest Pain|Finding|true|false||chest painnull|null|Attribute|true|false||chest painnull|Chest problem|Finding|true|false||chestnull|Chest|Anatomy|true|false||chest
null|Anterior thoracic region|Anatomy|true|false||chestnull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|null|Time|true|false||priornull|History of present illness (finding)|Finding|true|false||history
null|History of previous events|Finding|true|false||history
null|Historical aspects qualifier|Finding|true|false||history
null|Medical History|Finding|true|false||history
null|Concept History|Finding|true|false||historynull|History|Subject|true|false||historynull|Melena|Finding|true|false||melenanull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Poor appetite question|Finding|false|false||poor appetite
null|Decrease in appetite|Finding|false|false||poor appetitenull|null|Attribute|false|false||poor appetitenull|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group|Finding|false|false||poor
null|Patient Condition Code - Poor|Finding|false|false||poornull|Poverty|Subject|false|false||poornull|Language Proficiency - Poor|Modifier|false|false||poor
null|Specimen Quality - Poor|Modifier|false|false||poor
null|Poor - grade|Modifier|false|false||poor
null|Poor - qualifier|Modifier|false|false||poornull|Desire for food|Finding|false|false||appetitenull|month|Time|false|false||monthsnull|Gastroesophageal reflux disease|Disorder|true|false||heartburnnull|Heartburn|Finding|true|false||heartburnnull|Deglutition Disorders|Disorder|true|false||dysphagianull|Metastatic non-small cell lung cancer|Disorder|false|false||Stage IV nonsmall cell lung cancernull|Stage level 4|Finding|false|false||Stage IVnull|Tumor stage|Attribute|false|false||Stagenull|Stage|Time|false|false||Stage
null|Phase|Time|false|false||Stagenull|CELP gene|Finding|false|false||cell
null|CEL gene|Finding|false|false||cellnull|Cells|Anatomy|false|false||cellnull|Cell Device|Device|false|false||cell
null|Cellular Phone|Device|false|false||cellnull|Cell (compartment)|Modifier|false|false||cellnull|Adenocarcinoma of lung (disorder)|Disorder|false|false||lung cancer, adenocarcinomanull|Malignant neoplasm of lung|Disorder|false|false||lung cancer
null|Carcinoma of lung|Disorder|false|false||lung cancernull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Adenocarcinoma|Disorder|false|false||adenocarcinoma
null|Malignant adenomatous neoplasm|Disorder|false|false||adenocarcinomanull|EGFR protein, human|Drug|false|false||EGFR
null|Epidermal Growth Factor Receptor|Drug|false|false||EGFR
null|Epidermal Growth Factor Receptor|Drug|false|false||EGFR
null|Soluble ErbB-1|Drug|false|false||EGFRnull|EGFR protein, human|Finding|false|false||EGFR
null|Epidermal Growth Factor Receptor|Finding|false|false||EGFR
null|epidermal growth factor receptor activity|Finding|false|false||EGFR
null|Soluble ErbB-1|Finding|false|false||EGFR
null|EGFR gene|Finding|false|false||EGFRnull|Estimated Glomerular Filtration Rate|Procedure|false|false||EGFRnull|Type - ParameterizedDataType|Finding|false|false||type
null|SGCG gene|Finding|false|false||typenull|null|Modifier|false|false||typenull|KRAS protein, human|Drug|false|false||KRAS
null|KRAS protein, human|Drug|false|false||KRASnull|KRAS gene|Finding|false|false||KRAS
null|K-ras Oncogene|Finding|false|false||KRAS
null|Human Oncogene K-Ras|Finding|false|false||KRASnull|Mutation Abnormality|Disorder|false|false||mutatednull|Gene Variant Positive|Lab|false|false||mutatednull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Coronary Artery Bypass Surgery|Procedure|false|false||CABGnull|SERPINA5 protein, human|Drug|false|false||PCI
null|SERPINA5 protein, human|Drug|false|false||PCInull|Peritoneal Cancer Index|Finding|false|false||PCI
null|SERPINA5 wt Allele|Finding|false|false||PCI
null|SERPINA5 gene|Finding|false|false||PCInull|Percutaneous Coronary Intervention|Procedure|false|false||PCI
null|photochemical internalization|Procedure|false|false||PCI
null|Prophylactic Cranial Irradiation|Procedure|false|false||PCInull|Picocurie|LabModifier|false|false||PCInull|Leukocyte adhesion deficiency type 1|Disorder|false|false||LAD
null|Leukocyte adhesion deficiency|Disorder|false|false||LADnull|ITGB2 wt Allele|Finding|false|false||LAD
null|DLD gene|Finding|false|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false||LADnull|Ladino Language|Entity|false|false||LADnull|Chronic Kidney Insufficiency|Disorder|false|false||Chronic renal insufficiencynull|Chronic - Admission Level of Care Code|Finding|false|false||Chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||Chronicnull|chronic|Time|false|false||Chronicnull|Renal Insufficiency|Disorder|false|false||renal insufficiency
null|Kidney Failure|Disorder|false|false||renal insufficiencynull|Urologic Diseases|Disorder|false|false||renalnull|Kidney|Anatomy|false|false||renalnull|Insufficiency|Finding|false|false||insufficiencynull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|With glomerular filtration rate|Modifier|false|false||with GFRnull|RAPGEF5 gene|Finding|false|false||GFRnull|Glomerular Filtration Rate|LabModifier|false|false||GFRnull|Cyclophosphamide/Doxorubicin/Vincristine|Drug|false|false||CVAnull|Acute ill-defined cerebrovascular disease|Disorder|false|false||CVA
null|Cerebrovascular accident|Disorder|false|false||CVAnull|Small|LabModifier|false|false||smallnull|Left posterior|Modifier|false|false||left posteriornull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Posterior pituitary disease|Disorder|false|false||posteriornull|Dorsal|Modifier|false|false||posteriornull|Coronal (qualifier value)|Modifier|false|false||frontalnull|Infarction|Finding|false|false||infarctnull|Hypercholesterolemia|Disorder|false|false||Hypercholesterolemianull|Hypercholesterolemia result|Finding|false|false||Hypercholesterolemianull|Age related macular degeneration|Disorder|false|false||Macular Degeneration
null|Macular degeneration|Disorder|false|false||Macular Degenerationnull|macular|Modifier|false|false||Macularnull|biologic degeneration|Finding|false|false||Degeneration
null|Abnormal degeneration|Finding|false|false||Degenerationnull|Indirect exposure mechanism - Father|Finding|false|false||father
null|Relationship - Father|Finding|false|false||father
null|Father - courtesy title|Finding|false|false||fathernull|Father (person)|Subject|false|false||fathernull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|Relationship - Mother|Finding|false|false||mothernull|Mother (person)|Subject|false|false||mothernull|Neoplasm of uncertain or unknown behavior of stomach|Disorder|false|false||stomach
null|Stomach Diseases|Disorder|false|false||stomach
null|Benign neoplasm of stomach|Disorder|false|false||stomach
null|Carcinoma in situ of stomach|Disorder|false|false||stomachnull|Stomach problem|Finding|false|false||stomachnull|Procedure on stomach|Procedure|false|false||stomachnull|Stomach structure|Anatomy|false|false||stomach
null|Abdomen>Stomach|Anatomy|false|false||stomach
null|Stomach|Anatomy|false|false||stomachnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Osteosarcoma of bone|Disorder|false|false||osteosarcoma
null|Osteosarcoma|Disorder|false|false||osteosarcomanull|RB1 gene|Finding|false|false||osteosarcomanull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Generalnull|General medical service|Procedure|false|false||Generalnull|Generalized|Modifier|false|false||Generalnull|Elderly (population group)|Subject|false|false||Elderlynull|Old age|Time|false|false||Elderlynull|Chronically Ill|Disorder|false|false||chronically illnull|Patient appears chronically ill|Finding|false|false||chronically illnull|Malaise|Finding|false|false||illnull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|HEENT|Anatomy|false|false||HEENTnull|Scleral Diseases|Disorder|false|false||scleranull|examination of sclera|Procedure|false|false||scleranull|Sclera|Anatomy|false|false||scleranull|Anicteric|Finding|false|false||anictericnull|Myelofibrosis|Disorder|false|false||MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false||MMMnull|Passive joint movement of neck (finding)|Finding|false|false||Neck
null|Neck problem|Finding|false|false||Necknull|dendritic spine neck|Anatomy|false|false||Neck
null|Neck|Anatomy|false|false||Necknull|Supple|Finding|true|false||supplenull|Jugular venous pressure|Finding|true|false||JVPnull|Firm|Modifier|true|false||firmnull|Bilateral|Modifier|true|false||bilateralnull|Submandibular|Modifier|true|false||submandibularnull|Leukocyte adhesion deficiency type 1|Disorder|false|false||LAD
null|Leukocyte adhesion deficiency|Disorder|false|false||LADnull|ITGB2 wt Allele|Finding|false|false||LAD
null|DLD gene|Finding|false|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false||LADnull|Ladino Language|Entity|false|false||LADnull|Lung|Anatomy|false|false||Lungsnull|Dental Percussion|Procedure|false|false||percussion
null|Percussion|Procedure|false|false||percussionnull|Right lung|Anatomy|false|false||right lungnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|null|Attribute|false|false||breath sounds
null|Respiratory Sounds|Attribute|false|false||breath soundsnull|Breath|Finding|false|false||breathnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|Basilar Rales|Finding|false|false||crackles
null|Rales|Finding|false|false||cracklesnull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|lobe|Anatomy|false|false||lobesnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Wheezing|Finding|false|false||wheezingnull|Regular|Modifier|false|false||Regularnull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Rhythm|Finding|true|false||rhythm
null|rhythmic process (biological)|Finding|true|false||rhythmnull|Heart murmur|Finding|true|false||murmursnull|Pericardial friction rub|Finding|true|false||rubsnull|Malignant neoplasm of abdomen|Disorder|false|false||Abdomennull|Abdomen problem|Finding|false|false||Abdomennull|Abdomen|Anatomy|false|false||Abdomen
null|Abdominal Cavity|Anatomy|false|false||Abdomennull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|Bowel sounds|Finding|true|false||bowel soundsnull|Intestines|Anatomy|true|false||bowelnull|null|Device|true|false||soundsnull|null|Phenomenon|true|false||soundsnull|Present|Finding|true|false||present
null|Presentation|Finding|true|false||presentnull|Rebound tenderness|Finding|true|false||rebound tendernessnull|Emotional tenderness|Finding|true|false||tenderness
null|Sore to touch|Finding|true|false||tendernessnull|Protective muscle spasm|Finding|true|false||guardingnull|Organomegaly|Finding|true|false||organomegalynull|Hereditary Multiple Exostoses|Disorder|true|false||Extnull|EXT1 wt Allele|Finding|true|false||Ext
null|EXT1 gene|Finding|true|false||Extnull|Feels warm|Finding|false|false||warmnull|warming process|Phenomenon|false|false||warmnull|Well (answer to question)|Finding|true|false||wellnull|Well (container)|Device|true|false||wellnull|Microplate Well|Modifier|true|false||well
null|Good|Modifier|true|false||well
null|Healthy|Modifier|true|false||wellnull|null|Drug|true|false||pulsesnull|Physiologic pulse|Finding|true|false||pulsesnull|Pulse taking|Procedure|true|false||pulsesnull|Clubbing|Disorder|true|false||clubbingnull|Cyanosis|Finding|true|false||cyanosisnull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Certificate Status - Expired|Finding|false|false||expired
null|Referral status - Expired|Finding|false|false||expired
null|Cessation of life|Finding|false|false||expired
null|Expiration, Respiratory|Finding|false|false||expired
null|Expiration|Finding|false|false||expirednull|Specimen Reject Reason - Expired|Modifier|false|false||expirednull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Lymph|Finding|false|false||Lymphsnull|Monos|Drug|false|false||Monos
null|Mono-S|Drug|false|false||Monos
null|Monos|Drug|false|false||Monosnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||Eos
null|Familial eosinophilia|Disorder|false|false||Eosnull|PRSS33 gene|Finding|false|false||Eos
null|IKZF4 gene|Finding|false|false||Eosnull|Eos <Loriini>|Entity|false|false||Eosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||ASTnull|Atypical Spitz Nevus|Disorder|false|false||ASTnull|SLC17A5 wt Allele|Finding|false|false||AST
null|SLC17A5 gene|Finding|false|false||AST
null|GOT1 gene|Finding|false|false||ASTnull|Asterion|Anatomy|false|false||ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Lactate Dehydrogenase|Drug|false|false||LDH
null|Lactate Dehydrogenase|Drug|false|false||LDHnull|Lifetime Drinking History|Finding|false|false||LDHnull|Lactate dehydrogenase measurement|Procedure|false|false||LDHnull|Creatine Kinase|Drug|false|false||CPK
null|Creatine Kinase|Drug|false|false||CPKnull|PIK3C2A gene|Finding|false|false||CPKnull|Creatine kinase measurement|Procedure|false|false||CPKnull|Alkaline Phosphatase|Drug|false|false||AlkPhos
null|Alkaline Phosphatase|Drug|false|false||AlkPhosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MB
null|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MBnull|creatine kinase activity|Finding|false|false||CK-MBnull|Serum creatine phosphokinase MB isoenzyme measurement|Procedure|false|false||CK-MB
null|Creatine kinase MB measurement|Procedure|false|false||CK-MBnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MB
null|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MBnull|creatine kinase activity|Finding|false|false||CK-MBnull|Serum creatine phosphokinase MB isoenzyme measurement|Procedure|false|false||CK-MB
null|Creatine kinase MB measurement|Procedure|false|false||CK-MBnull|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Partial pressure of Oxygen|Finding|false|false||pO2
null|US Military enlisted E5|Finding|false|false||pO2null|PO2 measurement|Procedure|false|false||pO2null|Carbon dioxide measurement, partial pressure|Procedure|false|false||pCO2null|Carbon dioxide, partial pressure|Lab|false|false||pCO2null|nitrogenous base|Drug|false|false||Base
null|Base|Drug|false|false||Base
null|Dental Base|Drug|false|false||Base
null|base - RoleClass|Drug|false|false||Basenull|Base - General Qualifier|Finding|false|false||Base
null|BPIFA4P gene|Finding|false|false||Base
null|Base - RX Component Type|Finding|false|false||Basenull|Anatomical base|Anatomy|false|false||Basenull|Base - unit of product usage|LabModifier|false|false||Basenull|Published Comment|Finding|false|false||Comment
null|Comment|Finding|false|false||Commentnull|Green color|Modifier|false|false||GREENnull|Encounter due to blood type|Finding|false|false||BLOOD Type
null|Blood Group Systems|Finding|false|false||BLOOD Typenull|Blood group typing (procedure)|Procedure|false|false||BLOOD Typenull|Blood Type|Attribute|false|false||BLOOD Typenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Type - ParameterizedDataType|Finding|false|false||Type
null|SGCG gene|Finding|false|false||Typenull|null|Modifier|false|false||Typenull|artesunate|Drug|false|false||ART
null|artesunate|Drug|false|false||ARTnull|AGRP wt Allele|Finding|false|false||ART
null|AGRP gene|Finding|false|false||ARTnull|Assisted Reproductive Technologies|Procedure|false|false||ART
null|Antiretroviral therapy|Procedure|false|false||ARTnull|Artwork|Device|false|false||ARTnull|Arts|Subject|false|false||ARTnull|Partial pressure of Oxygen|Finding|false|false||pO2
null|US Military enlisted E5|Finding|false|false||pO2null|PO2 measurement|Procedure|false|false||pO2null|Carbon dioxide measurement, partial pressure|Procedure|false|false||pCO2null|Carbon dioxide, partial pressure|Lab|false|false||pCO2null|nitrogenous base|Drug|false|false||Base
null|Base|Drug|false|false||Base
null|Dental Base|Drug|false|false||Base
null|base - RoleClass|Drug|false|false||Basenull|Base - General Qualifier|Finding|false|false||Base
null|BPIFA4P gene|Finding|false|false||Base
null|Base - RX Component Type|Finding|false|false||Basenull|Anatomical base|Anatomy|false|false||Basenull|Base - unit of product usage|LabModifier|false|false||Basenull|lactate in blood (lab test)|Procedure|false|false||BLOOD Lactatenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|lactate|Drug|false|false||Lactate
null|lactate|Drug|false|false||Lactate
null|Lactates|Drug|false|false||Lactatenull|Lactic acid measurement|Procedure|false|false||Lactatenull|lactate in blood (lab test)|Procedure|false|false||BLOOD Lactatenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|lactate|Drug|false|false||Lactate
null|lactate|Drug|false|false||Lactate
null|Lactates|Drug|false|false||Lactatenull|Lactic acid measurement|Procedure|false|false||Lactatenull|lactate in blood (lab test)|Procedure|false|false||BLOOD Lactatenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|lactate|Drug|false|false||Lactate
null|lactate|Drug|false|false||Lactate
null|Lactates|Drug|false|false||Lactatenull|Lactic acid measurement|Procedure|false|false||Lactatenull|lactate in blood (lab test)|Procedure|false|false||BLOOD Lactatenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|lactate|Drug|false|false||Lactate
null|lactate|Drug|false|false||Lactate
null|Lactates|Drug|false|false||Lactatenull|Lactic acid measurement|Procedure|false|false||Lactatenull|Color of urine|Finding|false|false||URINE Colornull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|color additive|Drug|false|false||Color
null|Coloring Excipient|Drug|false|false||Colornull|color - solid dosage form|Modifier|false|false||Color
null|Color|Modifier|false|false||Colornull|Color quantity|LabModifier|false|false||Colornull|Cereal plant straw|Drug|false|false||Strawnull|Straw package type|Device|false|false||Strawnull|Straw Color|Modifier|false|false||Strawnull|Straw (unit of presentation)|LabModifier|false|false||Strawnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Hematuria|Disorder|false|false||URINE Bloodnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Blood and lymphatic system disorders|Disorder|false|false||Bloodnull|peripheral blood|Finding|false|false||Blood
null|Blood|Finding|false|false||Blood
null|In Blood|Finding|false|false||Bloodnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|nitrite ion|Drug|false|false||Nitrite
null|Nitrites|Drug|false|false||Nitrite
null|Nitrites|Drug|false|false||Nitrite
null|Nitrites|Drug|false|false||Nitrite
null|nitrite ion|Drug|false|false||Nitrite
null|nitrite ion|Drug|false|false||Nitritenull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Proteins|Drug|false|false||Protein
null|Proteins|Drug|false|false||Proteinnull|Protein Info|Finding|false|false||Proteinnull|Protein measurement|Procedure|false|false||Proteinnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Ketones|Drug|false|false||Ketonenull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|null|Lab|false|false||URINE RBC
null|Red blood cells urine positive|Lab|false|false||URINE RBCnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Leukocytes|Anatomy|true|false||WBCnull|Yeast, Dried|Drug|true|false||Yeast
null|Candida albicans allergenic extract|Drug|true|false||Yeast
null|Candida albicans allergenic extract|Drug|true|false||Yeast
null|Candida albicans allergenic extract|Drug|true|false||Yeastnull|Saccharomyces cerevisiae|Entity|true|false||Yeast
null|Yeasts|Entity|true|false||Yeastnull|Tissue Factor Pathway Inhibitor, human|Drug|true|false||Epi
null|epinephrine|Drug|true|false||Epi
null|epinephrine|Drug|true|false||Epi
null|epinephrine|Drug|true|false||Epi
null|Tissue Factor Pathway Inhibitor, human|Drug|true|false||Epinull|Exocrine pancreatic insufficiency|Disorder|true|false||Epinull|Eysenck personality inventory|Finding|true|false||Epi
null|TFPI wt Allele|Finding|true|false||Epi
null|TFPI gene|Finding|true|false||Epinull|Electronic Portal Imaging|Procedure|true|false||Epi
null|Echo-Planar Imaging|Procedure|true|false||Epinull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Hour|Time|false|false||Hoursnull|Random|Modifier|false|false||RANDOMnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Parameterized Data Type - Interval|Finding|false|false||Intervalnull|Interval|Time|false|false||Intervalnull|Enlargement (morphologic abnormality)|Disorder|false|false||enlargementnull|Hypertrophy|Finding|false|false||enlargementnull|Enlargement procedure|Procedure|false|false||enlargementnull|Massive|Modifier|false|false||massivenull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Pleural Diseases|Disorder|false|false||pleuralnull|Pleura|Anatomy|false|false||pleuralnull|Pleural|Modifier|false|false||pleuralnull|Effusion (substance)|Finding|false|false||effusion
null|null|Finding|false|false||effusion
null|effusion|Finding|false|false||effusionnull|Greater|LabModifier|false|false||larger
null|Large|LabModifier|false|false||largernull|Lung consolidation|Disorder|false|false||consolidationnull|Consolidation|Modifier|false|false||consolidationnull|Left lung|Anatomy|false|false||left lungnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|Possible|Finding|false|false||possiblynull|Possible diagnosis|Modifier|false|false||possiblynull|Extent|Modifier|false|false||extension ofnull|Telephone Extension Number|Finding|false|false||extension
null|Extension|Finding|false|false||extensionnull|Neoplasms|Disorder|false|false||tumornull|Tumor Mass|Finding|false|false||tumor
null|null|Finding|false|false||tumornull|Focal|Modifier|false|false||focalnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Administration Method - Infiltrate|Finding|false|false||infiltrate
null|null|Finding|false|false||infiltrate
null|Infiltration|Finding|false|false||infiltratenull|combination - answer to question|Finding|false|false||combinationnull|combination of objects|Entity|false|false||combinationnull|Combined|Modifier|false|false||combinationnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Biphasic Continuous Positive Airway Pressure|Procedure|false|false||BiPAPnull|Comfort brand of hydroxyethyl cellulose|Drug|false|false||comfort
null|Comfort brand of hydroxyethyl cellulose|Drug|false|false||comfortnull|Comfort|Finding|false|false||comfortnull|Oncologists|Subject|false|false||oncologistnull|Overnight|Time|false|false||overnightnull|Thoracentesis|Procedure|false|false||thoracentesisnull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Volume (publication)|Finding|false|false||volumenull|Volume|LabModifier|false|false||volumenull|Encounter due to palliative care|Finding|false|false||Palliative carenull|Palliative Care|Procedure|false|false||Palliative care
null|Palliative Nursing|Procedure|false|false||Palliative carenull|Palliative care service|Entity|false|false||Palliativenull|Palliative|Modifier|false|false||Palliativenull|Continuity Assessment Record and Evaluation|Finding|false|false||care
null|In care (finding)|Finding|false|false||carenull|care activity|Event|false|false||carenull|Decision|Finding|false|false||decisionnull|Has focus|Finding|false|false||focusnull|Focal|Modifier|false|false||focusnull|Comfort brand of hydroxyethyl cellulose|Drug|false|false||comfort
null|Comfort brand of hydroxyethyl cellulose|Drug|false|false||comfortnull|Comfort|Finding|false|false||comfortnull|Oncologists|Subject|false|false||oncologistnull|ErbB Receptors|Drug|false|false||her family
null|ErbB Receptors|Drug|false|false||her familynull|ErbB Receptors|Finding|false|false||her familynull|Entity Name Part Type - family|Finding|false|false||family
null|Last Name|Finding|false|false||family
null|Living Arrangement - Family|Finding|false|false||family
null|Family (taxonomic)|Finding|false|false||family
null|Family Collection|Finding|false|false||familynull|Family|Subject|false|false||familynull|Inventory of Callous-Unemotional Traits|Finding|false|false||ICUnull|Structure of intraculminate fissure|Anatomy|false|false||ICUnull|intensive care unit|Device|false|false||ICUnull|intensive care unit|Entity|false|false||ICUnull|Floor (anatomic)|Anatomy|false|false||floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Then|Time|false|false||soon afternull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|Robitussin|Drug|false|false||Robitussin
null|Robitussin|Drug|false|false||Robitussinnull|codeine|Drug|false|false||codeine
null|codeine|Drug|false|false||codeinenull|thrombospondin-1, human|Drug|false|false||tsp
null|Thrombospondins|Drug|false|false||tsp
null|Thrombospondins|Drug|false|false||tspnull|Tropical Spastic Paraparesis|Disorder|false|false||tspnull|THBS1 wt Allele|Finding|false|false||tsp
null|THBS1 gene|Finding|false|false||tspnull|Teaspoon Dosing Unit|LabModifier|false|false||tsp
null|Teaspoonful|LabModifier|false|false||tspnull|Once a day, at bedtime|Time|false|false||QHSnull|atorvastatin|Drug|false|false||ATORVASTATIN
null|atorvastatin|Drug|false|false||ATORVASTATINnull|Lipitor|Drug|false|false||LIPITOR
null|Lipitor|Drug|false|false||LIPITORnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Oral Route of Administration|Finding|true|false||by mouthnull|Oral cavity|Anatomy|true|false||mouth
null|Oral region|Anatomy|true|false||mouthnull|One Daily|Drug|true|false||one daily
null|One Daily|Drug|true|false||one daily
null|One Daily|Drug|true|false||one dailynull|Daily|Time|true|false||dailynull|Substitution - ActClass|Finding|true|false||Substitutionnull|Substitution - change|Event|true|false||Substitutionnull|benzonatate|Drug|true|false||BENZONATATE
null|benzonatate|Drug|true|false||BENZONATATEnull|capsule (pharmacologic)|Drug|true|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|true|false||Capsule
null|Structure of organ capsule|Anatomy|true|false||Capsulenull|Capsule Shape|Modifier|true|false||Capsulenull|Capsule (unit of presentation)|LabModifier|true|false||Capsule
null|Capsule Dosing Unit|LabModifier|true|false||Capsulenull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Thrice|LabModifier|false|false||three timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Calcitriol Drug Class|Drug|false|false||CALCITRIOL
null|calcitriol|Drug|false|false||CALCITRIOL
null|calcitriol|Drug|false|false||CALCITRIOL
null|calcitriol|Drug|false|false||CALCITRIOL
null|Calcitriol Drug Class|Drug|false|false||CALCITRIOLnull|microgram|LabModifier|false|false||mcgnull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Every - dosing instruction fragment|Finding|false|false||everynull|Every (qualifier)|Modifier|false|false||everynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|citalopram|Drug|false|false||CITALOPRAM
null|citalopram|Drug|false|false||CITALOPRAMnull|Transaction counts and value totals - provider|Finding|false|false||Provider
null|Provider|Finding|false|false||Providernull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|clopidogrel|Drug|false|false||CLOPIDOGREL
null|clopidogrel|Drug|false|false||CLOPIDOGRELnull|Plavix|Drug|false|false||PLAVIX
null|Plavix|Drug|false|false||PLAVIXnull|Transaction counts and value totals - provider|Finding|false|false||Provider
null|Provider|Finding|false|false||Providernull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|folic acid|Drug|false|false||FOLIC ACID
null|folic acid|Drug|false|false||FOLIC ACID
null|folic acid|Drug|false|false||FOLIC ACIDnull|Folic acid measurement|Procedure|false|false||FOLIC ACIDnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Oral Route of Administration|Finding|true|false||by mouthnull|Oral cavity|Anatomy|true|false||mouth
null|Oral region|Anatomy|true|false||mouthnull|One Daily|Drug|true|false||one daily
null|One Daily|Drug|true|false||one daily
null|One Daily|Drug|true|false||one dailynull|Daily|Time|true|false||dailynull|Substitution - ActClass|Finding|true|false||Substitutionnull|Substitution - change|Event|true|false||Substitutionnull|lorazepam|Drug|true|false||LORAZEPAM
null|lorazepam|Drug|true|false||LORAZEPAMnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Hour|Time|false|false||hoursnull|Nausea|Finding|false|false||Nauseanull|null|Attribute|false|false||Nauseanull|metoprolol tartrate|Drug|false|false||METOPROLOL TARTRATE
null|metoprolol tartrate|Drug|false|false||METOPROLOL TARTRATEnull|metoprolol|Drug|false|false||METOPROLOL
null|metoprolol|Drug|false|false||METOPROLOLnull|tartrate|Drug|false|false||TARTRATE
null|Tartrates|Drug|false|false||TARTRATE
null|tartrate|Drug|false|false||TARTRATEnull|Lopressor|Drug|false|false||LOPRESSOR
null|Lopressor|Drug|false|false||LOPRESSORnull|Transaction counts and value totals - provider|Finding|false|false||Provider
null|Provider|Finding|false|false||Providernull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Oral Route of Administration|Finding|true|false||by mouthnull|Oral cavity|Anatomy|true|false||mouth
null|Oral region|Anatomy|true|false||mouthnull|BID protein, human|Drug|true|false||BID
null|BID protein, human|Drug|true|false||BIDnull|Body integrity dysphoria|Disorder|true|false||BIDnull|BID gene|Finding|true|false||BIDnull|Twice a day|Time|true|false||BIDnull|Substitution - ActClass|Finding|true|false||Substitutionnull|Substitution - change|Event|true|false||Substitutionnull|tramadol|Drug|true|false||TRAMADOL
null|tramadol|Drug|true|false||TRAMADOLnull|Tramadol measurement (procedure)|Procedure|true|false||TRAMADOLnull|Transaction counts and value totals - provider|Finding|false|false||Provider
null|Provider|Finding|false|false||Providernull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Three times daily|Time|false|false||three times a daynull|Thrice|LabModifier|false|false||three timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|trazodone|Drug|false|false||TRAZODONE
null|trazodone|Drug|false|false||TRAZODONEnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Oral Route of Administration|Finding|true|false||by mouthnull|Oral cavity|Anatomy|true|false||mouth
null|Oral region|Anatomy|true|false||mouthnull|One Daily|Drug|true|false||one daily
null|One Daily|Drug|true|false||one daily
null|One Daily|Drug|true|false||one dailynull|Daily|Time|true|false||dailynull|Substitution - ActClass|Finding|true|false||Substitutionnull|Substitution - change|Event|true|false||Substitutionnull|aspirin|Drug|true|false||ASPIRIN
null|aspirin|Drug|true|false||ASPIRINnull|Transaction counts and value totals - provider|Finding|false|false||Provider
null|Provider|Finding|false|false||Providernull|Chewable Tablet|Drug|false|false||Tablet, Chewablenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Oral Route of Administration|Finding|true|false||by mouthnull|Oral cavity|Anatomy|true|false||mouth
null|Oral region|Anatomy|true|false||mouthnull|One Daily|Drug|true|false||one daily
null|One Daily|Drug|true|false||one daily
null|One Daily|Drug|true|false||one dailynull|Daily|Time|true|false||dailynull|Substitution - ActClass|Finding|true|false||Substitutionnull|Substitution - change|Event|true|false||Substitutionnull|ranitidine hydrochloride|Drug|true|false||RANITIDINE HCL
null|ranitidine hydrochloride|Drug|true|false||RANITIDINE HCLnull|ranitidine|Drug|true|false||RANITIDINE
null|ranitidine|Drug|true|false||RANITIDINEnull|Flinders medical centre-7 marker|Drug|true|false||HCL
null|hydrochloride|Drug|true|false||HCL
null|hydrochloride|Drug|true|false||HCLnull|Hairy Cell Leukemia|Disorder|true|false||HCLnull|Acid Control|Drug|true|false||ACID CONTROL
null|Acid Control|Drug|true|false||ACID CONTROLnull|Control brand of phenylpropanolamine|Drug|false|false||CONTROL
null|CONTROL veterinary product|Drug|false|false||CONTROL
null|control substance|Drug|false|false||CONTROL
null|Control brand of phenylpropanolamine|Drug|false|false||CONTROLnull|Control - Relationship modifier|Finding|false|false||CONTROL
null|Control function|Finding|false|false||CONTROL
null|Scientific Control|Finding|false|false||CONTROLnull|Control Groups|Subject|false|false||CONTROLnull|True Control Status|Modifier|false|false||CONTROL
null|control aspects|Modifier|false|false||CONTROLnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Oral cavity|Anatomy|true|false||mouth
null|Oral region|Anatomy|true|false||mouthnull|One Daily|Drug|true|false||one daily
null|One Daily|Drug|true|false||one daily
null|One Daily|Drug|true|false||one dailynull|Daily|Time|true|false||dailynull|Substitution - ActClass|Finding|true|false||Substitutionnull|Substitution - change|Event|true|false||Substitutionnull|Medication.discharge|Finding|true|false||Discharge Medicationsnull|Body Substance Discharge|Finding|true|false||Discharge
null|Discharge Body Fluid|Finding|true|false||Discharge
null|Body Fluid Discharge|Finding|true|false||Discharge
null|null|Finding|true|false||Dischargenull|Patient Discharge|Procedure|true|false||Dischargenull|Pharmaceutical Preparations|Drug|true|false||Medicationsnull|Medications|Finding|true|false||Medicationsnull|null|Attribute|true|false||Medications
null|null|Attribute|true|false||Medicationsnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Certificate Status - Expired|Finding|false|false||Expired
null|Referral status - Expired|Finding|false|false||Expired
null|Cessation of life|Finding|false|false||Expired
null|Expiration, Respiratory|Finding|false|false||Expired
null|Expiration|Finding|false|false||Expirednull|Specimen Reject Reason - Expired|Modifier|false|false||Expirednull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Small cell carcinoma of lung|Disorder|false|false||small cell lung cancernull|Small|LabModifier|false|false||smallnull|CELP gene|Finding|false|false||cell
null|CEL gene|Finding|false|false||cellnull|Cells|Anatomy|false|false||cellnull|Cell Device|Device|false|false||cell
null|Cellular Phone|Device|false|false||cellnull|Cell (compartment)|Modifier|false|false||cellnull|Malignant neoplasm of lung|Disorder|false|false||lung cancer
null|Carcinoma of lung|Disorder|false|false||lung cancernull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Melena|Finding|false|false||Melenanull|Certificate Status - Expired|Finding|false|false||Expired
null|Referral status - Expired|Finding|false|false||Expired
null|Cessation of life|Finding|false|false||Expired
null|Expiration, Respiratory|Finding|false|false||Expired
null|Expiration|Finding|false|false||Expirednull|Specimen Reject Reason - Expired|Modifier|false|false||Expirednull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions