 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|39,48|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|39,48|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|39,53|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|73,82|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|73,82|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|73,82|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|73,82|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|73,82|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|73,87|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|105,110|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|105,110|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|105,110|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|129,132|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|140,147|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|140,147|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|149,157|true|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|Allergies|181,190|true|false|false|C1717415||Allergies
Event|Event|Allergies|181,190|true|false|false|||Allergies
Finding|Pathologic Function|Allergies|181,190|true|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|Allergies|193,215|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|Allergies|201,205|true|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|Allergies|201,205|true|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|Allergies|201,215|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Event|Event|Allergies|206,215|true|false|false|||Reactions
Event|Event|Allergies|218,227|false|false|false|||Attending
Finding|Functional Concept|Allergies|218,227|false|false|false|C1999232|Attending (action)|Attending
Event|Event|Chief Complaint|253,262|false|false|false|||shortness
Attribute|Clinical Attribute|Chief Complaint|253,272|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|Chief Complaint|253,272|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|Chief Complaint|266,272|false|false|false|C0225386|Breath|breath
Finding|Classification|Chief Complaint|275,280|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|281,289|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|281,289|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|293,311|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|302,311|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|302,311|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|302,311|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|302,311|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|302,311|false|false|false|C0184661|Interventional procedure|Procedure
Finding|Body Substance|History of Present Illness|349,356|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|349,356|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|349,356|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|History of Present Illness|371,378|false|false|false|||history
Finding|Conceptual Entity|History of Present Illness|371,378|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|371,378|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|371,378|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|371,381|false|false|false|C0262926|Medical History|history of
Attribute|Clinical Attribute|History of Present Illness|371,405|false|false|false|C1881055|Personal History of Coronary Artery Disease|history of coronary artery disease
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|382,390|false|false|false|C0018787|Heart|coronary
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|382,397|false|false|false|C0205042|Coronary artery|coronary artery
Disorder|Disease or Syndrome|History of Present Illness|382,405|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|coronary artery disease
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|391,397|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|History of Present Illness|391,397|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Disorder|Disease or Syndrome|History of Present Illness|391,405|false|false|false|C0852949|Arteriopathic disease|artery disease
Disorder|Disease or Syndrome|History of Present Illness|398,405|false|false|false|C0012634|Disease|disease
Event|Event|History of Present Illness|398,405|false|false|false|||disease
Finding|Functional Concept|History of Present Illness|410,418|false|false|false|C0475224|Ischemic|ischemic
Disorder|Disease or Syndrome|History of Present Illness|426,429|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|426,429|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|History of Present Illness|426,429|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|History of Present Illness|426,429|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|History of Present Illness|426,429|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|History of Present Illness|426,429|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Event|Event|History of Present Illness|426,429|false|false|false|||DES
Finding|Gene or Genome|History of Present Illness|426,429|false|false|false|C1413980|DES gene|DES
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|433,436|false|false|false|C2987138|Methylcytosine Dioxygenase TET1|LCX
Drug|Enzyme|History of Present Illness|433,436|false|false|false|C2987138|Methylcytosine Dioxygenase TET1|LCX
Event|Event|History of Present Illness|433,436|false|false|false|||LCX
Finding|Gene or Genome|History of Present Illness|433,436|false|false|false|C1428863;C2987137|TET1 gene;TET1 wt Allele|LCX
Procedure|Diagnostic Procedure|History of Present Illness|442,445|false|false|false|C0430462|Transthoracic echocardiography|TTE
Finding|Intellectual Product|History of Present Illness|455,459|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Organ or Tissue Function|History of Present Illness|472,480|false|false|false|C0039155|Systole|systolic
Finding|Pathologic Function|History of Present Illness|472,492|false|false|false|C0749225|Systolic dysfunction|systolic dysfunction
Disorder|Disease or Syndrome|History of Present Illness|481,492|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Event|Event|History of Present Illness|481,492|false|false|false|||dysfunction
Finding|Conceptual Entity|History of Present Illness|481,492|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|History of Present Illness|481,492|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|History of Present Illness|481,492|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|495,500|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|History of Present Illness|495,500|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|History of Present Illness|495,500|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|History of Present Illness|495,508|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Event|Event|History of Present Illness|501,508|false|false|false|||failure
Finding|Functional Concept|History of Present Illness|501,508|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|History of Present Illness|501,508|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|History of Present Illness|501,508|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Attribute|Clinical Attribute|History of Present Illness|524,532|false|false|false|C0812388|Ejection time|ejection
Event|Event|History of Present Illness|524,532|false|false|false|||ejection
Finding|Daily or Recreational Activity|History of Present Illness|524,532|false|false|false|C0336969|Ejection as a Sports activity|ejection
Phenomenon|Phenomenon or Process|History of Present Illness|524,532|false|false|false|C0302131|Ejection as a Circumstance of Injury|ejection
Event|Event|History of Present Illness|533,541|false|false|false|||fraction
Finding|Intellectual Product|History of Present Illness|533,541|false|false|false|C1554103|MDFAttributeType - Fraction|fraction
Attribute|Clinical Attribute|History of Present Illness|543,547|false|false|false|C0428772|Left ventricular ejection fraction|LVEF
Event|Event|History of Present Illness|543,547|false|false|false|||LVEF
Procedure|Diagnostic Procedure|History of Present Illness|543,547|false|false|false|C3837267|LVEF (procedure)|LVEF
Disorder|Disease or Syndrome|History of Present Illness|557,584|false|false|false|C0085096|Peripheral Vascular Diseases|peripheral vascular disease
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|568,576|false|false|false|C0005847|Blood Vessel|vascular
Disorder|Disease or Syndrome|History of Present Illness|568,584|false|false|false|C0042373|Vascular Diseases|vascular disease
Disorder|Disease or Syndrome|History of Present Illness|577,584|false|false|false|C0012634|Disease|disease
Event|Event|History of Present Illness|577,584|false|false|false|||disease
Disorder|Disease or Syndrome|History of Present Illness|577,593|false|false|false|C0008679|Chronic disease|disease, chronic
Event|Event|History of Present Illness|586,593|false|false|false|||chronic
Finding|Intellectual Product|History of Present Illness|586,593|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|History of Present Illness|586,593|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|594,600|false|false|false|C0022646;C0227665|Both kidneys;Kidney|kidney
Disorder|Neoplastic Process|History of Present Illness|594,600|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|kidney
Event|Event|History of Present Illness|594,600|false|false|false|||kidney
Finding|Sign or Symptom|History of Present Illness|594,600|false|false|false|C0812426|Kidney problem|kidney
Procedure|Diagnostic Procedure|History of Present Illness|594,600|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|594,600|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Disorder|Disease or Syndrome|History of Present Illness|594,608|false|false|false|C0022658|Kidney Diseases|kidney disease
Disorder|Disease or Syndrome|History of Present Illness|601,608|false|false|false|C0012634|Disease|disease
Event|Event|History of Present Illness|601,608|false|false|false|||disease
Attribute|Clinical Attribute|History of Present Illness|610,615|false|true|false|C1300072|Tumor stage|stage
Anatomy|Body Location or Region|History of Present Illness|638,641|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|History of Present Illness|638,641|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|History of Present Illness|638,641|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Finding|Finding|History of Present Illness|646,652|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|History of Present Illness|646,652|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Event|Event|History of Present Illness|653,657|false|false|false|||UGIB
Disorder|Disease or Syndrome|History of Present Illness|671,674|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|History of Present Illness|671,674|false|false|false|||HTN
Disorder|Disease or Syndrome|History of Present Illness|676,688|false|false|false|C0242339|Dyslipidemias|dyslipidemia
Event|Event|History of Present Illness|676,688|false|false|false|||dyslipidemia
Event|Event|History of Present Illness|703,711|false|false|false|||presents
Finding|Finding|History of Present Illness|717,729|false|false|false|C3845714|Several days|several days
Event|Event|History of Present Illness|725,729|false|false|false|||days
Event|Event|History of Present Illness|733,742|false|false|false|||shortness
Attribute|Clinical Attribute|History of Present Illness|733,752|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|History of Present Illness|733,752|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|History of Present Illness|746,752|false|false|false|C0225386|Breath|breath
Event|Event|History of Present Illness|769,773|false|false|false|||says
Event|Event|History of Present Illness|789,796|false|false|false|||noticed
Finding|Intellectual Product|History of Present Illness|804,809|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Intellectual Product|History of Present Illness|804,815|false|false|false|C1272517|Sudden onset (contextual qualifier) (qualifier value)|acute onset
Event|Event|History of Present Illness|816,823|false|false|false|||dyspnea
Finding|Finding|History of Present Illness|816,823|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|History of Present Illness|816,823|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Event|Event|History of Present Illness|824,832|false|false|false|||starting
Event|Event|History of Present Illness|852,856|false|false|false|||walk
Event|Event|History of Present Illness|864,870|false|false|false|||stairs
Finding|Finding|History of Present Illness|864,870|false|false|false|C4300351|Prior functioning.stairs|stairs
Event|Event|History of Present Illness|878,882|false|false|false|||home
Finding|Idea or Concept|History of Present Illness|878,882|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|History of Present Illness|878,882|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|History of Present Illness|878,882|false|false|false|C1553498|home health encounter|home
Event|Event|History of Present Illness|897,900|false|false|false|||sit
Finding|Finding|History of Present Illness|897,900|false|false|false|C0277814;C0728713;C1539668;C1539774|Does sit;HHAT gene;SIT1 gene;Sitting position|sit
Finding|Gene or Genome|History of Present Illness|897,900|false|false|false|C0277814;C0728713;C1539668;C1539774|Does sit;HHAT gene;SIT1 gene;Sitting position|sit
Finding|Body Substance|History of Present Illness|920,926|false|false|false|C0225386|Breath|breath
Event|Event|History of Present Illness|961,965|false|false|false|||able
Finding|Finding|History of Present Illness|961,965|false|false|false|C1299581|Able (qualifier value)|able
Event|Event|History of Present Illness|969,974|true|false|false|||mount
Event|Event|History of Present Illness|982,988|true|false|false|||stairs
Finding|Finding|History of Present Illness|982,988|true|false|false|C4300351|Prior functioning.stairs|stairs
Event|Event|History of Present Illness|997,1007|true|false|false|||difficulty
Finding|Finding|History of Present Illness|997,1007|true|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Finding|Body Substance|History of Present Illness|1010,1017|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|1010,1017|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|1010,1017|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|History of Present Illness|1018,1024|true|false|false|||denies
Anatomy|Body Location or Region|History of Present Illness|1040,1045|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|1040,1045|true|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|1040,1050|true|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|1040,1050|true|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|1046,1050|true|false|false|C2598155||pain
Event|Event|History of Present Illness|1046,1050|true|false|false|||pain
Finding|Functional Concept|History of Present Illness|1046,1050|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1046,1050|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|1054,1066|true|false|false|||palpitations
Finding|Finding|History of Present Illness|1054,1066|true|false|false|C0030252|Palpitations|palpitations
Event|Event|History of Present Illness|1072,1081|true|false|false|||dizziness
Finding|Sign or Symptom|History of Present Illness|1072,1081|true|false|false|C0012833;C0042571|Dizziness;Vertigo|dizziness
Event|Event|History of Present Illness|1085,1100|true|false|false|||lightheadedness
Finding|Sign or Symptom|History of Present Illness|1085,1100|true|false|false|C0220870|Lightheadedness|lightheadedness
Finding|Body Substance|History of Present Illness|1103,1110|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|1103,1110|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|1103,1110|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|History of Present Illness|1119,1125|true|false|false|||denies
Drug|Organic Chemical|History of Present Illness|1130,1135|true|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|1130,1135|true|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|History of Present Illness|1130,1135|true|false|false|||cough
Finding|Sign or Symptom|History of Present Illness|1130,1135|true|false|false|C0010200|Coughing|cough
Event|Event|History of Present Illness|1137,1143|true|false|false|||fevers
Finding|Sign or Symptom|History of Present Illness|1137,1143|true|false|false|C0015967|Fever|fevers
Event|Event|History of Present Illness|1144,1150|true|false|false|||chills
Finding|Sign or Symptom|History of Present Illness|1144,1150|true|false|false|C0085593|Chills|chills
Anatomy|Body Location or Region|History of Present Illness|1165,1170|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|1165,1170|false|false|false|C0741025|Chest problem|chest
Finding|Sign or Symptom|History of Present Illness|1165,1181|false|false|false|C0235710|Chest discomfort|chest discomfort
Event|Event|History of Present Illness|1171,1181|false|false|false|||discomfort
Finding|Sign or Symptom|History of Present Illness|1171,1181|false|false|false|C2364135|Discomfort|discomfort
Event|Event|History of Present Illness|1212,1220|true|false|false|||symptoms
Finding|Functional Concept|History of Present Illness|1212,1220|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|History of Present Illness|1212,1220|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|History of Present Illness|1221,1231|true|false|false|||consistent
Finding|Idea or Concept|History of Present Illness|1221,1231|true|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|History of Present Illness|1221,1236|true|false|false|C0332290|Consistent with|consistent with
Event|Event|History of Present Illness|1237,1246|true|false|false|||orthopnea
Finding|Finding|History of Present Illness|1237,1246|true|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Finding|Sign or Symptom|History of Present Illness|1237,1246|true|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Disorder|Disease or Syndrome|History of Present Illness|1250,1253|true|false|false|C1956415|Paroxysmal nocturnal dyspnea|PND
Event|Event|History of Present Illness|1250,1253|true|false|false|||PND
Finding|Gene or Genome|History of Present Illness|1250,1253|true|false|false|C1417807;C4552608|NPPA gene;NPPA wt Allele|PND
Event|Event|History of Present Illness|1259,1268|true|false|false|||increased
Event|Event|History of Present Illness|1273,1281|true|false|false|||swelling
Finding|Finding|History of Present Illness|1273,1281|true|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|History of Present Illness|1273,1281|true|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Body Substance|History of Present Illness|1283,1290|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1283,1290|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1283,1290|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|1291,1296|false|false|false|||notes
Event|Event|History of Present Illness|1310,1321|false|false|false|||experienced
Finding|Body Substance|History of Present Illness|1343,1350|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|1343,1350|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|1343,1350|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|History of Present Illness|1351,1356|false|false|false|||takes
Attribute|Clinical Attribute|History of Present Illness|1361,1367|false|false|false|C0944911||weight
Event|Event|History of Present Illness|1361,1367|false|false|false|||weight
Finding|Finding|History of Present Illness|1361,1367|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|History of Present Illness|1361,1367|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|History of Present Illness|1361,1367|false|false|false|C1305866|Weighing patient|weight
Finding|Finding|History of Present Illness|1368,1384|false|false|false|C5202779|True or Present Nearly Every Day|nearly every day
Finding|Idea or Concept|History of Present Illness|1381,1384|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|History of Present Illness|1381,1384|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Attribute|Clinical Attribute|History of Present Illness|1400,1406|false|false|false|C0944911||weight
Event|Event|History of Present Illness|1400,1406|false|false|false|||weight
Finding|Finding|History of Present Illness|1400,1406|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|History of Present Illness|1400,1406|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|History of Present Illness|1400,1406|false|false|false|C1305866|Weighing patient|weight
Finding|Intellectual Product|History of Present Illness|1426,1430|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|History of Present Illness|1461,1471|false|false|false|||attributes
Drug|Organic Chemical|History of Present Illness|1526,1535|true|false|false|C0076840|torsemide|torsemide
Drug|Pharmacologic Substance|History of Present Illness|1526,1535|true|false|false|C0076840|torsemide|torsemide
Event|Event|History of Present Illness|1526,1535|true|false|false|||torsemide
Event|Event|History of Present Illness|1555,1560|true|false|false|||doses
Event|Event|History of Present Illness|1566,1572|true|false|false|||issues
Anatomy|Body Location or Region|History of Present Illness|1578,1587|true|false|false|C0000726|Abdomen|abdominal
Finding|Finding|History of Present Illness|1578,1596|true|false|false|C0000731;C1291077|Abdomen distended;Abdominal bloating|abdominal bloating
Finding|Sign or Symptom|History of Present Illness|1578,1596|true|false|false|C0000731;C1291077|Abdomen distended;Abdominal bloating|abdominal bloating
Event|Event|History of Present Illness|1588,1596|true|false|false|||bloating
Finding|Finding|History of Present Illness|1588,1596|true|false|false|C0000731;C1291077|Abdomen distended;Abdominal bloating|bloating
Finding|Sign or Symptom|History of Present Illness|1588,1596|true|false|false|C0000731;C1291077|Abdomen distended;Abdominal bloating|bloating
Event|Event|History of Present Illness|1600,1612|true|false|false|||constipation
Finding|Sign or Symptom|History of Present Illness|1600,1612|true|false|false|C0009806|Constipation|constipation
Event|Event|History of Present Illness|1625,1631|true|false|false|||travel
Finding|Daily or Recreational Activity|History of Present Illness|1625,1631|true|false|false|C0040802|travel|travel
Procedure|Health Care Activity|History of Present Illness|1625,1631|true|false|false|C1555670|travel charge|travel
Finding|Body Substance|History of Present Illness|1635,1642|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|1635,1642|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|1635,1642|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|History of Present Illness|1658,1667|false|false|false|||recovered
Finding|Functional Concept|History of Present Illness|1675,1680|false|false|false|C0521026|Viral|viral
Disorder|Disease or Syndrome|History of Present Illness|1681,1684|false|false|false|C0041912|Upper Respiratory Infections|URI
Event|Event|History of Present Illness|1681,1684|false|false|false|||URI
Finding|Gene or Genome|History of Present Illness|1681,1684|false|false|false|C1421895;C1548524;C3272713|URI1 gene;URI1 wt Allele;Uniform Resource Identifier|URI
Finding|Intellectual Product|History of Present Illness|1681,1684|false|false|false|C1421895;C1548524;C3272713|URI1 gene;URI1 wt Allele;Uniform Resource Identifier|URI
Finding|Idea or Concept|History of Present Illness|1705,1712|false|false|false|C1555582|Initial (abbreviation)|initial
Event|Event|History of Present Illness|1752,1756|false|false|false|||Exam
Finding|Functional Concept|History of Present Illness|1752,1756|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|History of Present Illness|1752,1756|false|false|false|C0582103|Medical Examination|Exam
Event|Event|History of Present Illness|1788,1796|false|false|false|||wheezing
Finding|Sign or Symptom|History of Present Illness|1788,1796|false|false|false|C0043144|Wheezing|wheezing
Event|Event|History of Present Illness|1807,1813|true|false|false|||volume
Finding|Intellectual Product|History of Present Illness|1807,1813|true|false|false|C1705102|Volume (publication)|volume
Finding|Pathologic Function|History of Present Illness|1807,1822|true|false|false|C0546817|Hypervolemia (finding)|volume overload
Event|Event|History of Present Illness|1814,1822|true|false|false|||overload
Event|Event|History of Present Illness|1827,1830|false|false|false|||EKG
Finding|Intellectual Product|History of Present Illness|1827,1830|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|History of Present Illness|1827,1830|false|false|false|C1623258|Electrocardiography|EKG
Event|Event|History of Present Illness|1832,1835|false|false|false|||NSR
Finding|Molecular Function|History of Present Illness|1832,1835|false|false|false|C1704493;C2700623|Neutral Sidebent Rotated|NSR
Finding|Pathologic Function|History of Present Illness|1832,1835|false|false|false|C1704493;C2700623|Neutral Sidebent Rotated|NSR
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1852,1856|false|false|false|C0004457|Axis vertebra|axis
Disorder|Injury or Poisoning|History of Present Illness|1852,1856|false|false|false|C0349013|Fracture of second cervical vertebra|axis
Event|Event|History of Present Illness|1872,1881|false|false|false|||intervals
Phenomenon|Natural Phenomenon or Process|History of Present Illness|1894,1899|false|false|false|C0678544||waves
Event|Event|History of Present Illness|1909,1913|false|false|false|||TWIs
Event|Event|History of Present Illness|1929,1934|true|false|false|||submm
Disorder|Disease or Syndrome|History of Present Illness|1943,1947|true|false|false|C0036916|Sexually Transmitted Diseases|STDs
Event|Event|History of Present Illness|1943,1947|true|false|false|||STDs
Event|Event|History of Present Illness|1953,1957|true|false|false|||STEs
Event|Event|History of Present Illness|1960,1964|false|false|false|||Labs
Lab|Laboratory or Test Result|History of Present Illness|1960,1964|false|false|false|C0587081|Laboratory test finding|Labs
Event|Event|History of Present Illness|1965,1971|false|false|false|||showed
Anatomy|Cell Component|History of Present Illness|1975,1978|false|false|false|C2263086|Nuclear cap binding complex location|CBC
Procedure|Laboratory Procedure|History of Present Illness|1975,1978|false|false|false|C0009555|Complete Blood Count|CBC
Disorder|Virus|History of Present Illness|2009,2012|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|History of Present Illness|2009,2012|false|false|false|||MCV
Lab|Laboratory or Test Result|History of Present Illness|2009,2012|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|History of Present Illness|2009,2012|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|2009,2012|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|2017,2020|false|false|false|C0053932|Bone Morphogenetic Proteins|BMP
Drug|Biologically Active Substance|History of Present Illness|2017,2020|false|false|false|C0053932|Bone Morphogenetic Proteins|BMP
Event|Event|History of Present Illness|2017,2020|false|false|false|||BMP
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|2017,2020|false|false|false|C0279266|carmustine/methotrexate/procarbazine protocol|BMP
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|2055,2061|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Drug|Hormone|History of Present Illness|2055,2061|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Event|Event|History of Present Illness|2067,2070|false|false|false|||VBG
Drug|Biologically Active Substance|History of Present Illness|2101,2113|false|false|false|C0042052|Urobilinogen|urobilinogen
Drug|Organic Chemical|History of Present Illness|2101,2113|false|false|false|C0042052|Urobilinogen|urobilinogen
Event|Event|History of Present Illness|2101,2113|false|false|false|||urobilinogen
Procedure|Laboratory Procedure|History of Present Illness|2101,2113|false|false|false|C0202241|Urobilinogen measurement|urobilinogen
Event|Event|History of Present Illness|2114,2117|false|false|false|||NEG
Finding|Finding|History of Present Illness|2114,2117|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|History of Present Illness|2119,2128|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|bilirubin
Drug|Organic Chemical|History of Present Illness|2119,2128|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|bilirubin
Drug|Pharmacologic Substance|History of Present Illness|2119,2128|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|bilirubin
Event|Event|History of Present Illness|2119,2128|false|false|false|||bilirubin
Procedure|Laboratory Procedure|History of Present Illness|2119,2128|false|false|false|C0201913;C0863174|Bilirubin, total measurement;blood bilirubin level test|bilirubin
Event|Event|History of Present Illness|2129,2132|false|false|false|||NEG
Finding|Finding|History of Present Illness|2129,2132|false|false|false|C5848551|Neg - answer|NEG
Event|Event|History of Present Illness|2139,2142|false|false|false|||NEG
Finding|Finding|History of Present Illness|2139,2142|false|false|false|C5848551|Neg - answer|NEG
Disorder|Disease or Syndrome|History of Present Illness|2144,2149|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|History of Present Illness|2144,2149|false|false|false|||blood
Finding|Body Substance|History of Present Illness|2144,2149|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Event|History of Present Illness|2150,2153|false|false|false|||NEG
Finding|Finding|History of Present Illness|2150,2153|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|History of Present Illness|2155,2162|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|nitrite
Drug|Inorganic Chemical|History of Present Illness|2155,2162|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|nitrite
Drug|Pharmacologic Substance|History of Present Illness|2155,2162|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|nitrite
Event|Event|History of Present Illness|2163,2166|false|false|false|||NEG
Finding|Finding|History of Present Illness|2163,2166|false|false|false|C5848551|Neg - answer|NEG
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|2168,2175|false|false|false|C0033684|Proteins|protein
Drug|Biologically Active Substance|History of Present Illness|2168,2175|false|false|false|C0033684|Proteins|protein
Event|Event|History of Present Illness|2168,2175|false|false|false|||protein
Finding|Conceptual Entity|History of Present Illness|2168,2175|false|false|false|C1521746|Protein Info|protein
Procedure|Laboratory Procedure|History of Present Illness|2168,2175|false|false|false|C0202202|Protein measurement|protein
Drug|Biologically Active Substance|History of Present Illness|2181,2188|false|false|false|C0017725|glucose|glucose
Drug|Organic Chemical|History of Present Illness|2181,2188|false|false|false|C0017725|glucose|glucose
Drug|Pharmacologic Substance|History of Present Illness|2181,2188|false|false|false|C0017725|glucose|glucose
Lab|Laboratory or Test Result|History of Present Illness|2181,2188|false|false|false|C5781949|Glucose^1.5H post dose glucagon|glucose
Procedure|Laboratory Procedure|History of Present Illness|2181,2188|false|false|false|C0337438|Glucose measurement|glucose
Event|Event|History of Present Illness|2189,2192|false|false|false|||NEG
Finding|Finding|History of Present Illness|2189,2192|false|false|false|C5848551|Neg - answer|NEG
Disorder|Injury or Poisoning|History of Present Illness|2194,2201|false|false|false|C0497010|Toxic effect of ketones|ketones
Drug|Organic Chemical|History of Present Illness|2194,2201|false|false|false|C0022634|Ketones|ketones
Event|Event|History of Present Illness|2194,2201|false|false|false|||ketones
Procedure|Laboratory Procedure|History of Present Illness|2194,2201|false|false|false|C0202110;C0555179|Ketone bodies measurement, quantitative;Urine ketone test|ketones
Event|Event|History of Present Illness|2202,2205|false|false|false|||NEG
Finding|Finding|History of Present Illness|2202,2205|false|false|false|C5848551|Neg - answer|NEG
Anatomy|Cell|History of Present Illness|2207,2210|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|History of Present Illness|2207,2210|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|History of Present Illness|2207,2210|false|false|false|C0014792|Erythrocytes|RBC
Anatomy|Cell|History of Present Illness|2214,2217|false|false|false|C0023516|Leukocytes|WBC
Event|Event|History of Present Illness|2225,2233|false|false|false|||bacteria
Finding|Functional Concept|History of Present Illness|2225,2233|false|false|false|C1510439|bacteria aspects|bacteria
Event|Event|History of Present Illness|2235,2242|false|false|false|||Imaging
Finding|Finding|History of Present Illness|2235,2242|false|false|false|C0740845|Imaging problem|Imaging
Procedure|Diagnostic Procedure|History of Present Illness|2235,2242|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|Imaging
Event|Event|History of Present Illness|2243,2249|false|false|false|||showed
Event|Event|History of Present Illness|2252,2255|false|false|false|||CXR
Procedure|Diagnostic Procedure|History of Present Illness|2252,2255|false|false|false|C0039985|Plain chest X-ray|CXR
Anatomy|Body Part, Organ, or Organ Component|Findings|2272,2277|false|false|false|C0024109|Lung|Lungs
Finding|Finding|Findings|2282,2292|false|false|false|C4085643;C5201148;C5962468|Moderate;Moderate Effect;Moderate Response|moderately
Finding|Finding|Findings|2293,2297|false|false|false|C5575035|Well (answer to question)|well
Event|Event|Findings|2298,2306|false|false|false|||expanded
Event|Event|Findings|2331,2336|false|false|false|||right
Finding|Functional Concept|Findings|2331,2336|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|Findings|2337,2342|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|Findings|2337,2342|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Location or Region|Findings|2343,2347|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Findings|2343,2347|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Findings|2343,2347|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Findings|2343,2347|false|false|false|C0740941|Lung Problem|lung
Finding|Finding|Findings|2343,2355|false|false|false|C4728208|Lung opacity|lung opacity
Event|Event|Findings|2348,2355|false|false|false|||opacity
Finding|Finding|Findings|2348,2355|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacity
Finding|Pathologic Function|Findings|2348,2355|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacity
Event|Event|Findings|2357,2360|false|false|false|||new
Finding|Finding|Findings|2357,2360|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Findings|2357,2360|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Anatomy|Body Part, Organ, or Organ Component|Findings|2375,2380|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Findings|2375,2380|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Event|Event|Findings|2375,2380|false|false|false|||heart
Finding|Sign or Symptom|Findings|2375,2380|false|false|false|C0795691|HEART PROBLEM|heart
Event|Event|Findings|2396,2404|false|false|false|||enlarged
Procedure|Therapeutic or Preventive Procedure|Findings|2396,2404|false|false|false|C1293134|Enlargement procedure|enlarged
Finding|Intellectual Product|Findings|2418,2422|false|false|false|C1547225|Mild Severity of Illness Code|mild
Anatomy|Body Part, Organ, or Organ Component|Findings|2423,2432|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Findings|2423,2432|false|false|false|C2707265||pulmonary
Finding|Finding|Findings|2423,2432|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Disorder|Disease or Syndrome|Findings|2423,2452|false|false|false|C5849517|Pulmonary vascular congestion|pulmonary vascular congestion
Anatomy|Body Part, Organ, or Organ Component|Findings|2433,2441|false|false|false|C0005847|Blood Vessel|vascular
Event|Event|Findings|2442,2452|false|false|false|||congestion
Finding|Pathologic Function|Findings|2442,2452|false|false|false|C0700148|Congestion|congestion
Anatomy|Tissue|Findings|2457,2464|true|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|Findings|2457,2464|true|false|false|C0032226|Pleural Diseases|pleural
Finding|Body Substance|Findings|2457,2473|true|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Finding|Findings|2457,2473|true|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Pathologic Function|Findings|2457,2473|true|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Event|Event|Findings|2465,2473|true|false|false|||effusion
Finding|Body Substance|Findings|2465,2473|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|Findings|2465,2473|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|Findings|2465,2473|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Disorder|Disease or Syndrome|Findings|2477,2489|true|false|false|C0032326|Pneumothorax|pneumothorax
Event|Event|Findings|2477,2489|true|false|false|||pneumothorax
Finding|Functional Concept|Impression|2506,2511|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Part, Organ, or Organ Component|Impression|2506,2522|false|false|false|C1261075|Structure of right lower lobe of lung|Right lower lobe
Anatomy|Body Location or Region|Impression|2512,2517|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|Impression|2512,2517|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|Impression|2512,2522|false|false|false|C0225758|Structure of lower lobe of lung|lower lobe
Anatomy|Body Part, Organ, or Organ Component|Impression|2518,2522|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|Impression|2518,2522|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Event|Event|Impression|2523,2530|false|false|false|||opacity
Finding|Finding|Impression|2523,2530|false|true|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacity
Finding|Pathologic Function|Impression|2523,2530|false|true|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacity
Event|Event|Impression|2537,2546|false|false|false|||represent
Disorder|Disease or Syndrome|Impression|2547,2556|false|true|false|C0032285|Pneumonia|pneumonia
Event|Event|Impression|2547,2556|false|false|false|||pneumonia
Finding|Functional Concept|Impression|2564,2569|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Finding|Intellectual Product|Impression|2570,2578|false|false|false|C1315013|Clinical NEC (not elsewhere classified in LNC)|clinical
Event|Event|Impression|2579,2586|false|false|false|||setting
Finding|Mental Process|Impression|2579,2586|false|false|false|C0542559|contextual factors|setting
Event|Event|Impression|2597,2608|false|false|false|||atelectasis
Finding|Pathologic Function|Impression|2597,2608|false|false|false|C0004144|Atelectasis|atelectasis
Anatomy|Body Part, Organ, or Organ Component|Impression|2623,2632|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Impression|2623,2632|false|false|false|C2707265||pulmonary
Finding|Finding|Impression|2623,2632|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Attribute|Clinical Attribute|Impression|2633,2638|false|false|false|C1717255||edema
Event|Event|Impression|2633,2638|false|false|false|||edema
Finding|Pathologic Function|Impression|2633,2638|false|false|false|C0013604|Edema|edema
Event|Event|Impression|2645,2652|false|false|false|||account
Event|Event|Impression|2662,2669|false|false|false|||finding
Finding|Finding|Impression|2662,2669|false|true|false|C0037088;C0243095;C2825141|Experimental Finding;Finding;Signs and Symptoms|finding
Finding|Sign or Symptom|Impression|2662,2669|false|true|false|C0037088;C0243095;C2825141|Experimental Finding;Finding;Signs and Symptoms|finding
Event|Event|Impression|2696,2701|false|false|false|||views
Event|Event|Impression|2711,2718|false|false|false|||helpful
Event|Activity|Impression|2731,2741|false|true|false|C1516048|Assessed|assessment
Event|Event|Impression|2731,2741|false|false|false|||assessment
Finding|Intellectual Product|Impression|2731,2741|false|true|false|C0679207|Knowledge acquisition using a method of assessment|assessment
Procedure|Diagnostic Procedure|Impression|2731,2741|false|true|false|C0028708;C0031809;C0220825;C0542573;C0549068;C0549070;C0549071;C0549072;C0549073;C0549074;C0549075;C0549076;C0549078;C0549079;C0549080;C1161151;C1261322;C2237115|Evaluation;Evaluation procedure;Nutrition Assessment;Personal care assessment;Physical Examination;assessment of cognitive functions|assessment
Procedure|Health Care Activity|Impression|2731,2741|false|true|false|C0028708;C0031809;C0220825;C0542573;C0549068;C0549070;C0549071;C0549072;C0549073;C0549074;C0549075;C0549076;C0549078;C0549079;C0549080;C1161151;C1261322;C2237115|Evaluation;Evaluation procedure;Nutrition Assessment;Personal care assessment;Physical Examination;assessment of cognitive functions|assessment
Event|Event|Impression|2746,2754|false|false|false|||Consults
Procedure|Health Care Activity|Impression|2746,2754|false|false|false|C0009818|Consultation|Consults
Finding|Body Substance|Impression|2764,2771|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Impression|2764,2771|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Impression|2764,2771|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Impression|2772,2780|true|false|false|||received
Drug|Organic Chemical|Impression|2797,2806|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|Impression|2797,2806|false|false|false|C0001927|albuterol|Albuterol
Drug|Amino Acid, Peptide, or Protein|Impression|2814,2817|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|Impression|2814,2817|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|Impression|2814,2817|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Finding|Cell Function|Impression|2814,2817|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|Impression|2814,2817|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|Impression|2825,2828|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|Impression|2825,2828|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|Impression|2825,2828|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|Impression|2825,2828|false|false|false|||NEB
Finding|Cell Function|Impression|2825,2828|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Impression|2825,2828|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Drug|Organic Chemical|Impression|2844,2853|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|Impression|2844,2853|false|false|false|C0001927|albuterol|Albuterol
Drug|Amino Acid, Peptide, or Protein|Impression|2861,2864|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|Impression|2861,2864|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|Impression|2861,2864|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Finding|Cell Function|Impression|2861,2864|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|Impression|2861,2864|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|Impression|2872,2875|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|Impression|2872,2875|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|Impression|2872,2875|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|Impression|2872,2875|false|false|false|||NEB
Finding|Cell Function|Impression|2872,2875|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Impression|2872,2875|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Drug|Organic Chemical|Impression|2891,2902|false|false|false|C0027235|ipratropium|Ipratropium
Drug|Pharmacologic Substance|Impression|2891,2902|false|false|false|C0027235|ipratropium|Ipratropium
Drug|Organic Chemical|Impression|2891,2910|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Pharmacologic Substance|Impression|2891,2910|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Inorganic Chemical|Impression|2903,2910|false|false|false|C0006222|Bromides|Bromide
Event|Event|Impression|2903,2910|false|false|false|||Bromide
Procedure|Laboratory Procedure|Impression|2903,2910|false|false|false|C0202341|Bromides measurement|Bromide
Drug|Amino Acid, Peptide, or Protein|Impression|2911,2914|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|Impression|2911,2914|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|Impression|2911,2914|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Finding|Cell Function|Impression|2911,2914|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|Impression|2911,2914|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|Impression|2917,2920|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|Impression|2917,2920|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|Impression|2917,2920|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|Impression|2917,2920|false|false|false|||NEB
Finding|Cell Function|Impression|2917,2920|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Impression|2917,2920|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Drug|Organic Chemical|Impression|2936,2945|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|Impression|2936,2945|false|false|false|C0001927|albuterol|Albuterol
Drug|Amino Acid, Peptide, or Protein|Impression|2953,2956|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|Impression|2953,2956|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|Impression|2953,2956|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Finding|Cell Function|Impression|2953,2956|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|Impression|2953,2956|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|Impression|2964,2967|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|Impression|2964,2967|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|Impression|2964,2967|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|Impression|2964,2967|false|false|false|||NEB
Finding|Cell Function|Impression|2964,2967|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Impression|2964,2967|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Drug|Organic Chemical|Impression|2982,2993|false|false|false|C0027235|ipratropium|Ipratropium
Drug|Pharmacologic Substance|Impression|2982,2993|false|false|false|C0027235|ipratropium|Ipratropium
Drug|Organic Chemical|Impression|2982,3001|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Pharmacologic Substance|Impression|2982,3001|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Inorganic Chemical|Impression|2994,3001|false|false|false|C0006222|Bromides|Bromide
Event|Event|Impression|2994,3001|false|false|false|||Bromide
Procedure|Laboratory Procedure|Impression|2994,3001|false|false|false|C0202341|Bromides measurement|Bromide
Drug|Amino Acid, Peptide, or Protein|Impression|3002,3005|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|Impression|3002,3005|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|Impression|3002,3005|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Event|Event|Impression|3002,3005|false|false|false|||Neb
Finding|Cell Function|Impression|3002,3005|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|Impression|3002,3005|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|Impression|3008,3011|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|Impression|3008,3011|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|Impression|3008,3011|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|Impression|3008,3011|false|false|false|||NEB
Finding|Cell Function|Impression|3008,3011|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Impression|3008,3011|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Drug|Antibiotic|Impression|3026,3038|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Drug|Clinical Drug|Impression|3026,3038|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Drug|Organic Chemical|Impression|3026,3038|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Event|Event|Impression|3026,3038|false|false|false|||Azithromycin
Drug|Antibiotic|Impression|3053,3064|false|false|false|C0007561|ceftriaxone|CefTRIAXone
Drug|Organic Chemical|Impression|3053,3064|false|false|false|C0007561|ceftriaxone|CefTRIAXone
Event|Event|Impression|3053,3064|false|false|false|||CefTRIAXone
Drug|Hormone|Impression|3078,3088|false|false|false|C0032952|prednisone|PredniSONE
Drug|Organic Chemical|Impression|3078,3088|false|false|false|C0032952|prednisone|PredniSONE
Drug|Pharmacologic Substance|Impression|3078,3088|false|false|false|C0032952|prednisone|PredniSONE
Drug|Organic Chemical|Impression|3108,3118|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|Impression|3108,3118|false|false|false|C0016860|furosemide|Furosemide
Event|Event|Impression|3108,3118|false|false|false|||Furosemide
Drug|Antibiotic|Impression|3139,3150|false|false|false|C0007561|ceftriaxone|CefTRIAXone
Drug|Organic Chemical|Impression|3139,3150|false|false|false|C0007561|ceftriaxone|CefTRIAXone
Drug|Antibiotic|Impression|3171,3183|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Drug|Clinical Drug|Impression|3171,3183|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Drug|Organic Chemical|Impression|3171,3183|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Event|Event|Impression|3171,3183|false|false|false|||Azithromycin
Drug|Organic Chemical|Impression|3242,3252|false|false|false|C0054836|carvedilol|Carvedilol
Drug|Pharmacologic Substance|Impression|3242,3252|false|false|false|C0054836|carvedilol|Carvedilol
Event|Event|Impression|3242,3252|false|false|false|||Carvedilol
Drug|Organic Chemical|Impression|3272,3282|false|false|false|C0028066|nifedipine|NIFEdipine
Drug|Pharmacologic Substance|Impression|3272,3282|false|false|false|C0028066|nifedipine|NIFEdipine
Event|Event|Impression|3272,3282|false|false|false|||NIFEdipine
Finding|Finding|Impression|3284,3292|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Impression|3284,3292|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Impression|3293,3300|false|false|false|||Release
Finding|Functional Concept|Impression|3293,3300|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Impression|3293,3300|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Impression|3293,3300|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Impression|3322,3331|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|Impression|3322,3331|false|false|false|C0001927|albuterol|Albuterol
Drug|Amino Acid, Peptide, or Protein|Impression|3339,3342|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|Impression|3339,3342|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|Impression|3339,3342|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Finding|Cell Function|Impression|3339,3342|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|Impression|3339,3342|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|Impression|3350,3353|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|Impression|3350,3353|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|Impression|3350,3353|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|Impression|3350,3353|false|false|false|||NEB
Finding|Cell Function|Impression|3350,3353|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Impression|3350,3353|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Drug|Organic Chemical|Impression|3368,3379|false|false|false|C0027235|ipratropium|Ipratropium
Drug|Pharmacologic Substance|Impression|3368,3379|false|false|false|C0027235|ipratropium|Ipratropium
Drug|Organic Chemical|Impression|3368,3387|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Pharmacologic Substance|Impression|3368,3387|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Inorganic Chemical|Impression|3380,3387|false|false|false|C0006222|Bromides|Bromide
Event|Event|Impression|3380,3387|false|false|false|||Bromide
Procedure|Laboratory Procedure|Impression|3380,3387|false|false|false|C0202341|Bromides measurement|Bromide
Drug|Amino Acid, Peptide, or Protein|Impression|3388,3391|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|Impression|3388,3391|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|Impression|3388,3391|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Finding|Cell Function|Impression|3388,3391|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|Impression|3388,3391|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|Impression|3394,3397|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|Impression|3394,3397|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|Impression|3394,3397|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|Impression|3394,3397|false|false|false|||NEB
Finding|Cell Function|Impression|3394,3397|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Impression|3394,3397|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Drug|Organic Chemical|Impression|3414,3424|false|false|false|C0060926|gabapentin|Gabapentin
Drug|Pharmacologic Substance|Impression|3414,3424|false|false|false|C0060926|gabapentin|Gabapentin
Event|Event|Impression|3414,3424|false|false|false|||Gabapentin
Drug|Amino Acid, Peptide, or Protein|Impression|3445,3452|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Hormone|Impression|3445,3452|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Pharmacologic Substance|Impression|3445,3452|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Event|Event|Impression|3445,3452|false|false|false|||Insulin
Finding|Gene or Genome|Impression|3445,3452|false|false|false|C1337112|INS gene|Insulin
Procedure|Laboratory Procedure|Impression|3445,3452|false|false|false|C0202098|Insulin measurement|Insulin
Event|Event|Impression|3455,3460|false|false|false|||Units
Event|Event|Impression|3462,3470|false|false|false|||Transfer
Finding|Functional Concept|Impression|3462,3470|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|Transfer
Finding|Idea or Concept|Impression|3462,3470|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|Transfer
Procedure|Health Care Activity|Impression|3462,3470|false|false|false|C4706767|Transfer (immobility management)|Transfer
Event|Activity|Impression|3517,3524|false|false|false|C1706079||arrival
Event|Event|Impression|3517,3524|false|false|false|||arrival
Finding|Functional Concept|Impression|3517,3524|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Anatomy|Anatomical Structure|Impression|3532,3537|false|false|false|C3714591|Floor (anatomic)|floor
Finding|Body Substance|Impression|3539,3546|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Impression|3539,3546|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Impression|3539,3546|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Impression|3547,3555|false|false|false|||recounts
Event|Event|Impression|3560,3567|false|false|false|||history
Finding|Conceptual Entity|Impression|3560,3567|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Impression|3560,3567|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Impression|3560,3567|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Idea or Concept|Impression|3571,3576|false|false|false|C1552828|Table Frame - above|above
Event|Event|Impression|3583,3587|false|false|false|||says
Event|Event|Impression|3597,3602|false|false|false|||feels
Event|Event|Impression|3603,3611|true|false|false|||improved
Finding|Finding|Impression|3603,3611|true|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Finding|Intellectual Product|Impression|3603,3611|true|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Procedure|Health Care Activity|Impression|3612,3627|true|false|false|C0001758|Aftercare|after treatment
Event|Event|Impression|3618,3627|true|false|false|||treatment
Finding|Conceptual Entity|Impression|3618,3627|true|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Impression|3618,3627|true|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Impression|3618,3627|true|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Impression|3618,3627|true|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Event|Event|Impression|3642,3649|true|false|false|||ongoing
Finding|Idea or Concept|Impression|3642,3649|true|false|false|C0549178|Continuous|ongoing
Event|Event|Impression|3650,3653|true|false|false|||SOB
Finding|Sign or Symptom|Impression|3650,3653|true|false|false|C0013404|Dyspnea|SOB
Anatomy|Body Space or Junction|Impression|3667,3670|false|false|false|C0262327|rostral sulcus|ROS
Drug|Biologically Active Substance|Impression|3667,3670|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Element, Ion, or Isotope|Impression|3667,3670|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Organic Chemical|Impression|3667,3670|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Pharmacologic Substance|Impression|3667,3670|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Event|Event|Impression|3667,3670|false|false|false|||ROS
Finding|Gene or Genome|Impression|3667,3670|false|false|false|C0812281;C1709820|ROS1 gene;ROS1 wt Allele|ROS
Procedure|Health Care Activity|Impression|3667,3670|false|false|false|C0489633|Review of systems (procedure)|ROS
Event|Event|Impression|3684,3692|false|false|false|||NEGATIVE
Finding|Classification|Impression|3684,3692|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Finding|Finding|Impression|3684,3692|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Lab|Laboratory or Test Result|Impression|3684,3692|false|false|false|C5237010|Expression Negative|NEGATIVE
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|3719,3727|false|false|false|C0018787|Heart|Coronary
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|3719,3734|false|false|false|C0205042|Coronary artery|Coronary artery
Disorder|Disease or Syndrome|Past Medical History|3719,3742|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|Coronary artery disease
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|3728,3734|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|Past Medical History|3728,3734|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Disorder|Disease or Syndrome|Past Medical History|3728,3742|false|false|false|C0852949|Arteriopathic disease|artery disease
Disorder|Disease or Syndrome|Past Medical History|3735,3742|false|false|false|C0012634|Disease|disease
Event|Event|Past Medical History|3735,3742|false|false|false|||disease
Disorder|Disease or Syndrome|Past Medical History|3743,3770|false|false|false|C0085096|Peripheral Vascular Diseases|Peripheral vascular disease
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|3754,3762|false|false|false|C0005847|Blood Vessel|vascular
Disorder|Disease or Syndrome|Past Medical History|3754,3770|false|false|false|C0042373|Vascular Diseases|vascular disease
Disorder|Disease or Syndrome|Past Medical History|3763,3770|false|false|false|C0012634|Disease|disease
Event|Event|Past Medical History|3763,3770|false|false|false|||disease
Finding|Gene or Genome|Past Medical History|3771,3775|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|Type
Finding|Intellectual Product|Past Medical History|3771,3775|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|Type
Disorder|Disease or Syndrome|Past Medical History|3771,3787|false|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|Type II Diabetes
Disorder|Disease or Syndrome|Past Medical History|3771,3796|false|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|Type II Diabetes Mellitus
Disorder|Disease or Syndrome|Past Medical History|3779,3787|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|Diabetes
Event|Event|Past Medical History|3779,3787|false|false|false|||Diabetes
Disorder|Disease or Syndrome|Past Medical History|3779,3796|false|false|false|C0011849|Diabetes Mellitus|Diabetes Mellitus
Finding|Finding|Past Medical History|3801,3809|false|false|false|C0241863|Diabetic|diabetic
Disorder|Disease or Syndrome|Past Medical History|3801,3821|false|false|false|C0011884|Diabetic Retinopathy|diabetic retinopathy
Disorder|Disease or Syndrome|Past Medical History|3810,3821|false|false|false|C0035309|Retinal Diseases|retinopathy
Event|Event|Past Medical History|3810,3821|false|false|false|||retinopathy
Disorder|Disease or Syndrome|Past Medical History|3822,3829|false|false|false|C0028754|Obesity|Obesity
Event|Event|Past Medical History|3822,3829|false|false|false|||Obesity
Finding|Finding|Past Medical History|3822,3829|false|false|false|C4759928|BODY MASS INDEX QUANTITATIVE TRAIT LOCUS 20|Obesity
Disorder|Disease or Syndrome|Past Medical History|3830,3840|false|false|false|C0014852|Esophageal Diseases|Esophageal
Disorder|Disease or Syndrome|Past Medical History|3830,3845|false|false|false|C0267081|Terminal esophageal web|Esophageal ring
Drug|Biomedical or Dental Material|Past Medical History|3841,3845|false|false|false|C1882953|Ring Dosage Form|ring
Event|Event|Past Medical History|3841,3845|false|false|false|||ring
Disorder|Disease or Syndrome|Past Medical History|3846,3858|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|Past Medical History|3846,3858|false|false|false|||Hypertension
Disorder|Disease or Syndrome|Past Medical History|3859,3871|false|false|false|C0242339|Dyslipidemias|Dyslipidemia
Event|Event|Past Medical History|3859,3871|false|false|false|||Dyslipidemia
Disorder|Disease or Syndrome|Past Medical History|3893,3902|false|false|false|C0751438|Posterior pituitary disease|posterior
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|3903,3909|false|false|false|C0040184|Bone structure of tibia|tibial
Disorder|Disease or Syndrome|Past Medical History|3910,3914|false|false|false|C0151950|Deep thrombophlebitis|DVTs
Event|Event|Past Medical History|3910,3914|false|false|false|||DVTs
Finding|Finding|Past Medical History|3934,3940|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Past Medical History|3934,3940|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|Past Medical History|3946,3949|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Event|Event|Past Medical History|3946,3949|false|false|false|||CKD
Attribute|Clinical Attribute|Past Medical History|3950,3955|false|false|false|C1300072|Tumor stage|Stage
Finding|Intellectual Product|Past Medical History|3950,3958|false|false|false|C0441772|Stage level 4|Stage IV
Event|Event|Past Medical History|3956,3958|false|false|false|||IV
Disorder|Disease or Syndrome|Past Medical History|3966,3969|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|Past Medical History|3966,3969|false|false|false|||HTN
Disorder|Neoplastic Process|Past Medical History|3971,3980|false|false|false|C0027627|Neoplasm Metastasis|secondary
Event|Event|Past Medical History|3971,3980|false|false|false|||secondary
Finding|Functional Concept|Past Medical History|3971,3980|false|false|false|C1522484|metastatic qualifier|secondary
Disorder|Disease or Syndrome|Past Medical History|3971,4000|false|false|false|C0020503|Hyperparathyroidism, Secondary|secondary hyperparathyroidism
Disorder|Disease or Syndrome|Past Medical History|3981,4000|false|false|false|C0020502|Hyperparathyroidism|hyperparathyroidism
Event|Event|Past Medical History|3981,4000|false|false|false|||hyperparathyroidism
Disorder|Disease or Syndrome|Past Medical History|4001,4007|false|false|false|C0002871|Anemia|Anemia
Event|Event|Past Medical History|4001,4007|false|false|false|||Anemia
Disorder|Disease or Syndrome|Past Medical History|4008,4012|false|false|false|C0018099|Gout|Gout
Event|Event|Past Medical History|4008,4012|false|false|false|||Gout
Event|Activity|Family Medical History|4066,4070|false|false|false|C1947906|Sorting|sort
Event|Event|Family Medical History|4066,4070|false|false|false|||sort
Finding|Cell Function|Family Medical History|4066,4070|false|false|false|C0237886;C0700314|Sorting (Cognition);Sorting - Cell Movement|sort
Finding|Mental Process|Family Medical History|4066,4070|false|false|false|C0237886;C0700314|Sorting (Cognition);Sorting - Cell Movement|sort
Disorder|Neoplastic Process|Family Medical History|4074,4080|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Family Medical History|4074,4080|false|false|false|||cancer
Finding|Conceptual Entity|Family Medical History|4082,4088|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|Family Medical History|4082,4088|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Event|Event|Family Medical History|4089,4093|false|false|false|||died
Anatomy|Body Location or Region|Family Medical History|4113,4117|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|4113,4117|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Family Medical History|4113,4117|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Family Medical History|4113,4117|false|false|false|C0740941|Lung Problem|lung
Disorder|Disease or Syndrome|Family Medical History|4113,4125|false|false|false|C0024115|Lung diseases|lung disease
Disorder|Disease or Syndrome|Family Medical History|4118,4125|false|false|false|C0012634|Disease|disease
Event|Event|Family Medical History|4118,4125|false|false|false|||disease
Finding|Idea or Concept|Family Medical History|4127,4133|false|false|false|C1546508|Relationship - Mother|Mother
Event|Event|Family Medical History|4134,4138|false|false|false|||died
Drug|Amino Acid, Peptide, or Protein|Family Medical History|4160,4167|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Immunologic Factor|Family Medical History|4160,4167|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Pharmacologic Substance|Family Medical History|4160,4167|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Event|Event|Family Medical History|4160,4167|false|false|false|||unknown
Finding|Finding|Family Medical History|4160,4167|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Functional Concept|Family Medical History|4160,4167|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Idea or Concept|Family Medical History|4160,4167|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Intellectual Product|Family Medical History|4160,4167|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Event|Event|Family Medical History|4168,4173|false|false|false|||cause
Finding|Conceptual Entity|Family Medical History|4168,4173|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Finding|Functional Concept|Family Medical History|4168,4173|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Disorder|Disease or Syndrome|Family Medical History|4185,4188|true|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Family Medical History|4185,4188|true|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Family Medical History|4185,4188|true|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Family Medical History|4185,4188|true|false|false|||CAD
Finding|Gene or Genome|Family Medical History|4185,4188|true|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Family Medical History|4185,4188|true|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Family Medical History|4185,4188|true|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Family Medical History|4185,4188|true|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Finding|Pathologic Function|Family Medical History|4192,4212|true|false|false|C0085298|Sudden Cardiac Death|sudden cardiac death
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|4199,4206|true|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|Family Medical History|4199,4206|true|false|false|C1314974|Cardiac attachment|cardiac
Finding|Pathologic Function|Family Medical History|4199,4212|true|false|false|C0376297|Cardiac Death|cardiac death
Event|Event|Family Medical History|4207,4212|true|false|false|||death
Finding|Finding|Family Medical History|4207,4212|true|false|false|C0011065;C1306577;C1546949|Cessation of life;Death (finding);Event Consequence - Death|death
Finding|Idea or Concept|Family Medical History|4207,4212|true|false|false|C0011065;C1306577;C1546949|Cessation of life;Death (finding);Event Consequence - Death|death
Finding|Organism Function|Family Medical History|4207,4212|true|false|false|C0011065;C1306577;C1546949|Cessation of life;Death (finding);Event Consequence - Death|death
Event|Event|Family Medical History|4229,4236|true|false|false|||history
Finding|Conceptual Entity|Family Medical History|4229,4236|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|4229,4236|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Family Medical History|4229,4236|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|4229,4239|true|false|false|C0262926|Medical History|history of
Disorder|Neoplastic Process|Family Medical History|4241,4247|true|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Family Medical History|4241,4247|true|false|false|||cancer
Procedure|Health Care Activity|General Exam|4299,4308|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|General Exam|4309,4317|false|false|false|||PHYSICAL
Finding|Finding|General Exam|4309,4317|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|General Exam|4309,4317|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|General Exam|4309,4317|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|General Exam|4309,4322|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|General Exam|4309,4322|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Event|Event|General Exam|4318,4322|false|false|false|||EXAM
Finding|Functional Concept|General Exam|4318,4322|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|4318,4322|false|false|false|C0582103|Medical Examination|EXAM
Event|Event|General Exam|4385,4392|false|false|false|||GENERAL
Finding|Classification|General Exam|4385,4392|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|General Exam|4385,4392|false|false|false|C3812897|General medical service|GENERAL
Event|Event|General Exam|4394,4402|false|false|false|||Pleasant
Finding|Mental Process|General Exam|4394,4402|false|false|false|C2987187|Pleasant|Pleasant
Attribute|Clinical Attribute|General Exam|4444,4447|false|false|false|C1114365||age
Drug|Biologically Active Substance|General Exam|4444,4447|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|General Exam|4444,4447|false|false|false|C0162574|Glycation End Products, Advanced|age
Event|Event|General Exam|4444,4447|false|false|false|||age
Event|Event|General Exam|4449,4455|false|false|false|||taking
Attribute|Clinical Attribute|General Exam|4456,4460|false|false|false|C4318566|Deep Resection Margin|deep
Event|Event|General Exam|4461,4468|false|false|false|||breaths
Finding|Body Substance|General Exam|4461,4468|false|false|false|C0225386|Breath|breaths
Event|Event|General Exam|4475,4483|false|false|false|||speaking
Anatomy|Body Location or Region|General Exam|4486,4491|false|false|false|C1512338|HEENT|HEENT
Event|Event|General Exam|4493,4497|false|false|false|||EOMI
Event|Event|General Exam|4499,4504|false|false|false|||PERRL
Finding|Finding|General Exam|4499,4504|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Finding|Finding|General Exam|4506,4515|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|General Exam|4516,4522|false|false|false|C0036410|Sclera|sclera
Disorder|Disease or Syndrome|General Exam|4516,4522|false|false|false|C0036412|Scleral Diseases|sclera
Event|Event|General Exam|4516,4522|false|false|false|||sclera
Procedure|Health Care Activity|General Exam|4516,4522|false|false|false|C2228481|examination of sclera|sclera
Anatomy|Body Part, Organ, or Organ Component|General Exam|4529,4540|false|false|false|C0009758;C0229274|Structure of palpebral conjunctiva;conjunctiva|conjunctiva
Disorder|Disease or Syndrome|General Exam|4529,4540|false|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|conjunctiva
Disorder|Neoplastic Process|General Exam|4529,4540|false|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|conjunctiva
Event|Event|General Exam|4529,4540|false|false|false|||conjunctiva
Finding|Body Substance|General Exam|4529,4540|false|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|conjunctiva
Finding|Intellectual Product|General Exam|4529,4540|false|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|conjunctiva
Procedure|Health Care Activity|General Exam|4529,4540|false|false|false|C0872390;C2228431|Procedure on conjunctiva;examination of conjunctiva|conjunctiva
Anatomy|Body Part, Organ, or Organ Component|General Exam|4542,4545|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|General Exam|4542,4545|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Location or Region|General Exam|4549,4553|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|General Exam|4549,4553|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|General Exam|4549,4553|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|General Exam|4555,4558|false|false|false|||JVD
Finding|Finding|General Exam|4555,4558|false|false|false|C0425687|Jugular venous engorgement|JVD
Anatomy|Body Part, Organ, or Organ Component|General Exam|4567,4572|false|false|false|C0018787;C4037974|Chest>Heart;Heart|HEART
Disorder|Neoplastic Process|General Exam|4567,4572|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|HEART
Event|Event|General Exam|4567,4572|false|false|false|||HEART
Finding|Sign or Symptom|General Exam|4567,4572|false|false|false|C0795691|HEART PROBLEM|HEART
Event|Event|General Exam|4574,4577|true|false|false|||RRR
Event|Event|General Exam|4589,4596|true|false|false|||murmurs
Finding|Finding|General Exam|4589,4596|true|false|false|C0018808|Heart murmur|murmurs
Event|Event|General Exam|4598,4605|true|false|false|||gallops
Event|Event|General Exam|4610,4614|true|false|false|||rubs
Finding|Finding|General Exam|4610,4614|true|false|false|C0232267|Pericardial friction rub|rubs
Anatomy|Body Part, Organ, or Organ Component|General Exam|4618,4623|false|false|false|C0024109|Lung|LUNGS
Drug|Organic Chemical|General Exam|4625,4629|true|false|false|C0951233|cetrimonium bromide|CTAB
Event|Event|General Exam|4625,4629|true|false|false|||CTAB
Event|Event|General Exam|4634,4641|true|false|false|||wheezes
Finding|Sign or Symptom|General Exam|4634,4641|true|false|false|C0043144|Wheezing|wheezes
Anatomy|Body Location or Region|General Exam|4644,4651|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|General Exam|4644,4651|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|General Exam|4644,4651|false|false|false|||ABDOMEN
Finding|Finding|General Exam|4644,4651|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|General Exam|4653,4658|false|false|false|C0028754|Obesity|Obese
Event|Event|General Exam|4653,4658|false|false|false|||Obese
Finding|Finding|General Exam|4653,4666|false|false|false|C0426650|Obese abdomen|Obese abdomen
Anatomy|Body Location or Region|General Exam|4659,4666|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|General Exam|4659,4666|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Event|Event|General Exam|4659,4666|false|false|false|||abdomen
Finding|Finding|General Exam|4659,4666|false|false|false|C0941288|Abdomen problem|abdomen
Event|Event|General Exam|4709,4718|true|false|false|||nontender
Event|Event|General Exam|4748,4756|true|false|false|||guarding
Finding|Finding|General Exam|4748,4756|true|false|false|C0427198|Protective muscle spasm|guarding
Event|Event|General Exam|4758,4760|true|false|false|||no
Event|Event|General Exam|4761,4779|true|false|false|||hepatosplenomegaly
Finding|Sign or Symptom|General Exam|4761,4779|true|false|false|C0019214|Hepatosplenomegaly|hepatosplenomegaly
Anatomy|Body Part, Organ, or Organ Component|General Exam|4783,4794|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Event|Event|General Exam|4799,4807|true|false|false|||cyanosis
Finding|Sign or Symptom|General Exam|4799,4807|true|false|false|C0010520|Cyanosis|cyanosis
Disorder|Anatomical Abnormality|General Exam|4809,4817|true|false|false|C0149651|Clubbing|clubbing
Event|Event|General Exam|4809,4817|true|false|false|||clubbing
Attribute|Clinical Attribute|General Exam|4822,4827|true|false|false|C1717255||edema
Event|Event|General Exam|4822,4827|true|false|false|||edema
Finding|Pathologic Function|General Exam|4822,4827|true|false|false|C0013604|Edema|edema
Drug|Food|General Exam|4831,4837|false|false|false|C5890763||PULSES
Event|Event|General Exam|4831,4837|false|false|false|||PULSES
Finding|Physiologic Function|General Exam|4831,4837|false|false|false|C0391850|Physiologic pulse|PULSES
Procedure|Health Care Activity|General Exam|4831,4837|false|false|false|C0034107|Pulse taking|PULSES
Finding|Conceptual Entity|General Exam|4842,4848|false|false|false|C0442038;C0920847|Circumpennate;Radial|radial
Drug|Food|General Exam|4849,4855|false|false|false|C5890763||pulses
Event|Event|General Exam|4849,4855|false|false|false|||pulses
Finding|Physiologic Function|General Exam|4849,4855|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|4849,4855|false|false|false|C0034107|Pulse taking|pulses
Event|Event|General Exam|4885,4891|false|false|false|||moving
Anatomy|Body Part, Organ, or Organ Component|General Exam|4898,4909|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Drug|Organic Chemical|General Exam|4915,4922|false|false|false|C1995603|PURPOSE (pharmacologic preparation)|purpose
Drug|Pharmacologic Substance|General Exam|4915,4922|false|false|false|C1995603|PURPOSE (pharmacologic preparation)|purpose
Event|Event|General Exam|4915,4922|false|false|false|||purpose
Finding|Functional Concept|General Exam|4915,4922|false|false|false|C1285529|Purpose|purpose
Anatomy|Body System|General Exam|4926,4930|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|General Exam|4926,4930|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|General Exam|4926,4930|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|General Exam|4926,4930|false|false|false|||SKIN
Finding|Body Substance|General Exam|4926,4930|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|General Exam|4926,4930|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Event|Event|General Exam|4932,4936|true|false|false|||Warm
Finding|Finding|General Exam|4932,4936|true|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|4932,4936|true|false|false|C0687712|warming process|Warm
Finding|Finding|General Exam|4941,4945|true|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|4946,4954|true|false|false|||perfused
Disorder|Injury or Poisoning|General Exam|4959,4971|true|false|false|C0015256|Excoriation|excoriations
Event|Event|General Exam|4959,4971|true|false|false|||excoriations
Event|Event|General Exam|4975,4982|true|false|false|||lesions
Finding|Finding|General Exam|4975,4982|true|false|false|C0221198|Lesion|lesions
Event|Event|General Exam|4987,4993|true|false|false|||rashes
Finding|Sign or Symptom|General Exam|4987,4993|true|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Finding|Body Substance|General Exam|5030,5039|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|5030,5039|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|5030,5039|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|5030,5039|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|General Exam|5040,5048|false|false|false|||PHYSICAL
Finding|Finding|General Exam|5040,5048|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|General Exam|5040,5048|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|General Exam|5040,5048|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|General Exam|5040,5053|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|General Exam|5040,5053|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Event|Event|General Exam|5049,5053|false|false|false|||EXAM
Finding|Functional Concept|General Exam|5049,5053|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|5049,5053|false|false|false|C0582103|Medical Examination|EXAM
Event|Event|General Exam|5124,5127|false|false|false|||GEN
Finding|Classification|General Exam|5124,5127|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|GEN
Finding|Gene or Genome|General Exam|5124,5127|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|GEN
Finding|Finding|General Exam|5129,5133|false|false|false|C5575035|Well (answer to question)|Well
Event|Event|General Exam|5134,5143|false|false|false|||appearing
Disorder|Disease or Syndrome|General Exam|5147,5150|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|5147,5150|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|5147,5150|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|5147,5150|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|5147,5150|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|General Exam|5147,5150|false|false|false|||NAD
Finding|Finding|General Exam|5147,5150|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|General Exam|5151,5155|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|General Exam|5151,5155|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|General Exam|5151,5155|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|General Exam|5161,5164|true|false|false|||JVD
Finding|Finding|General Exam|5161,5164|true|false|false|C0425687|Jugular venous engorgement|JVD
Event|Event|General Exam|5165,5176|true|false|false|||appreciated
Event|Event|General Exam|5181,5184|true|false|false|||RRR
Anatomy|Body Part, Organ, or Organ Component|General Exam|5198,5205|true|false|false|C0007272|Carotid Arteries|carotid
Finding|Finding|General Exam|5198,5212|true|false|false|C0007280|Carotid bruit|carotid bruits
Event|Event|General Exam|5206,5212|true|false|false|||bruits
Finding|Finding|General Exam|5206,5212|true|false|false|C0006318|Bruit|bruits
Event|Event|General Exam|5213,5224|true|false|false|||appreciated
Event|Event|General Exam|5225,5229|true|false|false|||PULM
Procedure|Health Care Activity|General Exam|5225,5229|true|false|false|C1315068|Pulmonary ventilator management|PULM
Drug|Organic Chemical|General Exam|5231,5235|true|false|false|C0951233|cetrimonium bromide|CTAB
Event|Event|General Exam|5231,5235|true|false|false|||CTAB
Event|Event|General Exam|5239,5246|true|false|false|||wheezes
Finding|Sign or Symptom|General Exam|5239,5246|true|false|false|C0043144|Wheezing|wheezes
Event|Event|General Exam|5248,5253|true|false|false|||rales
Finding|Finding|General Exam|5248,5253|true|false|false|C0034642;C0240859|Basilar Rales;Rales|rales
Event|Event|General Exam|5258,5266|true|false|false|||crackles
Finding|Finding|General Exam|5258,5266|true|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Finding|Conceptual Entity|General Exam|5269,5278|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|Symmetric
Finding|Finding|General Exam|5269,5278|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|Symmetric
Disorder|Congenital Abnormality|General Exam|5289,5292|false|false|false|C0015306|Hereditary Multiple Exostoses|EXT
Event|Event|General Exam|5289,5292|false|false|false|||EXT
Finding|Gene or Genome|General Exam|5289,5292|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|EXT
Finding|Finding|General Exam|5294,5298|true|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|General Exam|5294,5298|true|false|false|C0687712|warming process|warm
Finding|Finding|General Exam|5299,5303|true|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|5304,5312|true|false|false|||perfused
Finding|Functional Concept|General Exam|5317,5324|true|false|false|C0205323|Pitting|pitting
Finding|Finding|General Exam|5317,5330|true|false|false|C0333243|Pitting edema|pitting edema
Attribute|Clinical Attribute|General Exam|5325,5330|true|false|false|C1717255||edema
Event|Event|General Exam|5325,5330|true|false|false|||edema
Finding|Pathologic Function|General Exam|5325,5330|true|false|false|C0013604|Edema|edema
Procedure|Health Care Activity|General Exam|5385,5394|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|General Exam|5395,5399|false|false|false|||LABS
Lab|Laboratory or Test Result|General Exam|5395,5399|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|General Exam|5443,5448|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|5443,5448|false|false|false|||BLOOD
Finding|Body Substance|General Exam|5443,5448|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|5449,5452|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|5457,5460|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|5457,5460|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|5457,5460|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|5467,5470|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|5467,5470|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|5467,5470|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|5467,5470|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|5476,5479|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|5476,5479|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|5487,5490|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|5487,5490|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|5487,5490|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|5487,5490|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|5487,5490|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|5494,5497|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|5494,5497|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|5494,5497|false|false|false|||MCH
Finding|Gene or Genome|General Exam|5494,5497|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|5494,5497|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|5494,5497|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|5503,5507|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|5503,5507|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|5534,5537|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|5554,5559|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|5554,5559|false|false|false|||BLOOD
Finding|Body Substance|General Exam|5554,5559|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Event|General Exam|5572,5578|false|false|false|||Lymphs
Finding|Body Substance|General Exam|5572,5578|false|false|false|C0024202|Lymph|Lymphs
Drug|Antibiotic|General Exam|5585,5590|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|General Exam|5585,5590|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|General Exam|5585,5590|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|General Exam|5597,5600|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Event|Event|General Exam|5597,5600|false|false|false|||Eos
Finding|Gene or Genome|General Exam|5597,5600|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|General Exam|5699,5704|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|5699,5704|false|false|false|||BLOOD
Finding|Body Substance|General Exam|5699,5704|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|5709,5712|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|General Exam|5709,5712|false|false|false|||PTT
Procedure|Laboratory Procedure|General Exam|5709,5712|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|General Exam|5734,5739|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|5734,5739|false|false|false|||BLOOD
Finding|Body Substance|General Exam|5734,5739|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|5734,5747|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|5734,5747|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|5734,5747|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|5740,5747|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|5740,5747|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|5740,5747|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|5740,5747|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|5740,5747|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|5740,5747|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|5795,5799|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|5795,5799|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|5795,5799|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|5825,5830|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|5825,5830|false|false|false|||BLOOD
Finding|Body Substance|General Exam|5825,5830|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|5831,5837|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Drug|Hormone|General Exam|5831,5837|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Disorder|Disease or Syndrome|General Exam|5856,5861|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|5856,5861|false|false|false|||BLOOD
Finding|Body Substance|General Exam|5856,5861|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|General Exam|5888,5893|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|5888,5893|false|false|false|||BLOOD
Finding|Body Substance|General Exam|5888,5893|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|5894,5899|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|General Exam|5894,5899|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|General Exam|5894,5899|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|General Exam|5894,5899|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Drug|Pharmacologic Substance|General Exam|5897,5901|false|false|false|C4722362|MB-6|MB-6
Disorder|Disease or Syndrome|General Exam|5928,5933|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|5928,5933|false|false|false|||BLOOD
Finding|Body Substance|General Exam|5928,5933|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|5934,5939|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|General Exam|5934,5939|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|General Exam|5934,5939|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|General Exam|5934,5939|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Drug|Organic Chemical|General Exam|5937,5941|false|false|false|C0602256|MB 5|MB-5
Disorder|Disease or Syndrome|General Exam|5968,5973|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|5968,5973|false|false|false|||BLOOD
Finding|Body Substance|General Exam|5968,5973|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|5968,5981|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|General Exam|5974,5981|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|5974,5981|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|5974,5981|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|5974,5981|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|5974,5981|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|General Exam|5974,5981|false|false|false|||Calcium
Finding|Physiologic Function|General Exam|5974,5981|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|5974,5981|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|General Exam|6014,6019|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|6014,6019|false|false|false|||BLOOD
Finding|Body Substance|General Exam|6014,6019|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Event|General Exam|6024,6027|false|false|false|||pO2
Finding|Classification|General Exam|6024,6027|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|pO2
Finding|Molecular Function|General Exam|6024,6027|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|pO2
Procedure|Laboratory Procedure|General Exam|6024,6027|false|false|false|C1283004|PO2 measurement|pO2
Lab|Laboratory or Test Result|General Exam|6032,6036|false|false|false|C0391839|Carbon dioxide, partial pressure|pCO2
Procedure|Laboratory Procedure|General Exam|6032,6036|false|false|false|C0201931|Carbon dioxide measurement, partial pressure|pCO2
Anatomy|Body Location or Region|General Exam|6061,6065|false|false|false|C2987514|Anatomical base|Base
Drug|Biomedical or Dental Material|General Exam|6061,6065|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Drug|Chemical Viewed Functionally|General Exam|6061,6065|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|6061,6065|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Finding|Gene or Genome|General Exam|6061,6065|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|Base
Finding|Idea or Concept|General Exam|6061,6065|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|Base
Event|Event|General Exam|6106,6113|false|false|false|||IMAGING
Finding|Finding|General Exam|6106,6113|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|General Exam|6106,6113|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Event|Event|General Exam|6145,6148|false|false|false|||TTE
Procedure|Diagnostic Procedure|General Exam|6145,6148|false|false|false|C0430462|Transthoracic echocardiography|TTE
Finding|Functional Concept|General Exam|6158,6162|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Finding|General Exam|6158,6176|false|false|false|C2059558||left atrial volume
Anatomy|Body Part, Organ, or Organ Component|General Exam|6163,6169|false|false|false|C0018792|Heart Atrium|atrial
Finding|Intellectual Product|General Exam|6170,6176|false|false|false|C1705102|Volume (publication)|volume
Event|Event|General Exam|6177,6182|false|false|false|||index
Finding|Idea or Concept|General Exam|6177,6182|false|false|false|C0600653;C0918012;C1552854|Html Link Type - index;Index;Indexes|index
Finding|Intellectual Product|General Exam|6177,6182|false|false|false|C0600653;C0918012;C1552854|Html Link Type - index;Index;Indexes|index
Event|Event|General Exam|6193,6202|false|false|false|||increased
Finding|Functional Concept|General Exam|6219,6224|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Attribute|Clinical Attribute|General Exam|6219,6240|false|false|false|C0456165;C4050168|Right atrial pressure|right atrial pressure
Anatomy|Body Part, Organ, or Organ Component|General Exam|6225,6231|false|false|false|C0018792|Heart Atrium|atrial
Finding|Finding|General Exam|6225,6240|false|false|false|C0428877|Atrial Pressure|atrial pressure
Event|Event|General Exam|6232,6240|false|false|false|||pressure
Finding|Finding|General Exam|6232,6240|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|General Exam|6232,6240|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|General Exam|6232,6240|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|General Exam|6232,6240|false|false|false|C0033095||pressure
Finding|Functional Concept|General Exam|6254,6258|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|General Exam|6260,6271|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Part, Organ, or Organ Component|General Exam|6260,6276|false|false|false|C0507618|Wall of ventricle|ventricular wall
Event|Event|General Exam|6277,6288|false|false|false|||thicknesses
Anatomy|Body Space or Junction|General Exam|6293,6299|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|General Exam|6293,6299|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|General Exam|6293,6299|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Event|Event|General Exam|6300,6304|false|false|false|||size
Event|Event|General Exam|6309,6315|false|false|false|||normal
Finding|Intellectual Product|General Exam|6327,6331|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Functional Concept|General Exam|6341,6345|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Disorder|Disease or Syndrome|General Exam|6341,6378|false|false|false|C1277187|Left ventricular systolic dysfunction|left ventricular systolic dysfunction
Anatomy|Body Part, Organ, or Organ Component|General Exam|6346,6357|false|false|false|C0018827|Heart Ventricle|ventricular
Finding|Organ or Tissue Function|General Exam|6358,6366|false|false|false|C0039155|Systole|systolic
Finding|Pathologic Function|General Exam|6358,6378|false|false|false|C0749225|Systolic dysfunction|systolic dysfunction
Disorder|Disease or Syndrome|General Exam|6367,6378|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Event|Event|General Exam|6367,6378|false|false|false|||dysfunction
Finding|Conceptual Entity|General Exam|6367,6378|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|General Exam|6367,6378|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|General Exam|6367,6378|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Event|Event|General Exam|6391,6403|false|false|false|||inferoseptal
Event|Event|General Exam|6405,6413|false|false|false|||inferior
Finding|Social Behavior|General Exam|6405,6413|false|false|false|C0678975|inferiority|inferior
Finding|Finding|General Exam|6432,6436|false|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|6445,6453|false|false|false|||inferior
Finding|Social Behavior|General Exam|6445,6453|false|false|false|C0678975|inferiority|inferior
Attribute|Clinical Attribute|General Exam|6467,6478|false|false|false|C1980023|Wall motion|wall motion
Phenomenon|Natural Phenomenon or Process|General Exam|6472,6478|false|false|false|C0026597|Motion|motion
Disorder|Congenital Abnormality|General Exam|6479,6492|false|false|false|C0000768|Congenital Abnormality|abnormalities
Event|Event|General Exam|6479,6492|false|false|false|||abnormalities
Finding|Functional Concept|General Exam|6479,6492|false|false|false|C0000769|teratologic|abnormalities
Procedure|Diagnostic Procedure|General Exam|6494,6501|false|false|false|C0554756|Doppler studies|Doppler
Event|Event|General Exam|6503,6513|false|false|false|||parameters
Finding|Finding|General Exam|6503,6513|false|false|false|C0449381|Observation parameter|parameters
Event|Event|General Exam|6523,6533|false|false|false|||consistent
Finding|Idea or Concept|General Exam|6523,6533|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|General Exam|6523,6538|false|false|false|C0332290|Consistent with|consistent with
Finding|Classification|General Exam|6534,6544|false|false|false|C0441800|Grade|with Grade
Finding|Classification|General Exam|6539,6544|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|Grade
Finding|Finding|General Exam|6539,6544|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|Grade
Finding|Classification|General Exam|6539,6547|false|false|false|C0441802;C0475270;C1522446;C4049999|Clavien-Dindo Grade II;Disease Grade 2;G2 stage (tumor staging);Grade two rank|Grade II
Finding|Intellectual Product|General Exam|6539,6547|false|false|false|C0441802;C0475270;C1522446;C4049999|Clavien-Dindo Grade II;Disease Grade 2;G2 stage (tumor staging);Grade two rank|Grade II
Finding|Finding|General Exam|6549,6557|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|General Exam|6549,6557|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Functional Concept|General Exam|6559,6563|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|General Exam|6565,6576|false|false|false|C0018827|Heart Ventricle|ventricular
Attribute|Clinical Attribute|General Exam|6577,6586|false|false|false|C0012000|Diastole|diastolic
Finding|Pathologic Function|General Exam|6577,6598|false|false|false|C0520863|Diastolic dysfunction|diastolic dysfunction
Disorder|Disease or Syndrome|General Exam|6587,6598|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Event|Event|General Exam|6587,6598|false|false|false|||dysfunction
Finding|Conceptual Entity|General Exam|6587,6598|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|General Exam|6587,6598|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|General Exam|6587,6598|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|General Exam|6600,6605|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Part, Organ, or Organ Component|General Exam|6606,6617|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Part, Organ, or Organ Component|General Exam|6618,6625|false|false|false|C0935616|chamber [body part]|chamber
Event|Event|General Exam|6636,6640|false|false|false|||free
Finding|Functional Concept|General Exam|6636,6640|false|false|false|C0332296|Free of (attribute)|free
Attribute|Clinical Attribute|General Exam|6641,6652|false|false|false|C1980023|Wall motion|wall motion
Event|Event|General Exam|6646,6652|false|false|false|||motion
Phenomenon|Natural Phenomenon or Process|General Exam|6646,6652|false|false|false|C0026597|Motion|motion
Event|Event|General Exam|6657,6663|false|false|false|||normal
Event|Event|General Exam|6669,6678|false|false|false|||diameters
Anatomy|Body Part, Organ, or Organ Component|General Exam|6682,6687|false|false|false|C0003483;C4037978|Aorta;Chest+Abdomen>Aorta|aorta
Procedure|Health Care Activity|General Exam|6682,6687|false|false|false|C0869784|Procedure on aorta|aorta
Anatomy|Body Space or Junction|General Exam|6696,6701|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|General Exam|6696,6701|false|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|General Exam|6696,6701|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|General Exam|6696,6701|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Event|Event|General Exam|6703,6712|false|false|false|||ascending
Finding|Functional Concept|General Exam|6703,6712|false|false|false|C1547175;C1962987|Ascend (action);Sequencing - Ascending|ascending
Anatomy|Body Location or Region|General Exam|6717,6721|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Anatomy|Body Part, Organ, or Organ Component|General Exam|6717,6721|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Anatomy|Body Space or Junction|General Exam|6717,6721|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Finding|Finding|General Exam|6717,6721|false|false|false|C1538146;C4722404|Age-Related Clonal Hematopoiesis;ZBTB8OS gene|arch
Finding|Gene or Genome|General Exam|6717,6721|false|false|false|C1538146;C4722404|Age-Related Clonal Hematopoiesis;ZBTB8OS gene|arch
Event|Event|General Exam|6722,6728|false|false|false|||levels
Event|Event|General Exam|6733,6739|false|false|false|||normal
Anatomy|Body Part, Organ, or Organ Component|General Exam|6745,6751|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|General Exam|6753,6758|false|false|false|C1186983|Anatomical valve|valve
Event|Event|General Exam|6759,6767|false|false|false|||leaflets
Event|Event|General Exam|6783,6792|false|false|false|||thickened
Anatomy|Body Part, Organ, or Organ Component|General Exam|6797,6803|true|false|false|C0003483|Aorta|aortic
Finding|Pathologic Function|General Exam|6797,6812|true|false|false|C0003507|Aortic Valve Stenosis|aortic stenosis
Event|Event|General Exam|6804,6812|true|false|false|||stenosis
Finding|Pathologic Function|General Exam|6804,6812|true|false|false|C1261287|Stenosis|stenosis
Event|Event|General Exam|6821,6828|true|false|false|||present
Finding|Finding|General Exam|6821,6828|true|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|General Exam|6821,6828|true|false|false|C0150312;C0449450|Present;Presentation|present
Anatomy|Body Part, Organ, or Organ Component|General Exam|6842,6848|true|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|General Exam|6842,6854|true|false|false|C0003501;C4533215|Aortic valve structure;Chest>Aortic valve|aortic valve
Disorder|Congenital Abnormality|General Exam|6842,6863|true|false|false|C5193127;C5700069|AORTIC VALVE DISEASE 3;Stenosis of aorta|aortic valve stenosis
Disorder|Disease or Syndrome|General Exam|6842,6863|true|false|false|C5193127;C5700069|AORTIC VALVE DISEASE 3;Stenosis of aorta|aortic valve stenosis
Finding|Pathologic Function|General Exam|6842,6863|true|false|false|C0003507|Aortic Valve Stenosis|aortic valve stenosis
Anatomy|Body Part, Organ, or Organ Component|General Exam|6849,6854|true|false|false|C1186983|Anatomical valve|valve
Event|Event|General Exam|6855,6863|true|false|false|||stenosis
Finding|Pathologic Function|General Exam|6855,6863|true|false|false|C1261287|Stenosis|stenosis
Finding|Functional Concept|General Exam|6865,6870|false|false|false|C1883002|Sequence Chromatogram|Trace
Anatomy|Body Part, Organ, or Organ Component|General Exam|6871,6877|false|false|false|C0003483|Aorta|aortic
Event|Event|General Exam|6879,6892|false|false|false|||regurgitation
Finding|Finding|General Exam|6879,6892|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|General Exam|6879,6892|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|General Exam|6879,6892|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Event|Event|General Exam|6896,6900|false|false|false|||seen
Anatomy|Body Part, Organ, or Organ Component|General Exam|6906,6918|false|false|false|C0026264|Mitral Valve|mitral valve
Anatomy|Body Part, Organ, or Organ Component|General Exam|6913,6918|false|false|false|C1186983|Anatomical valve|valve
Event|Event|General Exam|6919,6927|false|false|false|||leaflets
Finding|Finding|General Exam|6932,6942|false|false|false|C4085643;C5201148;C5962468|Moderate;Moderate Effect;Moderate Response|moderately
Event|Event|General Exam|6944,6953|false|false|false|||thickened
Finding|Intellectual Product|General Exam|6955,6959|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Disorder|Disease or Syndrome|General Exam|6965,6985|false|false|false|C0026266|Mitral Valve Insufficiency|mitral regurgitation
Event|Event|General Exam|6972,6985|false|false|false|||regurgitation
Finding|Finding|General Exam|6972,6985|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|General Exam|6972,6985|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|General Exam|6972,6985|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Event|Event|General Exam|6989,6993|false|false|false|||seen
Anatomy|Body Part, Organ, or Organ Component|General Exam|7010,7015|false|false|false|C1186983|Anatomical valve|valve
Event|Event|General Exam|7016,7024|false|false|false|||leaflets
Event|Event|General Exam|7036,7045|false|false|false|||thickened
Finding|Intellectual Product|General Exam|7056,7060|false|false|false|C1547225|Mild Severity of Illness Code|mild
Anatomy|Body Part, Organ, or Organ Component|General Exam|7061,7070|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|General Exam|7061,7070|false|false|false|C2707265||pulmonary
Finding|Finding|General Exam|7061,7070|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Anatomy|Body Part, Organ, or Organ Component|General Exam|7072,7078|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|General Exam|7072,7078|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Finding|Organ or Tissue Function|General Exam|7079,7087|false|false|false|C0039155|Systole|systolic
Disorder|Disease or Syndrome|General Exam|7079,7100|false|false|false|C0221155|Systolic Hypertension|systolic hypertension
Disorder|Disease or Syndrome|General Exam|7088,7100|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|General Exam|7088,7100|false|false|false|||hypertension
Anatomy|Body Location or Region|General Exam|7114,7125|true|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|General Exam|7114,7125|true|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Disorder|Disease or Syndrome|General Exam|7114,7134|true|false|false|C0031039|Pericardial effusion|pericardial effusion
Finding|Body Substance|General Exam|7114,7134|true|false|false|C1253937|Pericardial effusion body substance|pericardial effusion
Event|Event|General Exam|7126,7134|true|false|false|||effusion
Finding|Body Substance|General Exam|7126,7134|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|General Exam|7126,7134|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|General Exam|7126,7134|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Event|Event|General Exam|7139,7149|false|false|false|||IMPRESSION
Finding|Intellectual Product|General Exam|7139,7149|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|General Exam|7139,7149|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Intellectual Product|General Exam|7156,7160|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Disorder|Disease or Syndrome|General Exam|7170,7193|false|false|false|C1277187|Left ventricular systolic dysfunction|LV systolic dysfunction
Finding|Organ or Tissue Function|General Exam|7173,7181|false|false|false|C0039155|Systole|systolic
Finding|Pathologic Function|General Exam|7173,7193|false|false|false|C0749225|Systolic dysfunction|systolic dysfunction
Disorder|Disease or Syndrome|General Exam|7182,7193|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Event|Event|General Exam|7182,7193|false|false|false|||dysfunction
Finding|Conceptual Entity|General Exam|7182,7193|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|General Exam|7182,7193|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|General Exam|7182,7193|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Finding|General Exam|7199,7226|false|false|false|C0155668|Old myocardial infarction|prior myocardial infarction
Anatomy|Tissue|General Exam|7205,7215|false|false|false|C0027061|Myocardium|myocardial
Attribute|Clinical Attribute|General Exam|7205,7226|false|false|false|C2926063||myocardial infarction
Disorder|Disease or Syndrome|General Exam|7205,7226|false|false|false|C0027051|Myocardial Infarction|myocardial infarction
Event|Event|General Exam|7216,7226|false|false|false|||infarction
Finding|Pathologic Function|General Exam|7216,7226|false|false|false|C0021308|Infarction|infarction
Event|Event|General Exam|7238,7247|false|false|false|||territory
Finding|Classification|General Exam|7254,7259|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|Grade
Finding|Finding|General Exam|7254,7259|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|Grade
Finding|Classification|General Exam|7254,7262|false|false|false|C0441802;C0475270;C1522446;C4049999|Clavien-Dindo Grade II;Disease Grade 2;G2 stage (tumor staging);Grade two rank|Grade II
Finding|Intellectual Product|General Exam|7254,7262|false|false|false|C0441802;C0475270;C1522446;C4049999|Clavien-Dindo Grade II;Disease Grade 2;G2 stage (tumor staging);Grade two rank|Grade II
Disorder|Disease or Syndrome|General Exam|7264,7288|false|false|false|C1273070|Left ventricular diastolic dysfunction|LV diastolic dysfunction
Attribute|Clinical Attribute|General Exam|7267,7276|false|false|false|C0012000|Diastole|diastolic
Finding|Pathologic Function|General Exam|7267,7288|false|false|false|C0520863|Diastolic dysfunction|diastolic dysfunction
Disorder|Disease or Syndrome|General Exam|7277,7288|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Event|Event|General Exam|7277,7288|false|false|false|||dysfunction
Finding|Conceptual Entity|General Exam|7277,7288|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|General Exam|7277,7288|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|General Exam|7277,7288|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Event|Event|General Exam|7315,7320|false|false|false|||study
Finding|Intellectual Product|General Exam|7315,7320|false|false|false|C1705923|Study Object|study
Procedure|Research Activity|General Exam|7315,7320|false|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|study
Event|Event|General Exam|7329,7337|false|false|false|||reviewed
Event|Event|General Exam|7359,7367|false|false|false|||function
Finding|Finding|General Exam|7359,7367|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|General Exam|7359,7367|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|General Exam|7359,7367|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|General Exam|7359,7367|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Event|Event|General Exam|7388,7396|false|false|false|||vigorous
Phenomenon|Natural Phenomenon or Process|General Exam|7413,7419|false|false|false|C0026597|Motion|motion
Disorder|Congenital Abnormality|General Exam|7420,7433|false|false|false|C0000768|Congenital Abnormality|abnormalities
Event|Event|General Exam|7420,7433|false|false|false|||abnormalities
Finding|Functional Concept|General Exam|7420,7433|false|false|false|C0000769|teratologic|abnormalities
Event|Event|General Exam|7464,7473|false|false|false|||territory
Event|Event|General Exam|7478,7481|false|false|false|||CXR
Procedure|Diagnostic Procedure|General Exam|7478,7481|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|General Exam|7482,7484|false|false|false|||PA
Drug|Amino Acid, Peptide, or Protein|General Exam|7487,7490|false|false|false|C1366678;C1433371;C4049852|L-Type Amino Acid Transporter;LAT protein, human;ORC3 protein, human|LAT
Drug|Biologically Active Substance|General Exam|7487,7490|false|false|false|C1366678;C1433371;C4049852|L-Type Amino Acid Transporter;LAT protein, human;ORC3 protein, human|LAT
Drug|Immunologic Factor|General Exam|7487,7490|false|false|false|C1366678;C1433371;C4049852|L-Type Amino Acid Transporter;LAT protein, human;ORC3 protein, human|LAT
Event|Event|General Exam|7487,7490|false|false|false|||LAT
Finding|Gene or Genome|General Exam|7487,7490|false|false|false|C1335085;C1425844;C1705279;C2240043|LAT gene;ORC3 gene;ORC3 wt Allele;SPNS1 gene|LAT
Disorder|Disease or Syndrome|General Exam|7505,7518|true|false|false|C0521530|Lung consolidation|consolidation
Event|Event|General Exam|7505,7518|true|false|false|||consolidation
Anatomy|Body Part, Organ, or Organ Component|General Exam|7522,7531|true|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|General Exam|7522,7531|true|false|false|C2707265||pulmonary
Finding|Finding|General Exam|7522,7531|true|false|false|C4522268|Pulmonary (intended site)|pulmonary
Attribute|Clinical Attribute|General Exam|7533,7538|true|false|false|C1717255||edema
Event|Event|General Exam|7533,7538|true|false|false|||edema
Finding|Pathologic Function|General Exam|7533,7538|true|false|false|C0013604|Edema|edema
Anatomy|Body Location or Region|General Exam|7551,7556|false|false|false|C1548802|Body Site Modifier - Lower|LOWER
Event|Activity|General Exam|7551,7556|false|false|false|C2003888|Lower (action)|LOWER
Anatomy|Body Part, Organ, or Organ Component|General Exam|7551,7566|false|false|false|C0023216|Lower Extremity|LOWER EXTREMITY
Anatomy|Body Part, Organ, or Organ Component|General Exam|7557,7566|false|false|false|C0015385|Limb structure|EXTREMITY
Procedure|Diagnostic Procedure|General Exam|7567,7574|false|false|false|C0554756|Doppler studies|DOPPLER
Procedure|Diagnostic Procedure|General Exam|7567,7585|false|false|false|C0162481|Doppler Ultrasound (procedure)|DOPPLER ULTRASOUND
Event|Event|General Exam|7575,7585|false|false|false|||ULTRASOUND
Finding|Functional Concept|General Exam|7575,7585|false|false|false|C0220934|Ultrasonic|ULTRASOUND
Phenomenon|Natural Phenomenon or Process|General Exam|7575,7585|false|false|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|ULTRASOUND
Procedure|Diagnostic Procedure|General Exam|7575,7585|false|false|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|ULTRASOUND
Event|Event|General Exam|7610,7620|false|false|false|||thrombosis
Finding|Pathologic Function|General Exam|7610,7620|false|false|false|C0040053|Thrombosis|thrombosis
Disorder|Disease or Syndrome|General Exam|7642,7651|false|false|false|C0751438|Posterior pituitary disease|posterior
Anatomy|Body Part, Organ, or Organ Component|General Exam|7652,7658|false|false|false|C0040184|Bone structure of tibia|tibial
Anatomy|Body Part, Organ, or Organ Component|General Exam|7660,7665|false|false|false|C0042449|Veins|veins
Event|Event|General Exam|7660,7665|false|false|false|||veins
Procedure|Therapeutic or Preventive Procedure|General Exam|7660,7665|false|false|false|C0398102|Procedure on vein|veins
Anatomy|Body Location or Region|General Exam|7683,7688|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|7683,7688|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|General Exam|7683,7700|false|false|false|C0023216|Lower Extremity|lower extremities
Anatomy|Body Part, Organ, or Organ Component|General Exam|7689,7700|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Event|Event|General Exam|7724,7733|false|false|false|||unchanged
Finding|Finding|General Exam|7724,7733|false|false|false|C0442739||unchanged
Event|Event|General Exam|7734,7742|false|false|false|||compared
Anatomy|Body Location or Region|General Exam|7756,7761|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|7756,7761|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|General Exam|7756,7771|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|General Exam|7762,7771|false|false|false|C0015385|Limb structure|extremity
Event|Event|General Exam|7772,7782|false|false|false|||ultrasound
Finding|Functional Concept|General Exam|7772,7782|false|false|false|C0220934|Ultrasonic|ultrasound
Phenomenon|Natural Phenomenon or Process|General Exam|7772,7782|false|false|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|ultrasound
Procedure|Diagnostic Procedure|General Exam|7772,7782|false|false|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|ultrasound
Finding|Finding|General Exam|7792,7795|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|General Exam|7792,7795|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Attribute|Clinical Attribute|General Exam|7796,7800|true|false|false|C4318566|Deep Resection Margin|deep
Disorder|Disease or Syndrome|General Exam|7796,7818|true|false|false|C0149871|Deep Vein Thrombosis|deep venous thrombosis
Anatomy|Body Part, Organ, or Organ Component|General Exam|7801,7807|true|false|false|C0042449|Veins|venous
Finding|Finding|General Exam|7801,7818|true|false|false|C0042487;C0517555|Venous Thrombosis;Venous thrombosis after immobility|venous thrombosis
Finding|Pathologic Function|General Exam|7801,7818|true|false|false|C0042487;C0517555|Venous Thrombosis;Venous thrombosis after immobility|venous thrombosis
Event|Event|General Exam|7808,7818|true|false|false|||thrombosis
Finding|Pathologic Function|General Exam|7808,7818|true|false|false|C0040053|Thrombosis|thrombosis
Anatomy|Body Part, Organ, or Organ Component|General Exam|7830,7839|false|false|false|C0015385|Limb structure|extremity
Finding|Functional Concept|General Exam|7845,7850|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Disorder|Anatomical Abnormality|General Exam|7855,7859|false|false|false|C0010709|Cyst|cyst
Event|Event|General Exam|7855,7859|false|false|false|||cyst
Finding|Body Substance|General Exam|7855,7859|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Finding|Intellectual Product|General Exam|7855,7859|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Event|Event|General Exam|7860,7869|false|false|false|||measuring
Event|Event|General Exam|7912,7921|false|false|false|||unchanged
Finding|Finding|General Exam|7912,7921|false|false|false|C0442739||unchanged
Event|Event|General Exam|7983,7995|false|false|false|||MICROBIOLOGY
Finding|Functional Concept|General Exam|7983,7995|false|false|false|C0025953;C1571921;C4049106|Microbiological;Microbiology - Laboratory Class;Microbiology Diagnostic Service Section ID|MICROBIOLOGY
Finding|Intellectual Product|General Exam|7983,7995|false|false|false|C0025953;C1571921;C4049106|Microbiological;Microbiology - Laboratory Class;Microbiology Diagnostic Service Section ID|MICROBIOLOGY
Procedure|Laboratory Procedure|General Exam|7983,7995|false|false|false|C0085672|Microbiology procedure|MICROBIOLOGY
Finding|Body Substance|General Exam|8028,8033|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|8028,8033|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|8028,8033|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Procedure|Laboratory Procedure|General Exam|8028,8041|false|false|false|C0430404|Urine culture|URINE CULTURE
Drug|Biomedical or Dental Material|General Exam|8034,8041|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|General Exam|8034,8041|false|false|false|||CULTURE
Finding|Functional Concept|General Exam|8034,8041|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|General Exam|8034,8041|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|General Exam|8034,8041|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|General Exam|8060,8062|false|false|false|||SP
Disorder|Disease or Syndrome|General Exam|8086,8091|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|8086,8091|false|false|false|||BLOOD
Finding|Body Substance|General Exam|8086,8091|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|8086,8099|false|false|false|C0200949|Blood culture|BLOOD CULTURE
Drug|Biomedical or Dental Material|General Exam|8092,8099|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|General Exam|8092,8099|false|false|false|||CULTURE
Finding|Functional Concept|General Exam|8092,8099|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|General Exam|8092,8099|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|General Exam|8092,8099|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Disorder|Disease or Syndrome|General Exam|8105,8110|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Event|Event|General Exam|8105,8110|false|false|false|||Blood
Finding|Body Substance|General Exam|8105,8110|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Procedure|Laboratory Procedure|General Exam|8105,8118|false|false|false|C0200949|Blood culture|Blood Culture
Drug|Biomedical or Dental Material|General Exam|8111,8118|false|false|false|C1706355|Culture Dose Form|Culture
Event|Event|General Exam|8111,8118|false|false|false|||Culture
Finding|Functional Concept|General Exam|8111,8118|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|Culture
Finding|Idea or Concept|General Exam|8111,8118|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|Culture
Procedure|Laboratory Procedure|General Exam|8111,8118|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|Culture
Finding|Idea or Concept|General Exam|8120,8127|false|false|false|C1691786;C1704475|Pending - Allergy Clinical Status;Pending - referral status|PENDING
Disorder|Disease or Syndrome|General Exam|8130,8135|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|8130,8135|false|false|false|||BLOOD
Finding|Body Substance|General Exam|8130,8135|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|8130,8143|false|false|false|C0200949|Blood culture|BLOOD CULTURE
Drug|Biomedical or Dental Material|General Exam|8136,8143|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|General Exam|8136,8143|false|false|false|||CULTURE
Finding|Functional Concept|General Exam|8136,8143|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|General Exam|8136,8143|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|General Exam|8136,8143|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Disorder|Disease or Syndrome|General Exam|8149,8154|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Event|Event|General Exam|8149,8154|false|false|false|||Blood
Finding|Body Substance|General Exam|8149,8154|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Procedure|Laboratory Procedure|General Exam|8149,8162|false|false|false|C0200949|Blood culture|Blood Culture
Drug|Biomedical or Dental Material|General Exam|8155,8162|false|false|false|C1706355|Culture Dose Form|Culture
Event|Event|General Exam|8155,8162|false|false|false|||Culture
Finding|Functional Concept|General Exam|8155,8162|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|Culture
Finding|Idea or Concept|General Exam|8155,8162|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|Culture
Procedure|Laboratory Procedure|General Exam|8155,8162|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|Culture
Finding|Idea or Concept|General Exam|8164,8171|false|false|false|C1691786;C1704475|Pending - Allergy Clinical Status;Pending - referral status|PENDING
Finding|Body Substance|General Exam|8206,8215|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|8206,8215|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|8206,8215|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|8206,8215|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|General Exam|8216,8220|false|false|false|||LABS
Lab|Laboratory or Test Result|General Exam|8216,8220|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|General Exam|8264,8269|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|8264,8269|false|false|false|||BLOOD
Finding|Body Substance|General Exam|8264,8269|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|8270,8273|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|8278,8281|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|8278,8281|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|8278,8281|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|8288,8291|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|8288,8291|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|8288,8291|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|8288,8291|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|8297,8300|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|8297,8300|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|8308,8311|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|8308,8311|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|8308,8311|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|8308,8311|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|8308,8311|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|8315,8318|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|8315,8318|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|8315,8318|false|false|false|||MCH
Finding|Gene or Genome|General Exam|8315,8318|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|8315,8318|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|8315,8318|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|8324,8328|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|8324,8328|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|8355,8358|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|8375,8380|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|8375,8380|false|false|false|||BLOOD
Finding|Body Substance|General Exam|8375,8380|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|8375,8388|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|8375,8388|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|8375,8388|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|8381,8388|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|8381,8388|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|8381,8388|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|8381,8388|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|8381,8388|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|8381,8388|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|8436,8440|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|8436,8440|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|8436,8440|false|false|false|C0202059|Bicarbonate measurement|HCO3
Event|Event|General Exam|8460,8463|false|false|false|||PMH
Finding|Finding|General Exam|8460,8463|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|PMH
Disorder|Disease or Syndrome|General Exam|8464,8467|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|General Exam|8464,8467|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|General Exam|8464,8467|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|General Exam|8464,8467|false|false|false|||CAD
Finding|Gene or Genome|General Exam|8464,8467|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|General Exam|8464,8467|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|General Exam|8464,8467|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|General Exam|8464,8467|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Finding|Functional Concept|General Exam|8472,8480|false|false|false|C0475224|Ischemic|ischemic
Event|Event|General Exam|8481,8483|false|false|false|||MR
Disorder|Disease or Syndrome|General Exam|8488,8491|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|General Exam|8488,8491|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|General Exam|8488,8491|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|General Exam|8488,8491|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|General Exam|8488,8491|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|General Exam|8488,8491|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Event|Event|General Exam|8488,8491|false|false|false|||DES
Finding|Gene or Genome|General Exam|8488,8491|false|false|false|C1413980|DES gene|DES
Procedure|Diagnostic Procedure|General Exam|8504,8507|false|false|false|C0430462|Transthoracic echocardiography|TTE
Finding|Intellectual Product|General Exam|8518,8522|false|false|false|C1547225|Mild Severity of Illness Code|mild
Disorder|Disease or Syndrome|General Exam|8532,8555|false|false|false|C1277187|Left ventricular systolic dysfunction|LV systolic dysfunction
Finding|Organ or Tissue Function|General Exam|8535,8543|false|false|false|C0039155|Systole|systolic
Finding|Pathologic Function|General Exam|8535,8555|false|false|false|C0749225|Systolic dysfunction|systolic dysfunction
Disorder|Disease or Syndrome|General Exam|8544,8555|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Event|Event|General Exam|8544,8555|false|false|false|||dysfunction
Finding|Conceptual Entity|General Exam|8544,8555|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|General Exam|8544,8555|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|General Exam|8544,8555|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Attribute|Clinical Attribute|General Exam|8565,8569|false|false|false|C0428772|Left ventricular ejection fraction|LVEF
Event|Event|General Exam|8565,8569|false|false|false|||LVEF
Procedure|Diagnostic Procedure|General Exam|8565,8569|false|false|false|C3837267|LVEF (procedure)|LVEF
Anatomy|Anatomical Structure|General Exam|8580,8583|false|false|false|C3669270|Strucure of thick cushion of skin|PAD
Disorder|Disease or Syndrome|General Exam|8580,8583|false|false|false|C0332568;C1704436|Pad Mass;Peripheral Arterial Diseases|PAD
Disorder|Neoplastic Process|General Exam|8580,8583|false|false|false|C0332568;C1704436|Pad Mass;Peripheral Arterial Diseases|PAD
Drug|Biomedical or Dental Material|General Exam|8580,8583|false|false|false|C2347441|Pad Dosage Form|PAD
Event|Event|General Exam|8580,8583|false|false|false|||PAD
Finding|Gene or Genome|General Exam|8580,8583|false|false|false|C1425244;C1425478;C3540603|DHX40 gene;PADI4 gene;PADI4 wt Allele|PAD
Procedure|Therapeutic or Preventive Procedure|General Exam|8580,8583|false|false|false|C3814046|PAD Regimen|PAD
Disorder|Disease or Syndrome|General Exam|8585,8588|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Event|Event|General Exam|8585,8588|false|false|false|||CKD
Attribute|Clinical Attribute|General Exam|8590,8595|false|false|false|C1300072|Tumor stage|stage
Anatomy|Body Location or Region|General Exam|8607,8610|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|General Exam|8607,8610|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|General Exam|8607,8610|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Finding|Finding|General Exam|8615,8621|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|General Exam|8615,8621|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Event|Event|General Exam|8622,8626|false|false|false|||UGIV
Event|Event|General Exam|8640,8648|false|false|false|||presents
Event|Event|General Exam|8663,8666|false|false|false|||SOB
Finding|Sign or Symptom|General Exam|8663,8666|false|false|false|C0013404|Dyspnea|SOB
Attribute|Clinical Attribute|General Exam|8668,8674|false|false|false|C0944911||weight
Event|Event|General Exam|8668,8674|false|false|false|||weight
Finding|Finding|General Exam|8668,8674|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|General Exam|8668,8674|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|General Exam|8668,8674|false|false|false|C1305866|Weighing patient|weight
Finding|Finding|General Exam|8668,8679|false|false|false|C0043094;C3814804|Gaining Weight question;Weight Gain|weight gain
Finding|Intellectual Product|General Exam|8668,8679|false|false|false|C0043094;C3814804|Gaining Weight question;Weight Gain|weight gain
Event|Event|General Exam|8675,8679|false|false|false|||gain
Finding|Intellectual Product|General Exam|8685,8690|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Part, Organ, or Organ Component|General Exam|8691,8696|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|General Exam|8691,8696|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Event|Event|General Exam|8691,8696|false|false|false|||heart
Finding|Sign or Symptom|General Exam|8691,8696|false|false|false|C0795691|HEART PROBLEM|heart
Finding|Functional Concept|General Exam|8698,8705|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|General Exam|8698,8705|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|General Exam|8698,8705|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|General Exam|8706,8718|false|false|false|||exacerbation
Finding|Finding|General Exam|8706,8718|false|false|false|C4086268|Exacerbation|exacerbation
Event|Event|General Exam|8735,8743|false|false|false|||diuresis
Finding|Organ or Tissue Function|General Exam|8735,8743|false|false|false|C0012797|Diuresis|diuresis
Drug|Organic Chemical|General Exam|8752,8757|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|General Exam|8752,8757|false|false|false|C0699992|Lasix|Lasix
Event|Event|General Exam|8752,8757|false|false|false|||Lasix
Event|Event|General Exam|8789,8800|false|false|false|||improvement
Finding|Conceptual Entity|General Exam|8789,8800|false|false|false|C2986411|Improvement|improvement
Attribute|Clinical Attribute|General Exam|8804,8814|false|false|false|C2979880||subjective
Finding|Finding|General Exam|8804,8814|false|false|false|C2266644|subjective (symptom)|subjective
Event|Event|General Exam|8815,8822|false|false|false|||dyspnea
Finding|Finding|General Exam|8815,8822|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|General Exam|8815,8822|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Event|Event|General Exam|8830,8836|true|false|false|||showed
Finding|Intellectual Product|General Exam|8840,8845|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Disease or Syndrome|General Exam|8840,8849|true|false|false|C3536663|Acute deep venous thrombosis|acute DVT
Anatomy|Body Location or Region|General Exam|8846,8849|true|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|General Exam|8846,8849|true|false|false|C2926618||DVT
Disorder|Disease or Syndrome|General Exam|8846,8849|true|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|General Exam|8846,8849|true|false|false|||DVT
Event|Event|General Exam|8851,8854|true|false|false|||CXR
Procedure|Diagnostic Procedure|General Exam|8851,8854|true|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|General Exam|8863,8867|true|false|false|||sign
Finding|Finding|General Exam|8863,8867|true|false|false|C0311392;C1547188|Language Ability - Sign;Physical findings|sign
Finding|Idea or Concept|General Exam|8863,8867|true|false|false|C0311392;C1547188|Language Ability - Sign;Physical findings|sign
Disorder|Disease or Syndrome|General Exam|8871,8884|true|false|false|C0521530|Lung consolidation|consolidation
Event|Event|General Exam|8871,8884|true|false|false|||consolidation
Event|Event|General Exam|8898,8909|true|false|false|||improvement
Finding|Conceptual Entity|General Exam|8898,8909|true|false|false|C2986411|Improvement|improvement
Event|Event|General Exam|8913,8920|true|false|false|||dyspnea
Finding|Finding|General Exam|8913,8920|true|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|General Exam|8913,8920|true|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Functional Concept|General Exam|8925,8937|true|false|false|C2348609|Supplement|supplemental
Event|Event|General Exam|8942,8953|true|false|false|||requirement
Finding|Functional Concept|General Exam|8942,8953|true|false|false|C1514873|Requirement|requirement
Finding|Body Substance|General Exam|8959,8966|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|General Exam|8959,8966|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|General Exam|8959,8966|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|General Exam|8971,8981|false|false|false|||discharged
Event|Event|General Exam|8983,8984|false|false|false|||/
Drug|Pharmacologic Substance|General Exam|8986,8996|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|General Exam|8986,8996|false|false|false|||medication
Finding|Intellectual Product|General Exam|8986,8996|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|General Exam|8997,9004|false|false|false|||changes
Finding|Functional Concept|General Exam|8997,9004|false|false|false|C0392747|Changing|changes
Attribute|Clinical Attribute|General Exam|9009,9028|false|false|false|C2707305||Shortness of breath
Finding|Sign or Symptom|General Exam|9009,9028|false|false|false|C0013404|Dyspnea|Shortness of breath
Finding|Body Substance|General Exam|9022,9028|false|false|false|C0225386|Breath|breath
Finding|Finding|General Exam|9031,9038|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|Hypoxia
Finding|Pathologic Function|General Exam|9031,9038|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|Hypoxia
Finding|Intellectual Product|General Exam|9041,9046|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Finding|General Exam|9041,9059|false|false|false|C0743630|exacerbation acute|acute exacerbation
Event|Event|General Exam|9047,9059|false|false|false|||exacerbation
Finding|Finding|General Exam|9047,9059|false|false|false|C4086268|Exacerbation|exacerbation
Finding|Intellectual Product|General Exam|9063,9070|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|General Exam|9063,9070|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|General Exam|9063,9094|false|false|false|C2711480|Chronic diastolic heart failure|chronic diastolic heart failure
Attribute|Clinical Attribute|General Exam|9071,9080|false|false|false|C0012000|Diastole|diastolic
Disorder|Disease or Syndrome|General Exam|9071,9094|false|false|false|C1135196|Heart Failure, Diastolic|diastolic heart failure
Anatomy|Body Part, Organ, or Organ Component|General Exam|9081,9086|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|General Exam|9081,9086|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|General Exam|9081,9086|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|General Exam|9081,9094|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Event|Event|General Exam|9087,9094|false|false|false|||failure
Finding|Functional Concept|General Exam|9087,9094|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|General Exam|9087,9094|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|General Exam|9087,9094|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|General Exam|9101,9110|false|false|false|||preserved
Attribute|Clinical Attribute|General Exam|9111,9115|false|false|false|C0428772|Left ventricular ejection fraction|LVEF
Event|Event|General Exam|9111,9115|false|false|false|||LVEF
Procedure|Diagnostic Procedure|General Exam|9111,9115|false|false|false|C3837267|LVEF (procedure)|LVEF
Attribute|Clinical Attribute|General Exam|9126,9132|false|false|false|C0944911||weight
Event|Event|General Exam|9126,9132|false|false|false|||weight
Finding|Finding|General Exam|9126,9132|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|General Exam|9126,9132|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|General Exam|9126,9132|false|false|false|C1305866|Weighing patient|weight
Procedure|Laboratory Procedure|General Exam|9144,9147|false|false|false|C3161851|liquid-based cytology (procedure)|lbs
Procedure|Health Care Activity|General Exam|9150,9159|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|General Exam|9160,9166|false|false|false|C0944911||weight
Event|Event|General Exam|9160,9166|false|false|false|||weight
Finding|Finding|General Exam|9160,9166|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|General Exam|9160,9166|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|General Exam|9160,9166|false|false|false|C1305866|Weighing patient|weight
Drug|Biomedical or Dental Material|General Exam|9173,9181|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|General Exam|9173,9181|false|false|false|||baseline
Finding|Idea or Concept|General Exam|9173,9181|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Drug|Amino Acid, Peptide, or Protein|General Exam|9183,9186|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Hormone|General Exam|9183,9186|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Pharmacologic Substance|General Exam|9183,9186|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Event|Event|General Exam|9183,9186|false|false|false|||BNP
Finding|Gene or Genome|General Exam|9183,9186|false|false|false|C1417808;C2982014|NPPB gene;NPPB wt Allele|BNP
Procedure|Laboratory Procedure|General Exam|9183,9186|false|false|false|C1095989|Brain natriuretic peptide measurement|BNP
Event|Event|General Exam|9188,9196|false|false|false|||elevated
Attribute|Clinical Attribute|General Exam|9209,9216|false|false|false|C0032930|Precipitating Factors|trigger
Finding|Idea or Concept|General Exam|9218,9225|false|false|false|C0750491;C1571873|Allergy Clinical Status - Suspect;Suspected (qualifier value)|suspect
Drug|Food|General Exam|9226,9233|false|true|false|C0012155|Diet|dietary
Event|Event|General Exam|9226,9233|false|false|false|||dietary
Event|Event|General Exam|9237,9249|false|false|false|||uncontrolled
Event|Event|General Exam|9258,9261|true|false|false|||EKG
Finding|Intellectual Product|General Exam|9258,9261|true|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|General Exam|9258,9261|true|false|false|C1623258|Electrocardiography|EKG
Event|Event|General Exam|9262,9269|true|false|false|||changes
Finding|Functional Concept|General Exam|9262,9269|true|false|false|C0392747|Changing|changes
Anatomy|Body Space or Junction|General Exam|9274,9277|true|false|false|C0262187|anterior calcarine sulcus (human only)|ACS
Disorder|Disease or Syndrome|General Exam|9274,9277|true|false|false|C0742343;C0796147|Acrocallosal Syndrome;Acute Chest Syndrome|ACS
Drug|Amino Acid, Peptide, or Protein|General Exam|9274,9277|true|false|false|C4042561|ACSS2 protein, human|ACS
Drug|Enzyme|General Exam|9274,9277|true|false|false|C4042561|ACSS2 protein, human|ACS
Event|Event|General Exam|9274,9277|true|false|false|||ACS
Finding|Gene or Genome|General Exam|9274,9277|true|false|false|C1150760;C1424787;C1825842;C1842089;C2266615;C4318612;C5400867;C5551036|ACCS gene;ACS - Activity Card Sort;ACSS2 gene;ACSS2 wt Allele;American Community Survey;CO-methylating acetyl-CoA synthase activity;PLA2G15 gene;acetate-CoA ligase activity|ACS
Finding|Intellectual Product|General Exam|9274,9277|true|false|false|C1150760;C1424787;C1825842;C1842089;C2266615;C4318612;C5400867;C5551036|ACCS gene;ACS - Activity Card Sort;ACSS2 gene;ACSS2 wt Allele;American Community Survey;CO-methylating acetyl-CoA synthase activity;PLA2G15 gene;acetate-CoA ligase activity|ACS
Finding|Molecular Function|General Exam|9274,9277|true|false|false|C1150760;C1424787;C1825842;C1842089;C2266615;C4318612;C5400867;C5551036|ACCS gene;ACS - Activity Card Sort;ACSS2 gene;ACSS2 wt Allele;American Community Survey;CO-methylating acetyl-CoA synthase activity;PLA2G15 gene;acetate-CoA ligase activity|ACS
Event|Event|General Exam|9284,9292|true|false|false|||negative
Finding|Classification|General Exam|9284,9292|true|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|General Exam|9284,9292|true|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|General Exam|9284,9292|true|false|false|C5237010|Expression Negative|negative
Finding|Functional Concept|General Exam|9294,9300|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Event|Event|General Exam|9301,9304|false|false|false|||TTE
Procedure|Diagnostic Procedure|General Exam|9301,9304|true|false|false|C0430462|Transthoracic echocardiography|TTE
Event|Event|General Exam|9305,9311|false|false|false|||showed
Finding|Intellectual Product|General Exam|9313,9317|false|false|false|C1547225|Mild Severity of Illness Code|mild
Disorder|Disease or Syndrome|General Exam|9327,9350|false|false|false|C1277187|Left ventricular systolic dysfunction|LV systolic dysfunction
Finding|Organ or Tissue Function|General Exam|9330,9338|false|false|false|C0039155|Systole|systolic
Finding|Pathologic Function|General Exam|9330,9350|false|false|false|C0749225|Systolic dysfunction|systolic dysfunction
Disorder|Disease or Syndrome|General Exam|9339,9350|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Event|Event|General Exam|9339,9350|false|false|false|||dysfunction
Finding|Conceptual Entity|General Exam|9339,9350|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|General Exam|9339,9350|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|General Exam|9339,9350|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Anatomy|Tissue|General Exam|9361,9371|false|false|false|C0027061|Myocardium|myocardial
Event|Event|General Exam|9373,9383|false|false|false|||infarction
Finding|Pathologic Function|General Exam|9373,9383|false|false|false|C0021308|Infarction|infarction
Event|Event|General Exam|9395,9404|false|false|false|||territory
Finding|Finding|General Exam|9409,9413|false|false|false|C5575035|Well (answer to question)|well
Finding|Classification|General Exam|9417,9422|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|Grade
Finding|Finding|General Exam|9417,9422|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|Grade
Finding|Classification|General Exam|9417,9425|false|false|false|C0441802;C0475270;C1522446;C4049999|Clavien-Dindo Grade II;Disease Grade 2;G2 stage (tumor staging);Grade two rank|Grade II
Finding|Intellectual Product|General Exam|9417,9425|false|false|false|C0441802;C0475270;C1522446;C4049999|Clavien-Dindo Grade II;Disease Grade 2;G2 stage (tumor staging);Grade two rank|Grade II
Attribute|Clinical Attribute|General Exam|9430,9439|false|false|false|C0012000|Diastole|diastolic
Finding|Pathologic Function|General Exam|9430,9451|false|false|false|C0520863|Diastolic dysfunction|diastolic dysfunction
Disorder|Disease or Syndrome|General Exam|9440,9451|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Event|Event|General Exam|9440,9451|false|false|false|||dysfunction
Finding|Conceptual Entity|General Exam|9440,9451|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|General Exam|9440,9451|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|General Exam|9440,9451|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Event|Event|General Exam|9456,9463|false|false|false|||similar
Event|Event|General Exam|9477,9480|false|false|false|||TTE
Procedure|Diagnostic Procedure|General Exam|9477,9480|false|false|false|C0430462|Transthoracic echocardiography|TTE
Finding|Mental Process|General Exam|9482,9487|false|false|false|C0870444|doubt|Doubt
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|9488,9491|false|false|false|C0600500|Peptide Nucleic Acids|PNA
Event|Event|General Exam|9488,9491|false|false|false|||PNA
Event|Event|General Exam|9499,9502|false|false|false|||CXR
Procedure|Diagnostic Procedure|General Exam|9499,9502|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|General Exam|9507,9511|false|false|false|||lack
Drug|Organic Chemical|General Exam|9515,9520|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|General Exam|9515,9520|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|General Exam|9515,9520|false|false|false|||cough
Finding|Sign or Symptom|General Exam|9515,9520|false|false|false|C0010200|Coughing|cough
Event|Event|General Exam|9521,9526|false|false|false|||fever
Finding|Finding|General Exam|9521,9526|false|false|true|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|General Exam|9521,9526|false|false|true|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|General Exam|9528,9533|false|false|false|||doubt
Finding|Mental Process|General Exam|9528,9533|false|false|false|C0870444|doubt|doubt
Finding|Finding|General Exam|9543,9546|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|General Exam|9543,9546|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Disorder|Disease or Syndrome|General Exam|9547,9552|false|false|false|C0343101|Wells syndrome|Wells
Event|Event|General Exam|9555,9560|false|false|false|||score
Finding|Finding|General Exam|9555,9560|false|false|false|C0449820|Score|score
Event|Event|General Exam|9570,9576|false|false|false|||stable
Finding|Intellectual Product|General Exam|9570,9576|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Functional Concept|General Exam|9577,9583|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Event|Event|General Exam|9599,9607|false|false|false|||diuresis
Finding|Organ or Tissue Function|General Exam|9599,9607|false|false|false|C0012797|Diuresis|diuresis
Drug|Organic Chemical|General Exam|9617,9622|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|General Exam|9617,9622|false|false|false|C0699992|Lasix|Lasix
Event|Event|General Exam|9653,9664|false|false|false|||improvement
Finding|Conceptual Entity|General Exam|9653,9664|false|false|false|C2986411|Improvement|improvement
Attribute|Clinical Attribute|General Exam|9668,9678|false|false|false|C2979880||subjective
Finding|Finding|General Exam|9668,9678|false|false|false|C2266644|subjective (symptom)|subjective
Event|Event|General Exam|9680,9687|false|false|false|||dyspnea
Finding|Finding|General Exam|9680,9687|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|General Exam|9680,9687|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Event|Event|General Exam|9698,9702|false|false|false|||home
Finding|Idea or Concept|General Exam|9698,9702|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|General Exam|9698,9702|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|General Exam|9698,9702|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|General Exam|9703,9712|false|false|false|C0076840|torsemide|torsemide
Drug|Pharmacologic Substance|General Exam|9703,9712|false|false|false|C0076840|torsemide|torsemide
Drug|Organic Chemical|General Exam|9719,9729|false|false|false|C0028066|nifedipine|nifedipine
Drug|Pharmacologic Substance|General Exam|9719,9729|false|false|false|C0028066|nifedipine|nifedipine
Disorder|Mental or Behavioral Dysfunction|General Exam|9735,9738|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|General Exam|9735,9738|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|General Exam|9735,9738|false|false|false|C1530795|BID protein, human|BID
Event|Event|General Exam|9735,9738|false|false|false|||BID
Finding|Gene or Genome|General Exam|9735,9738|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|General Exam|9744,9754|false|false|false|C0054836|carvedilol|carvedilol
Drug|Pharmacologic Substance|General Exam|9744,9754|false|false|false|C0054836|carvedilol|carvedilol
Disorder|Mental or Behavioral Dysfunction|General Exam|9760,9763|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|General Exam|9760,9763|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|General Exam|9760,9763|false|false|false|C1530795|BID protein, human|BID
Event|Event|General Exam|9760,9763|false|false|false|||BID
Finding|Gene or Genome|General Exam|9760,9763|false|false|false|C1332410|BID gene|BID
Event|Event|General Exam|9770,9776|false|false|false|||stable
Finding|Intellectual Product|General Exam|9770,9776|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|General Exam|9792,9801|false|false|false|||discharge
Finding|Body Substance|General Exam|9792,9801|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|General Exam|9792,9801|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|General Exam|9792,9801|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|General Exam|9792,9801|false|false|false|C0030685|Patient Discharge|discharge
Disorder|Disease or Syndrome|General Exam|9806,9818|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|General Exam|9806,9818|false|false|false|||Hypertension
Finding|Body Substance|General Exam|9821,9828|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|General Exam|9821,9828|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|General Exam|9821,9828|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|General Exam|9829,9835|false|false|false|||missed
Attribute|Clinical Attribute|General Exam|9848,9859|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|General Exam|9848,9859|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|General Exam|9848,9859|false|false|false|||medications
Finding|Intellectual Product|General Exam|9848,9859|false|false|false|C4284232|Medications|medications
Finding|Idea or Concept|General Exam|9869,9872|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|General Exam|9869,9872|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|General Exam|9876,9885|false|false|false|||admission
Procedure|Health Care Activity|General Exam|9876,9885|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|General Exam|9887,9896|false|false|false|||Continued
Finding|Idea or Concept|General Exam|9897,9901|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|General Exam|9897,9901|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|General Exam|9897,9901|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|General Exam|9902,9912|false|false|false|C0054836|carvedilol|carvedilol
Drug|Pharmacologic Substance|General Exam|9902,9912|false|false|false|C0054836|carvedilol|carvedilol
Disorder|Mental or Behavioral Dysfunction|General Exam|9918,9921|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|General Exam|9918,9921|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|General Exam|9918,9921|false|false|false|C1530795|BID protein, human|BID
Event|Event|General Exam|9918,9921|false|false|false|||BID
Finding|Gene or Genome|General Exam|9918,9921|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|General Exam|9927,9937|false|false|false|C0028066|nifedipine|nifedipine
Drug|Pharmacologic Substance|General Exam|9927,9937|false|false|false|C0028066|nifedipine|nifedipine
Disorder|Mental or Behavioral Dysfunction|General Exam|9943,9946|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|General Exam|9943,9946|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|General Exam|9943,9946|false|false|false|C1530795|BID protein, human|BID
Event|Event|General Exam|9943,9946|false|false|false|||BID
Finding|Gene or Genome|General Exam|9943,9946|false|false|false|C1332410|BID gene|BID
Event|Event|General Exam|9960,9970|false|false|false|||parameters
Finding|Finding|General Exam|9960,9970|false|false|false|C0449381|Observation parameter|parameters
Event|Event|General Exam|9972,9979|false|false|false|||Appears
Event|Event|General Exam|9988,9993|false|false|false|||trial
Procedure|Research Activity|General Exam|9988,9993|false|false|false|C0008976|Clinical Trials|trial
Drug|Organic Chemical|General Exam|10004,10018|false|false|false|C0037982|spironolactone|spironolactone
Drug|Pharmacologic Substance|General Exam|10004,10018|false|false|false|C0037982|spironolactone|spironolactone
Event|Event|General Exam|10004,10018|false|false|false|||spironolactone
Event|Event|General Exam|10028,10035|false|false|false|||limited
Event|Event|General Exam|10040,10052|false|false|false|||hyperkalemia
Finding|Finding|General Exam|10040,10052|false|false|false|C0020461;C5700154|Hyperkalemia;Serum potassium level above reference range|hyperkalemia
Event|Event|General Exam|10066,10074|false|false|false|||deferred
Anatomy|Body Part, Organ, or Organ Component|General Exam|10084,10091|false|false|false|C0042027|Urinary tract|Urinary
Finding|Finding|General Exam|10084,10101|false|false|false|C0042023|Increased frequency of micturition|Urinary frequency
Event|Event|General Exam|10092,10101|false|false|false|||frequency
Finding|Intellectual Product|General Exam|10092,10101|false|false|false|C3898838;C4321352|Frequency;How Often|frequency
Finding|Finding|General Exam|10102,10119|false|false|false|C0150045|Urge Incontinence|urge incontinence
Disorder|Disease or Syndrome|General Exam|10107,10119|false|false|false|C0021167|Incontinence|incontinence
Event|Event|General Exam|10107,10119|false|false|false|||incontinence
Event|Event|General Exam|10121,10129|false|false|false|||occurred
Finding|Mental Process|General Exam|10133,10140|false|false|false|C0542559|contextual factors|setting
Event|Event|General Exam|10145,10153|false|false|false|||diuresis
Finding|Organ or Tissue Function|General Exam|10145,10153|false|false|false|C0012797|Diuresis|diuresis
Event|Event|General Exam|10167,10174|false|false|false|||ordered
Event|Event|General Exam|10190,10201|false|false|false|||enterococci
Finding|Finding|General Exam|10203,10209|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|General Exam|10203,10209|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|General Exam|10211,10223|false|false|false|||colonization
Finding|Finding|General Exam|10211,10223|false|false|false|C4289767|Colonization|colonization
Event|Event|General Exam|10228,10236|false|false|false|||symptoms
Finding|Functional Concept|General Exam|10228,10236|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|General Exam|10228,10236|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|General Exam|10237,10245|false|false|false|||persists
Event|Event|General Exam|10279,10286|false|false|false|||CHRONIC
Finding|Intellectual Product|General Exam|10279,10286|false|false|false|C1547296|Chronic - Admission Level of Care Code|CHRONIC
Procedure|Health Care Activity|General Exam|10279,10286|false|false|false|C1555457|Provision of recurring care for chronic illness|CHRONIC
Finding|Intellectual Product|General Exam|10287,10293|false|false|false|C1547311|Patient Condition Code - Stable|STABLE
Event|Event|General Exam|10294,10300|false|false|false|||ISSUES
Disorder|Disease or Syndrome|General Exam|10315,10321|false|false|false|C0002871|Anemia|anemia
Event|Event|General Exam|10315,10321|false|false|false|||anemia
Drug|Biomedical or Dental Material|General Exam|10330,10338|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|General Exam|10330,10338|false|false|false|||baseline
Finding|Idea or Concept|General Exam|10330,10338|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Drug|Biomedical or Dental Material|General Exam|10363,10371|true|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|General Exam|10363,10371|true|false|false|||baseline
Finding|Idea or Concept|General Exam|10363,10371|true|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|General Exam|10376,10381|true|false|false|||signs
Finding|Finding|General Exam|10376,10381|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|General Exam|10376,10381|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Event|Event|General Exam|10392,10400|true|false|false|||bleeding
Finding|Pathologic Function|General Exam|10392,10400|true|false|false|C0019080|Hemorrhage|bleeding
Finding|Finding|General Exam|10403,10409|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Idea or Concept|General Exam|10403,10409|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Event|Event|General Exam|10410,10424|false|false|false|||multifactorial
Finding|Finding|General Exam|10410,10424|false|true|false|C1837655|Multifactorial|multifactorial
Disorder|Disease or Syndrome|General Exam|10427,10433|false|false|false|C0002871|Anemia|anemia
Event|Event|General Exam|10427,10433|false|false|false|||anemia
Disorder|Disease or Syndrome|General Exam|10427,10452|false|false|false|C0002873|Anemia of chronic disease|anemia of chronic disease
Finding|Intellectual Product|General Exam|10437,10444|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|General Exam|10437,10444|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|General Exam|10437,10452|false|false|false|C0008679|Chronic disease|chronic disease
Disorder|Disease or Syndrome|General Exam|10445,10452|false|false|false|C0012634|Disease|disease
Event|Event|General Exam|10445,10452|false|false|false|||disease
Finding|Finding|General Exam|10456,10460|false|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|10474,10487|false|false|false|||erythropoiten
Event|Event|General Exam|10489,10499|false|false|false|||production
Event|Occupational Activity|General Exam|10489,10499|false|false|false|C0033268|production|production
Finding|Intellectual Product|General Exam|10489,10499|false|false|false|C1548180|Production Processing ID|production
Disorder|Disease or Syndrome|General Exam|10504,10507|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Event|Event|General Exam|10504,10507|false|false|false|||CKD
Drug|Element, Ion, or Isotope|General Exam|10517,10522|false|false|false|C0003075|Anions|anion
Attribute|Clinical Attribute|General Exam|10517,10526|false|false|false|C0003074|Anion Gap|anion gap
Lab|Laboratory or Test Result|General Exam|10517,10526|false|false|false|C1509129|Anion gap result|anion gap
Procedure|Laboratory Procedure|General Exam|10517,10526|false|false|false|C0201889;C2189246|Anion gap measurement;blood anion gap (lab test)|anion gap
Drug|Amino Acid, Peptide, or Protein|General Exam|10523,10526|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|gap
Drug|Biologically Active Substance|General Exam|10523,10526|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|gap
Event|Event|General Exam|10523,10526|false|false|false|||gap
Finding|Gene or Genome|General Exam|10523,10526|false|false|false|C1419277;C2984552|RASA1 gene;RASA1 wt Allele|gap
Event|Event|General Exam|10527,10536|false|false|false|||metabolic
Finding|Cell Function|General Exam|10527,10536|false|false|false|C0311400;C1524026|Metabolic;Metabolic Process, Cellular|metabolic
Finding|Functional Concept|General Exam|10527,10536|false|false|false|C0311400;C1524026|Metabolic;Metabolic Process, Cellular|metabolic
Procedure|Diagnostic Procedure|General Exam|10527,10536|false|false|false|C4263342|Multisection metabolic|metabolic
Finding|Pathologic Function|General Exam|10527,10545|false|false|false|C0220981|Metabolic acidosis|metabolic acidosis
Event|Event|General Exam|10537,10545|false|false|false|||acidosis
Finding|Pathologic Function|General Exam|10537,10545|false|false|false|C0001122|Acidosis|acidosis
Finding|Body Substance|General Exam|10548,10555|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|General Exam|10548,10555|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|General Exam|10548,10555|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Functional Concept|General Exam|10548,10559|false|false|false|C0332310|Has patient|Patient has
Event|Event|General Exam|10582,10587|false|false|false|||NAGMA
Event|Event|General Exam|10612,10620|true|false|false|||diarrhea
Finding|Finding|General Exam|10612,10620|true|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|General Exam|10612,10620|true|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Event|Event|General Exam|10627,10634|false|false|false|||suspect
Finding|Gene or Genome|General Exam|10635,10639|false|true|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|Type
Finding|Intellectual Product|General Exam|10635,10639|false|true|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|Type
Disorder|Disease or Syndrome|General Exam|10644,10647|false|false|false|C0001126|Renal tubular acidosis|RTA
Event|Event|General Exam|10644,10647|false|false|false|||RTA
Finding|Gene or Genome|General Exam|10644,10647|false|false|false|C1419304;C1428415;C3889271|HHV8 ORF50 Gene;MRGPRF gene;RBFOX2 gene|RTA
Event|Event|General Exam|10654,10662|false|false|false|||advanced
Attribute|Clinical Attribute|General Exam|10663,10666|false|false|false|C1114365||age
Drug|Biologically Active Substance|General Exam|10663,10666|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|General Exam|10663,10666|false|false|false|C0162574|Glycation End Products, Advanced|age
Event|Event|General Exam|10671,10678|false|false|false|||history
Finding|Conceptual Entity|General Exam|10671,10678|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|General Exam|10671,10678|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|General Exam|10671,10678|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|General Exam|10671,10681|false|false|false|C0262926|Medical History|history of
Event|Event|General Exam|10713,10726|false|false|false|||hyporeninemia
Attribute|Clinical Attribute|General Exam|10732,10737|false|false|false|C1300072|Tumor stage|Stage
Finding|Intellectual Product|General Exam|10732,10740|false|false|false|C0441772|Stage level 4|Stage IV
Finding|Intellectual Product|General Exam|10741,10748|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|General Exam|10741,10748|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Disorder|Disease or Syndrome|General Exam|10741,10763|false|false|false|C1561643|Chronic Kidney Diseases|Chronic Kidney Disease
Anatomy|Body Part, Organ, or Organ Component|General Exam|10749,10755|false|false|false|C0022646;C0227665|Both kidneys;Kidney|Kidney
Disorder|Neoplastic Process|General Exam|10749,10755|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|Kidney
Finding|Sign or Symptom|General Exam|10749,10755|false|false|false|C0812426|Kidney problem|Kidney
Procedure|Diagnostic Procedure|General Exam|10749,10755|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|Kidney
Procedure|Therapeutic or Preventive Procedure|General Exam|10749,10755|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|Kidney
Disorder|Disease or Syndrome|General Exam|10749,10763|false|false|false|C0022658|Kidney Diseases|Kidney Disease
Disorder|Disease or Syndrome|General Exam|10756,10763|false|false|false|C0012634|Disease|Disease
Event|Event|General Exam|10756,10763|false|false|false|||Disease
Drug|Biomedical or Dental Material|General Exam|10765,10773|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|General Exam|10765,10773|false|false|false|||baseline
Finding|Idea or Concept|General Exam|10765,10773|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Disorder|Disease or Syndrome|General Exam|10788,10791|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Event|Event|General Exam|10788,10791|false|false|false|||CKD
Disorder|Disease or Syndrome|General Exam|10797,10800|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|General Exam|10797,10800|false|false|false|||HTN
Drug|Biomedical or Dental Material|General Exam|10830,10838|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|General Exam|10830,10838|false|false|false|||baseline
Finding|Idea or Concept|General Exam|10830,10838|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Finding|General Exam|10840,10843|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|Low
Finding|Intellectual Product|General Exam|10840,10843|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|Low
Event|Event|General Exam|10844,10845|false|false|false|||K
Drug|Food|General Exam|10855,10859|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|General Exam|10855,10859|false|false|false|||diet
Finding|Functional Concept|General Exam|10855,10859|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|General Exam|10855,10859|false|false|false|C0012159|Diet therapy|diet
Event|Event|General Exam|10861,10870|false|false|false|||Continued
Finding|Idea or Concept|General Exam|10871,10875|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|General Exam|10871,10875|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|General Exam|10871,10875|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|General Exam|10876,10886|false|false|false|C0006674;C3714610|Calcitriol Drug Class;calcitriol|calcitriol
Drug|Pharmacologic Substance|General Exam|10876,10886|false|false|false|C0006674;C3714610|Calcitriol Drug Class;calcitriol|calcitriol
Drug|Vitamin|General Exam|10876,10886|false|false|false|C0006674;C3714610|Calcitriol Drug Class;calcitriol|calcitriol
Event|Event|General Exam|10876,10886|false|false|false|||calcitriol
Event|Event|General Exam|10922,10927|false|false|false|||dosed
Attribute|Clinical Attribute|General Exam|10932,10943|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|General Exam|10932,10943|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|General Exam|10932,10943|false|false|false|||medications
Finding|Intellectual Product|General Exam|10932,10943|false|false|false|C4284232|Medications|medications
Anatomy|Body Part, Organ, or Organ Component|General Exam|10948,10956|false|false|false|C0018787|Heart|Coronary
Anatomy|Body Part, Organ, or Organ Component|General Exam|10948,10963|false|false|false|C0205042|Coronary artery|Coronary artery
Disorder|Disease or Syndrome|General Exam|10948,10971|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|Coronary artery disease
Anatomy|Body Part, Organ, or Organ Component|General Exam|10957,10963|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|General Exam|10957,10963|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Disorder|Disease or Syndrome|General Exam|10957,10971|false|false|false|C0852949|Arteriopathic disease|artery disease
Disorder|Disease or Syndrome|General Exam|10964,10971|false|false|false|C0012634|Disease|disease
Event|Event|General Exam|10964,10971|false|false|false|||disease
Disorder|Disease or Syndrome|General Exam|10976,10979|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|General Exam|10976,10979|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|General Exam|10976,10979|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|General Exam|10976,10979|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|General Exam|10976,10979|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|General Exam|10976,10979|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Event|Event|General Exam|10976,10979|false|false|false|||DES
Finding|Gene or Genome|General Exam|10976,10979|false|false|false|C1413980|DES gene|DES
Drug|Amino Acid, Peptide, or Protein|General Exam|10983,10986|false|false|false|C2987138|Methylcytosine Dioxygenase TET1|LCX
Drug|Enzyme|General Exam|10983,10986|false|false|false|C2987138|Methylcytosine Dioxygenase TET1|LCX
Event|Event|General Exam|10983,10986|false|false|false|||LCX
Finding|Gene or Genome|General Exam|10983,10986|false|false|false|C1428863;C2987137|TET1 gene;TET1 wt Allele|LCX
Drug|Amino Acid, Peptide, or Protein|General Exam|10992,11001|false|false|false|C0041199|Troponin|troponins
Drug|Biologically Active Substance|General Exam|10992,11001|false|false|false|C0041199|Troponin|troponins
Event|Event|General Exam|10992,11001|false|false|false|||troponins
Event|Event|General Exam|11008,11015|false|false|false|||trended
Finding|Intellectual Product|General Exam|11044,11048|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|General Exam|11049,11056|false|false|false|||stopped
Drug|Amino Acid, Peptide, or Protein|General Exam|11058,11063|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|General Exam|11058,11063|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|General Exam|11058,11063|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|General Exam|11058,11063|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Event|Event|General Exam|11061,11063|false|false|false|||MB
Event|Event|General Exam|11069,11073|false|false|false|||flat
Finding|Body Substance|General Exam|11076,11083|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|General Exam|11076,11083|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|General Exam|11076,11083|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|General Exam|11084,11091|true|false|false|||deneied
Anatomy|Body Location or Region|General Exam|11096,11101|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|General Exam|11096,11101|true|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|General Exam|11096,11106|true|false|false|C2926613||chest pain
Finding|Sign or Symptom|General Exam|11096,11106|true|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|General Exam|11102,11106|true|false|false|C2598155||pain
Event|Event|General Exam|11102,11106|true|false|false|||pain
Finding|Functional Concept|General Exam|11102,11106|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|General Exam|11102,11106|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|General Exam|11110,11113|false|false|false|||TTE
Procedure|Diagnostic Procedure|General Exam|11110,11113|false|false|false|C0430462|Transthoracic echocardiography|TTE
Event|Event|General Exam|11114,11120|false|false|false|||showed
Finding|Intellectual Product|General Exam|11121,11125|false|false|false|C1547225|Mild Severity of Illness Code|mild
Disorder|Disease or Syndrome|General Exam|11136,11159|false|false|false|C1277187|Left ventricular systolic dysfunction|LV systolic dysfunction
Finding|Organ or Tissue Function|General Exam|11139,11147|false|false|false|C0039155|Systole|systolic
Finding|Pathologic Function|General Exam|11139,11159|false|false|false|C0749225|Systolic dysfunction|systolic dysfunction
Disorder|Disease or Syndrome|General Exam|11148,11159|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Event|Event|General Exam|11148,11159|false|false|false|||dysfunction
Finding|Conceptual Entity|General Exam|11148,11159|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|General Exam|11148,11159|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|General Exam|11148,11159|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Finding|General Exam|11164,11191|false|false|false|C0155668|Old myocardial infarction|prior myocardial infarction
Anatomy|Tissue|General Exam|11170,11180|false|false|false|C0027061|Myocardium|myocardial
Attribute|Clinical Attribute|General Exam|11170,11191|false|false|false|C2926063||myocardial infarction
Disorder|Disease or Syndrome|General Exam|11170,11191|false|false|false|C0027051|Myocardial Infarction|myocardial infarction
Event|Event|General Exam|11181,11191|false|false|false|||infarction
Finding|Pathologic Function|General Exam|11181,11191|false|false|false|C0021308|Infarction|infarction
Event|Event|General Exam|11204,11213|false|false|false|||territory
Event|Event|General Exam|11218,11225|false|false|false|||similar
Event|Event|General Exam|11239,11242|false|false|false|||TTE
Procedure|Diagnostic Procedure|General Exam|11239,11242|false|false|false|C0430462|Transthoracic echocardiography|TTE
Event|Event|General Exam|11244,11253|false|false|false|||Continued
Finding|Idea or Concept|General Exam|11255,11259|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|General Exam|11255,11259|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|General Exam|11255,11259|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|General Exam|11260,11267|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|General Exam|11260,11267|false|false|false|C0004057|aspirin|aspirin
Event|Event|General Exam|11260,11267|false|false|false|||aspirin
Finding|Idea or Concept|General Exam|11277,11281|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|General Exam|11277,11281|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|General Exam|11277,11281|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|General Exam|11282,11292|false|false|false|C0054836|carvedilol|carvedilol
Drug|Pharmacologic Substance|General Exam|11282,11292|false|false|false|C0054836|carvedilol|carvedilol
Disorder|Mental or Behavioral Dysfunction|General Exam|11298,11301|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|General Exam|11298,11301|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|General Exam|11298,11301|false|false|false|C1530795|BID protein, human|BID
Event|Event|General Exam|11298,11301|false|false|false|||BID
Finding|Gene or Genome|General Exam|11298,11301|false|false|false|C1332410|BID gene|BID
Event|Event|General Exam|11307,11314|false|false|false|||holding
Event|Event|General Exam|11316,11326|false|false|false|||parameters
Finding|Finding|General Exam|11316,11326|false|false|false|C0449381|Observation parameter|parameters
Finding|Idea or Concept|General Exam|11328,11332|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|General Exam|11328,11332|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|General Exam|11328,11332|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|General Exam|11333,11345|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|General Exam|11333,11345|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|General Exam|11333,11345|false|false|false|||atorvastatin
Event|Event|General Exam|11351,11354|false|false|false|||qHS
Finding|Gene or Genome|General Exam|11360,11364|false|true|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|Type
Finding|Intellectual Product|General Exam|11360,11364|false|true|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|Type
Disorder|Disease or Syndrome|General Exam|11360,11376|false|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|Type II Diabetes
Disorder|Disease or Syndrome|General Exam|11360,11385|false|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|Type II Diabetes Mellitus
Disorder|Disease or Syndrome|General Exam|11368,11376|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|Diabetes
Disorder|Disease or Syndrome|General Exam|11368,11385|false|false|false|C0011849|Diabetes Mellitus|Diabetes Mellitus
Event|Event|General Exam|11377,11385|false|false|false|||Mellitus
Drug|Amino Acid, Peptide, or Protein|General Exam|11392,11397|false|false|false|C0019018|Glycosylated hemoglobin A|HbA1C
Drug|Biologically Active Substance|General Exam|11392,11397|false|false|false|C0019018|Glycosylated hemoglobin A|HbA1C
Procedure|Laboratory Procedure|General Exam|11392,11397|false|false|false|C0202054|Glucohemoglobin measurement|HbA1C
Drug|Organic Chemical|General Exam|11426,11433|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|General Exam|11426,11433|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|General Exam|11426,11433|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Event|Event|General Exam|11426,11433|false|false|false|||control
Finding|Conceptual Entity|General Exam|11426,11433|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|General Exam|11426,11433|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|General Exam|11426,11433|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Disorder|Disease or Syndrome|General Exam|11456,11468|false|false|false|C0362046|Prediabetes syndrome|pre-diabetic
Event|Event|General Exam|11469,11474|false|false|false|||range
Finding|Intellectual Product|General Exam|11469,11474|false|false|false|C3542016|Concept model range (foundation metadata concept)|range
Event|Event|General Exam|11478,11486|false|false|false|||Continue
Finding|Idea or Concept|General Exam|11478,11486|false|false|false|C0549178|Continuous|Continue
Event|Event|General Exam|11487,11491|false|false|false|||home
Finding|Idea or Concept|General Exam|11487,11491|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|General Exam|11487,11491|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|General Exam|11487,11491|false|false|false|C1553498|home health encounter|home
Anatomy|Body Part, Organ, or Organ Component|General Exam|11506,11511|false|false|false|C0222045|Integumentary scale|scale
Event|Activity|General Exam|11506,11511|false|false|false|C1947916|Scaling|scale
Finding|Conceptual Entity|General Exam|11506,11511|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Finding|Intellectual Product|General Exam|11506,11511|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Finding|Daily or Recreational Activity|General Exam|11518,11524|false|false|false|C4048877|Dinner|dinner
Disorder|Disease or Syndrome|General Exam|11529,11534|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|General Exam|11529,11534|false|false|false|||blood
Finding|Body Substance|General Exam|11529,11534|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Organic Chemical|General Exam|11529,11540|false|false|false|C0005802|Blood Glucose|blood sugar
Procedure|Laboratory Procedure|General Exam|11529,11540|false|false|false|C0392201|Blood glucose measurement|blood sugar
Drug|Biomedical or Dental Material|General Exam|11535,11540|false|false|false|C0007004;C0242209;C3665462|Carbohydrates;Sugars;raw sugar|sugar
Drug|Organic Chemical|General Exam|11535,11540|false|false|false|C0007004;C0242209;C3665462|Carbohydrates;Sugars;raw sugar|sugar
Drug|Pharmacologic Substance|General Exam|11535,11540|false|false|false|C0007004;C0242209;C3665462|Carbohydrates;Sugars;raw sugar|sugar
Event|Event|General Exam|11535,11540|false|false|false|||sugar
Disorder|Disease or Syndrome|General Exam|11576,11581|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|General Exam|11576,11581|false|false|false|||blood
Finding|Body Substance|General Exam|11576,11581|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Organic Chemical|General Exam|11576,11587|false|false|false|C0005802|Blood Glucose|blood sugar
Procedure|Laboratory Procedure|General Exam|11576,11587|false|false|false|C0392201|Blood glucose measurement|blood sugar
Drug|Biomedical or Dental Material|General Exam|11582,11587|false|false|false|C0007004;C0242209;C3665462|Carbohydrates;Sugars;raw sugar|sugar
Drug|Organic Chemical|General Exam|11582,11587|false|false|false|C0007004;C0242209;C3665462|Carbohydrates;Sugars;raw sugar|sugar
Drug|Pharmacologic Substance|General Exam|11582,11587|false|false|false|C0007004;C0242209;C3665462|Carbohydrates;Sugars;raw sugar|sugar
Event|Event|General Exam|11582,11587|false|false|false|||sugar
Event|Event|General Exam|11588,11593|false|false|false|||under
Disorder|Disease or Syndrome|General Exam|11603,11615|false|false|false|C0242339|Dyslipidemias|Dyslipidemia
Event|Event|General Exam|11603,11615|false|false|false|||Dyslipidemia
Event|Event|General Exam|11617,11626|false|false|false|||continued
Finding|Idea or Concept|General Exam|11627,11631|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|General Exam|11627,11631|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|General Exam|11627,11631|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|General Exam|11632,11644|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|General Exam|11632,11644|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|General Exam|11632,11644|false|false|false|||atorvastatin
Drug|Pharmacologic Substance|General Exam|11648,11656|false|false|false|C1950154|Insomnia homeopathic medication|Insomnia
Event|Event|General Exam|11648,11656|false|false|false|||Insomnia
Finding|Sign or Symptom|General Exam|11648,11656|false|false|false|C0917801|Sleeplessness|Insomnia
Event|Event|General Exam|11658,11667|false|false|false|||continued
Finding|Idea or Concept|General Exam|11668,11672|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|General Exam|11668,11672|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|General Exam|11668,11672|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|General Exam|11673,11683|false|false|false|C0060926|gabapentin|gabapentin
Drug|Pharmacologic Substance|General Exam|11673,11683|false|false|false|C0060926|gabapentin|gabapentin
Event|Event|General Exam|11673,11683|false|false|false|||gabapentin
Disorder|Disease or Syndrome|General Exam|11687,11691|false|false|false|C0018099|Gout|Gout
Event|Event|General Exam|11687,11691|false|false|false|||Gout
Event|Event|General Exam|11693,11702|false|false|false|||continued
Finding|Idea or Concept|General Exam|11703,11707|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|General Exam|11703,11707|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|General Exam|11703,11707|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|General Exam|11708,11719|false|false|false|C0002144|allopurinol|allopurinol
Drug|Pharmacologic Substance|General Exam|11708,11719|false|false|false|C0002144|allopurinol|allopurinol
Event|Event|General Exam|11708,11719|false|false|false|||allopurinol
Finding|Idea or Concept|General Exam|11754,11766|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Event|Event|General Exam|11807,11816|false|false|false|||Discharge
Finding|Body Substance|General Exam|11807,11816|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|General Exam|11807,11816|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|General Exam|11807,11816|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|General Exam|11807,11816|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|General Exam|11817,11823|false|false|false|C0944911||weight
Event|Event|General Exam|11817,11823|false|false|false|||weight
Finding|Finding|General Exam|11817,11823|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|General Exam|11817,11823|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|General Exam|11817,11823|false|false|false|C1305866|Weighing patient|weight
Event|Event|General Exam|11834,11843|false|false|false|||Discharge
Finding|Body Substance|General Exam|11834,11843|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|General Exam|11834,11843|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|General Exam|11834,11843|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|General Exam|11834,11843|false|false|false|C0030685|Patient Discharge|Discharge
Drug|Biologically Active Substance|General Exam|11844,11854|false|false|false|C0010294|creatinine|creatinine
Drug|Organic Chemical|General Exam|11844,11854|false|false|false|C0010294|creatinine|creatinine
Event|Event|General Exam|11844,11854|false|false|false|||creatinine
Finding|Physiologic Function|General Exam|11844,11854|false|false|false|C4551889|Creatinine metabolic function|creatinine
Procedure|Laboratory Procedure|General Exam|11844,11854|false|false|false|C0201975|Creatinine measurement|creatinine
Event|Event|General Exam|11862,11871|false|false|false|||Discharge
Finding|Body Substance|General Exam|11862,11871|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|General Exam|11862,11871|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|General Exam|11862,11871|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|General Exam|11862,11871|false|false|false|C0030685|Patient Discharge|Discharge
Anatomy|Body Space or Junction|General Exam|11872,11876|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|General Exam|11872,11876|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|General Exam|11872,11876|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|General Exam|11872,11876|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Pharmacologic Substance|General Exam|11877,11885|false|false|false|C0012798;C5399719|Diuretic [APC];Diuretics|diuretic
Event|Event|General Exam|11877,11885|false|false|false|||diuretic
Drug|Organic Chemical|General Exam|11887,11896|false|false|false|C0076840|torsemide|torsemide
Drug|Pharmacologic Substance|General Exam|11887,11896|false|false|false|C0076840|torsemide|torsemide
Finding|Idea or Concept|General Exam|11910,11922|false|false|false|C1548597|Marketing basis - Transitional|Transitional
Event|Activity|General Exam|11923,11928|false|false|false|C5966184|Issue (action)|issue
Event|Event|General Exam|11923,11928|false|false|false|||issue
Finding|Finding|General Exam|11923,11928|false|false|false|C0033213;C1706387|Issue (document);Problem|issue
Finding|Intellectual Product|General Exam|11923,11928|false|false|false|C0033213;C1706387|Issue (document);Problem|issue
Event|Event|General Exam|11930,11938|false|false|false|||consider
Finding|Classification|General Exam|11939,11949|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|General Exam|11939,11949|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Drug|Amino Acid, Peptide, or Protein|General Exam|11950,11953|false|false|false|C0014822;C0357126;C2976467|EPO protein, human;Erythropoietin;epoetin alfa|epo
Drug|Biologically Active Substance|General Exam|11950,11953|false|false|false|C0014822;C0357126;C2976467|EPO protein, human;Erythropoietin;epoetin alfa|epo
Drug|Hormone|General Exam|11950,11953|false|false|false|C0014822;C0357126;C2976467|EPO protein, human;Erythropoietin;epoetin alfa|epo
Drug|Pharmacologic Substance|General Exam|11950,11953|false|false|false|C0014822;C0357126;C2976467|EPO protein, human;Erythropoietin;epoetin alfa|epo
Event|Event|General Exam|11950,11953|false|false|false|||epo
Finding|Gene or Genome|General Exam|11950,11953|false|false|false|C1366564;C1367459;C1414438;C1705819;C3496094|EPO gene;EPX gene;Exclusive Provider Organization Plan;TIMP1 gene;TIMP1 wt Allele|epo
Finding|Intellectual Product|General Exam|11950,11953|false|false|false|C1366564;C1367459;C1414438;C1705819;C3496094|EPO gene;EPX gene;Exclusive Provider Organization Plan;TIMP1 gene;TIMP1 wt Allele|epo
Anatomy|Body Part, Organ, or Organ Component|General Exam|11959,11964|false|false|false|C0022646|Kidney|renal
Disorder|Disease or Syndrome|General Exam|11959,11964|false|false|false|C0042075|Urologic Diseases|renal
Finding|Idea or Concept|General Exam|11968,11980|false|false|false|C1548597|Marketing basis - Transitional|Transitional
Event|Activity|General Exam|11981,11986|false|false|false|C5966184|Issue (action)|issue
Event|Event|General Exam|11981,11986|false|false|false|||issue
Finding|Finding|General Exam|11981,11986|false|false|false|C0033213;C1706387|Issue (document);Problem|issue
Finding|Intellectual Product|General Exam|11981,11986|false|false|false|C0033213;C1706387|Issue (document);Problem|issue
Event|Event|General Exam|11991,11995|false|false|false|||goal
Finding|Idea or Concept|General Exam|11991,11995|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Finding|Intellectual Product|General Exam|11991,11995|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Event|Event|General Exam|12010,12016|false|false|false|||accord
Finding|Social Behavior|General Exam|12010,12016|false|false|false|C0680240|Agreement|accord
Anatomy|Body Part, Organ, or Organ Component|General Exam|12037,12040|false|false|false|C0152325;C2954192|Gray matter of anterior cingulate gyrus;Structure of forceps minor|ACC
Anatomy|Tissue|General Exam|12037,12040|false|false|false|C0152325;C2954192|Gray matter of anterior cingulate gyrus;Structure of forceps minor|ACC
Disorder|Congenital Abnormality|General Exam|12037,12040|false|false|false|C0175754;C0206686;C0282160|Adrenocortical carcinoma;Agenesis of corpus callosum;Aplasia Cutis Congenita|ACC
Disorder|Neoplastic Process|General Exam|12037,12040|false|false|false|C0175754;C0206686;C0282160|Adrenocortical carcinoma;Agenesis of corpus callosum;Aplasia Cutis Congenita|ACC
Drug|Amino Acid, Peptide, or Protein|General Exam|12037,12040|false|false|false|C3541857;C4724142|Acetyl-CoA Carboxylase 1;Amorphous Calcium Carbonate|ACC
Drug|Enzyme|General Exam|12037,12040|false|false|false|C3541857;C4724142|Acetyl-CoA Carboxylase 1;Amorphous Calcium Carbonate|ACC
Drug|Pharmacologic Substance|General Exam|12037,12040|false|false|false|C3541857;C4724142|Acetyl-CoA Carboxylase 1;Amorphous Calcium Carbonate|ACC
Event|Event|General Exam|12037,12040|false|false|false|||ACC
Finding|Gene or Genome|General Exam|12037,12040|false|false|false|C1412104;C3541413|ACACA gene;ACACA wt Allele|ACC
Disorder|Disease or Syndrome|General Exam|12041,12044|false|false|false|C0002880;C0272325|Autoimmune hemolytic anemia;Factor 8 deficiency, acquired|AHA
Drug|Organic Chemical|General Exam|12041,12044|false|false|false|C0050451|acetohydroxamic acid|AHA
Drug|Pharmacologic Substance|General Exam|12041,12044|false|false|false|C0050451|acetohydroxamic acid|AHA
Event|Event|General Exam|12041,12044|false|false|false|||AHA
Event|Event|General Exam|12049,12059|false|false|false|||guidelines
Finding|Intellectual Product|General Exam|12049,12059|false|false|false|C0162791;C0220845;C0282423|Guideline (Publication Type);Guidelines;guiding characteristics|guidelines
Event|Event|General Exam|12079,12089|false|false|false|||difficulty
Finding|Finding|General Exam|12079,12089|false|true|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Finding|Functional Concept|General Exam|12101,12111|false|false|false|C1524062|Additional|additional
Event|Event|General Exam|12112,12118|false|false|false|||agents
Disorder|Disease or Syndrome|General Exam|12123,12126|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Event|Event|General Exam|12123,12126|false|false|false|||CKD
Finding|Functional Concept|General Exam|12128,12134|false|false|false|C0439801|Limited (extensiveness)|limits
Event|Event|General Exam|12135,12138|false|false|false|||use
Finding|Functional Concept|General Exam|12135,12138|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|General Exam|12135,12138|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Functional Concept|General Exam|12135,12141|false|false|false|C1524063|Use of|use of
Drug|Organic Chemical|General Exam|12142,12151|false|false|false|C0009014|clonidine|clonidine
Drug|Pharmacologic Substance|General Exam|12142,12151|false|false|false|C0009014|clonidine|clonidine
Event|Event|General Exam|12142,12151|false|false|false|||clonidine
Drug|Biomedical or Dental Material|General Exam|12158,12166|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|General Exam|12158,12166|false|false|false|||baseline
Finding|Idea or Concept|General Exam|12158,12166|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Drug|Biologically Active Substance|General Exam|12167,12176|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Element, Ion, or Isotope|General Exam|12167,12176|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Food|General Exam|12167,12176|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Inorganic Chemical|General Exam|12167,12176|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Pharmacologic Substance|General Exam|12167,12176|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Event|Event|General Exam|12167,12176|false|false|false|||potassium
Finding|Physiologic Function|General Exam|12167,12176|false|false|false|C4553027|Potassium metabolic function|potassium
Procedure|Laboratory Procedure|General Exam|12167,12176|false|false|false|C0202194|Potassium measurement|potassium
Finding|Finding|General Exam|12184,12190|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|General Exam|12184,12190|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|General Exam|12191,12196|false|false|false|||limit
Drug|Organic Chemical|General Exam|12205,12219|false|false|false|C0037982|spironolactone|spironolactone
Drug|Pharmacologic Substance|General Exam|12205,12219|false|false|false|C0037982|spironolactone|spironolactone
Event|Event|General Exam|12205,12219|false|false|false|||spironolactone
Event|Event|General Exam|12224,12227|false|false|false|||TTE
Procedure|Diagnostic Procedure|General Exam|12224,12227|false|false|false|C0430462|Transthoracic echocardiography|TTE
Event|Event|General Exam|12228,12234|false|false|false|||showed
Event|Event|General Exam|12244,12255|false|false|false|||hypokinesis
Finding|Finding|General Exam|12244,12255|false|false|false|C0086439|Hypokinesia|hypokinesis
Event|Event|General Exam|12263,12271|false|false|false|||consider
Event|Event|General Exam|12272,12276|false|false|false|||MIBI
Procedure|Laboratory Procedure|General Exam|12272,12276|false|false|false|C5557372|Multiplexed Ion Beam Imaging|MIBI
Event|Event|General Exam|12281,12291|false|false|false|||outpatient
Finding|Classification|General Exam|12281,12291|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|General Exam|12281,12291|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Functional Concept|General Exam|12292,12307|false|false|false|C0205464|pharmacological|pharmacological
Phenomenon|Phenomenon or Process|General Exam|12292,12314|false|false|false|C0449421|Pharmacological stress|pharmacological stress
Attribute|Clinical Attribute|General Exam|12308,12314|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|General Exam|12308,12314|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|General Exam|12308,12314|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Event|Event|General Exam|12308,12314|false|false|false|||stress
Finding|Finding|General Exam|12308,12314|false|false|false|C0038435|Stress|stress
Procedure|Diagnostic Procedure|General Exam|12308,12319|false|false|false|C0015260;C3494508|Exercise stress test;Stress Test|stress test
Anatomy|Body Location or Region|General Exam|12315,12319|false|false|false|C4318744|Test - temporal region|test
Event|Event|General Exam|12315,12319|false|false|false|||test
Finding|Functional Concept|General Exam|12315,12319|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|General Exam|12315,12319|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|General Exam|12315,12319|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|General Exam|12315,12319|false|false|false|C0022885|Laboratory Procedures|test
Anatomy|Body Part, Organ, or Organ Component|General Exam|12331,12338|false|false|false|C0042027|Urinary tract|urinary
Attribute|Clinical Attribute|General Exam|12331,12348|false|false|false|C5700171|Bladder retention of urine|urinary retention
Finding|Functional Concept|General Exam|12331,12348|false|false|false|C0080274|Urinary Retention|urinary retention
Attribute|Clinical Attribute|General Exam|12339,12348|false|false|false|C1318143|Retention - dental|retention
Event|Event|General Exam|12339,12348|false|false|false|||retention
Finding|Cell Function|General Exam|12339,12348|false|false|false|C0035280;C0080274;C0333117;C1753315|Retention (Psychology);Retention of content;Urinary Retention;cellular entity retention|retention
Finding|Functional Concept|General Exam|12339,12348|false|false|false|C0035280;C0080274;C0333117;C1753315|Retention (Psychology);Retention of content;Urinary Retention;cellular entity retention|retention
Finding|Mental Process|General Exam|12339,12348|false|false|false|C0035280;C0080274;C0333117;C1753315|Retention (Psychology);Retention of content;Urinary Retention;cellular entity retention|retention
Disorder|Disease or Syndrome|General Exam|12349,12361|false|false|false|C0021167|Incontinence|incontinence
Event|Event|General Exam|12349,12361|false|false|false|||incontinence
Event|Event|General Exam|12383,12391|false|false|false|||diuresis
Finding|Organ or Tissue Function|General Exam|12383,12391|false|false|false|C0012797|Diuresis|diuresis
Event|Event|General Exam|12398,12404|false|false|false|||assess
Event|Event|General Exam|12419,12427|false|false|false|||symptoms
Finding|Functional Concept|General Exam|12419,12427|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|General Exam|12419,12427|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|General Exam|12431,12438|false|false|false|||routine
Finding|Idea or Concept|General Exam|12431,12438|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|routine
Finding|Intellectual Product|General Exam|12431,12438|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|routine
Procedure|Laboratory Procedure|General Exam|12431,12438|false|false|false|C1979801|Routine coag|routine
Finding|Classification|General Exam|12440,12450|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|General Exam|12440,12450|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Procedure|Health Care Activity|General Exam|12440,12457|false|false|false|C0545084|Outpatient visits|outpatient visits
Event|Event|General Exam|12451,12457|false|false|false|||visits
Finding|Social Behavior|General Exam|12451,12457|false|false|false|C0545082|Visit|visits
Procedure|Health Care Activity|General Exam|12451,12457|false|false|false|C1512346|Patient Visit|visits
Event|Event|General Exam|12460,12464|false|false|false|||CODE
Event|Occupational Activity|General Exam|12460,12464|false|false|false|C0009219|Coding|CODE
Finding|Intellectual Product|General Exam|12460,12464|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|CODE
Event|Event|General Exam|12472,12481|false|false|false|||confirmed
Event|Activity|General Exam|12486,12493|false|false|false|C3812666|Personal Contact|CONTACT
Event|Event|General Exam|12486,12493|false|false|false|||CONTACT
Finding|Functional Concept|General Exam|12486,12493|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Idea or Concept|General Exam|12486,12493|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Intellectual Product|General Exam|12486,12493|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Phenomenon|Phenomenon or Process|General Exam|12486,12493|false|false|false|C0392367|Physical contact|CONTACT
Attribute|Clinical Attribute|General Exam|12515,12526|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|General Exam|12515,12526|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|General Exam|12515,12526|false|false|false|||Medications
Finding|Intellectual Product|General Exam|12515,12526|false|false|false|C4284232|Medications|Medications
Finding|Finding|General Exam|12515,12539|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|General Exam|12530,12539|false|false|false|||Admission
Procedure|Health Care Activity|General Exam|12530,12539|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|General Exam|12558,12568|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|General Exam|12558,12568|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|General Exam|12558,12573|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|General Exam|12569,12573|false|false|false|||list
Finding|Intellectual Product|General Exam|12569,12573|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|General Exam|12577,12585|false|false|false|||accurate
Drug|Organic Chemical|General Exam|12590,12598|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|General Exam|12590,12598|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|General Exam|12590,12598|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|General Exam|12590,12598|false|false|false|||complete
Finding|Functional Concept|General Exam|12590,12598|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|General Exam|12590,12598|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|General Exam|12603,12614|false|false|false|C0002144|allopurinol|Allopurinol
Drug|Pharmacologic Substance|General Exam|12603,12614|false|false|false|C0002144|allopurinol|Allopurinol
Event|Event|General Exam|12637,12640|false|false|false|||DAY
Finding|Idea or Concept|General Exam|12637,12640|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|DAY
Finding|Intellectual Product|General Exam|12637,12640|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|DAY
Drug|Organic Chemical|General Exam|12645,12657|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|General Exam|12645,12657|false|false|false|C0286651|atorvastatin|Atorvastatin
Event|Event|General Exam|12667,12670|false|false|false|||QPM
Drug|Organic Chemical|General Exam|12675,12685|false|false|false|C0006674;C3714610|Calcitriol Drug Class;calcitriol|Calcitriol
Drug|Pharmacologic Substance|General Exam|12675,12685|false|false|false|C0006674;C3714610|Calcitriol Drug Class;calcitriol|Calcitriol
Drug|Vitamin|General Exam|12675,12685|false|false|false|C0006674;C3714610|Calcitriol Drug Class;calcitriol|Calcitriol
Event|Event|General Exam|12675,12685|false|false|false|||Calcitriol
Drug|Organic Chemical|General Exam|12707,12717|false|false|false|C0054836|carvedilol|Carvedilol
Drug|Pharmacologic Substance|General Exam|12707,12717|false|false|false|C0054836|carvedilol|Carvedilol
Disorder|Mental or Behavioral Dysfunction|General Exam|12727,12730|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|General Exam|12727,12730|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|General Exam|12727,12730|false|false|false|C1530795|BID protein, human|BID
Event|Event|General Exam|12727,12730|false|false|false|||BID
Finding|Gene or Genome|General Exam|12727,12730|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|General Exam|12735,12745|false|false|false|C0060926|gabapentin|Gabapentin
Drug|Pharmacologic Substance|General Exam|12735,12745|false|false|false|C0060926|gabapentin|Gabapentin
Drug|Organic Chemical|General Exam|12764,12774|false|false|false|C0028066|nifedipine|NIFEdipine
Drug|Pharmacologic Substance|General Exam|12764,12774|false|false|false|C0028066|nifedipine|NIFEdipine
Event|Event|General Exam|12764,12774|false|false|false|||NIFEdipine
Finding|Finding|General Exam|12776,12784|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|General Exam|12776,12784|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|General Exam|12785,12792|false|false|false|||Release
Finding|Functional Concept|General Exam|12785,12792|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|General Exam|12785,12792|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|General Exam|12785,12792|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Disorder|Mental or Behavioral Dysfunction|General Exam|12803,12806|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|General Exam|12803,12806|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|General Exam|12803,12806|false|false|false|C1530795|BID protein, human|BID
Event|Event|General Exam|12803,12806|false|false|false|||BID
Finding|Gene or Genome|General Exam|12803,12806|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|General Exam|12811,12820|false|false|false|C0076840|torsemide|Torsemide
Drug|Pharmacologic Substance|General Exam|12811,12820|false|false|false|C0076840|torsemide|Torsemide
Drug|Organic Chemical|General Exam|12840,12853|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Pharmacologic Substance|General Exam|12840,12853|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Event|Event|General Exam|12840,12853|false|false|false|||Nitroglycerin
Finding|Gene or Genome|General Exam|12873,12876|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Location or Region|General Exam|12877,12882|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|General Exam|12877,12882|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|General Exam|12877,12887|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|General Exam|12877,12887|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|General Exam|12883,12887|false|false|false|C2598155||pain
Event|Event|General Exam|12883,12887|false|false|false|||pain
Finding|Functional Concept|General Exam|12883,12887|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|General Exam|12883,12887|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|General Exam|12892,12905|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|General Exam|12892,12905|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|General Exam|12892,12905|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|General Exam|12892,12905|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|General Exam|12924,12927|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|General Exam|12928,12932|false|false|false|C2598155||Pain
Event|Event|General Exam|12928,12932|false|false|false|||Pain
Finding|Functional Concept|General Exam|12928,12932|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|General Exam|12928,12932|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Intellectual Product|General Exam|12935,12939|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Drug|Organic Chemical|General Exam|12945,12952|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|General Exam|12945,12952|false|false|false|C0004057|aspirin|Aspirin
Drug|Amino Acid, Peptide, or Protein|General Exam|12973,12980|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Hormone|General Exam|12973,12980|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Pharmacologic Substance|General Exam|12973,12980|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Event|Event|General Exam|12973,12980|false|false|false|||Insulin
Finding|Gene or Genome|General Exam|12973,12980|false|false|false|C1337112|INS gene|Insulin
Procedure|Laboratory Procedure|General Exam|12973,12980|false|false|false|C0202098|Insulin measurement|Insulin
Finding|Functional Concept|General Exam|12991,12998|false|false|false|C0332246|Sliding|Sliding
Procedure|Therapeutic or Preventive Procedure|General Exam|12991,13004|false|false|false|C2937251|sliding scale|Sliding Scale
Anatomy|Body Part, Organ, or Organ Component|General Exam|12999,13004|false|false|false|C0222045|Integumentary scale|Scale
Event|Activity|General Exam|12999,13004|false|false|false|C1947916|Scaling|Scale
Finding|Conceptual Entity|General Exam|12999,13004|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|Scale
Finding|Intellectual Product|General Exam|12999,13004|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|Scale
Drug|Amino Acid, Peptide, or Protein|General Exam|13005,13012|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Hormone|General Exam|13005,13012|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Pharmacologic Substance|General Exam|13005,13012|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Event|Event|General Exam|13005,13012|false|false|false|||Insulin
Finding|Gene or Genome|General Exam|13005,13012|false|false|false|C1337112|INS gene|Insulin
Procedure|Laboratory Procedure|General Exam|13005,13012|false|false|false|C0202098|Insulin measurement|Insulin
Finding|Functional Concept|General Exam|13016,13023|false|false|false|C0332246|Sliding|Sliding
Procedure|Therapeutic or Preventive Procedure|General Exam|13016,13029|false|false|false|C2937251|sliding scale|Sliding Scale
Anatomy|Body Part, Organ, or Organ Component|General Exam|13024,13029|false|false|false|C0222045|Integumentary scale|Scale
Event|Activity|General Exam|13024,13029|false|false|false|C1947916|Scaling|Scale
Event|Event|General Exam|13024,13029|false|false|false|||Scale
Finding|Conceptual Entity|General Exam|13024,13029|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|Scale
Finding|Intellectual Product|General Exam|13024,13029|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|Scale
Drug|Amino Acid, Peptide, or Protein|General Exam|13042,13049|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Hormone|General Exam|13042,13049|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Pharmacologic Substance|General Exam|13042,13049|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Event|Event|General Exam|13042,13049|false|false|false|||Insulin
Finding|Gene or Genome|General Exam|13042,13049|false|false|false|C1337112|INS gene|Insulin
Procedure|Laboratory Procedure|General Exam|13042,13049|false|false|false|C0202098|Insulin measurement|Insulin
Event|Event|General Exam|13053,13062|false|false|false|||Discharge
Finding|Body Substance|General Exam|13053,13062|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|General Exam|13053,13062|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|General Exam|13053,13062|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|General Exam|13053,13062|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|General Exam|13053,13074|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|General Exam|13063,13074|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|General Exam|13063,13074|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|General Exam|13063,13074|false|false|false|||Medications
Finding|Intellectual Product|General Exam|13063,13074|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|General Exam|13080,13093|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|General Exam|13080,13093|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|General Exam|13080,13093|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|General Exam|13080,13093|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|General Exam|13112,13115|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|General Exam|13116,13120|false|false|false|C2598155||Pain
Event|Event|General Exam|13116,13120|false|false|false|||Pain
Finding|Functional Concept|General Exam|13116,13120|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|General Exam|13116,13120|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Intellectual Product|General Exam|13123,13127|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Drug|Organic Chemical|General Exam|13134,13145|false|false|false|C0002144|allopurinol|Allopurinol
Drug|Pharmacologic Substance|General Exam|13134,13145|false|false|false|C0002144|allopurinol|Allopurinol
Event|Event|General Exam|13168,13171|false|false|false|||DAY
Finding|Idea or Concept|General Exam|13168,13171|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|DAY
Finding|Intellectual Product|General Exam|13168,13171|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|DAY
Drug|Organic Chemical|General Exam|13178,13185|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|General Exam|13178,13185|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|General Exam|13207,13219|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|General Exam|13207,13219|false|false|false|C0286651|atorvastatin|Atorvastatin
Event|Event|General Exam|13229,13232|false|false|false|||QPM
Drug|Organic Chemical|General Exam|13239,13249|false|false|false|C0006674;C3714610|Calcitriol Drug Class;calcitriol|Calcitriol
Drug|Pharmacologic Substance|General Exam|13239,13249|false|false|false|C0006674;C3714610|Calcitriol Drug Class;calcitriol|Calcitriol
Drug|Vitamin|General Exam|13239,13249|false|false|false|C0006674;C3714610|Calcitriol Drug Class;calcitriol|Calcitriol
Drug|Organic Chemical|General Exam|13273,13283|false|false|false|C0054836|carvedilol|Carvedilol
Drug|Pharmacologic Substance|General Exam|13273,13283|false|false|false|C0054836|carvedilol|Carvedilol
Disorder|Mental or Behavioral Dysfunction|General Exam|13293,13296|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|General Exam|13293,13296|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|General Exam|13293,13296|false|false|false|C1530795|BID protein, human|BID
Event|Event|General Exam|13293,13296|false|false|false|||BID
Finding|Gene or Genome|General Exam|13293,13296|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|General Exam|13303,13313|false|false|false|C0060926|gabapentin|Gabapentin
Drug|Pharmacologic Substance|General Exam|13303,13313|false|false|false|C0060926|gabapentin|Gabapentin
Drug|Amino Acid, Peptide, or Protein|General Exam|13334,13341|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Hormone|General Exam|13334,13341|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Pharmacologic Substance|General Exam|13334,13341|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Event|Event|General Exam|13334,13341|false|false|false|||Insulin
Finding|Gene or Genome|General Exam|13334,13341|false|false|false|C1337112|INS gene|Insulin
Procedure|Laboratory Procedure|General Exam|13334,13341|false|false|false|C0202098|Insulin measurement|Insulin
Finding|Functional Concept|General Exam|13352,13359|false|false|false|C0332246|Sliding|Sliding
Procedure|Therapeutic or Preventive Procedure|General Exam|13352,13365|false|false|false|C2937251|sliding scale|Sliding Scale
Anatomy|Body Part, Organ, or Organ Component|General Exam|13360,13365|false|false|false|C0222045|Integumentary scale|Scale
Event|Activity|General Exam|13360,13365|false|false|false|C1947916|Scaling|Scale
Finding|Conceptual Entity|General Exam|13360,13365|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|Scale
Finding|Intellectual Product|General Exam|13360,13365|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|Scale
Drug|Amino Acid, Peptide, or Protein|General Exam|13366,13373|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Hormone|General Exam|13366,13373|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Pharmacologic Substance|General Exam|13366,13373|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Event|Event|General Exam|13366,13373|false|false|false|||Insulin
Finding|Gene or Genome|General Exam|13366,13373|false|false|false|C1337112|INS gene|Insulin
Procedure|Laboratory Procedure|General Exam|13366,13373|false|false|false|C0202098|Insulin measurement|Insulin
Finding|Functional Concept|General Exam|13377,13384|false|false|false|C0332246|Sliding|Sliding
Procedure|Therapeutic or Preventive Procedure|General Exam|13377,13390|false|false|false|C2937251|sliding scale|Sliding Scale
Anatomy|Body Part, Organ, or Organ Component|General Exam|13385,13390|false|false|false|C0222045|Integumentary scale|Scale
Event|Activity|General Exam|13385,13390|false|false|false|C1947916|Scaling|Scale
Event|Event|General Exam|13385,13390|false|false|false|||Scale
Finding|Conceptual Entity|General Exam|13385,13390|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|Scale
Finding|Intellectual Product|General Exam|13385,13390|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|Scale
Drug|Amino Acid, Peptide, or Protein|General Exam|13403,13410|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Hormone|General Exam|13403,13410|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Pharmacologic Substance|General Exam|13403,13410|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Event|Event|General Exam|13403,13410|false|false|false|||Insulin
Finding|Gene or Genome|General Exam|13403,13410|false|false|false|C1337112|INS gene|Insulin
Procedure|Laboratory Procedure|General Exam|13403,13410|false|false|false|C0202098|Insulin measurement|Insulin
Drug|Organic Chemical|General Exam|13416,13426|false|false|false|C0028066|nifedipine|NIFEdipine
Drug|Pharmacologic Substance|General Exam|13416,13426|false|false|false|C0028066|nifedipine|NIFEdipine
Event|Event|General Exam|13416,13426|false|false|false|||NIFEdipine
Finding|Finding|General Exam|13428,13436|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|General Exam|13428,13436|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|General Exam|13437,13444|false|false|false|||Release
Finding|Functional Concept|General Exam|13437,13444|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|General Exam|13437,13444|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|General Exam|13437,13444|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Disorder|Mental or Behavioral Dysfunction|General Exam|13455,13458|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|General Exam|13455,13458|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|General Exam|13455,13458|false|false|false|C1530795|BID protein, human|BID
Event|Event|General Exam|13455,13458|false|false|false|||BID
Finding|Gene or Genome|General Exam|13455,13458|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|General Exam|13466,13479|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Pharmacologic Substance|General Exam|13466,13479|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Event|Event|General Exam|13466,13479|false|false|false|||Nitroglycerin
Finding|Gene or Genome|General Exam|13499,13502|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Location or Region|General Exam|13503,13508|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|General Exam|13503,13508|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|General Exam|13503,13513|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|General Exam|13503,13513|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|General Exam|13509,13513|false|true|false|C2598155||pain
Event|Event|General Exam|13509,13513|false|false|false|||pain
Finding|Functional Concept|General Exam|13509,13513|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|General Exam|13509,13513|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|General Exam|13521,13530|false|false|false|C0076840|torsemide|Torsemide
Drug|Pharmacologic Substance|General Exam|13521,13530|false|false|false|C0076840|torsemide|Torsemide
Event|Event|General Exam|13551,13560|false|false|false|||Discharge
Finding|Body Substance|General Exam|13551,13560|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|General Exam|13551,13560|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|General Exam|13551,13560|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|General Exam|13551,13560|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|General Exam|13551,13572|false|false|false|C4019243||Discharge Disposition
Finding|Finding|General Exam|13551,13572|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|General Exam|13561,13572|false|false|false|C2926604||Disposition
Event|Event|General Exam|13561,13572|false|false|false|||Disposition
Procedure|Health Care Activity|General Exam|13561,13572|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|General Exam|13574,13578|false|false|false|||Home
Finding|Idea or Concept|General Exam|13574,13578|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|General Exam|13574,13578|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|General Exam|13574,13578|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|General Exam|13584,13591|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|General Exam|13584,13591|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|General Exam|13594,13602|false|false|false|||Facility
Finding|Intellectual Product|General Exam|13594,13602|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|General Exam|13610,13619|false|false|false|||Discharge
Finding|Body Substance|General Exam|13610,13619|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|General Exam|13610,13619|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|General Exam|13610,13619|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|General Exam|13610,13619|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|General Exam|13610,13629|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|General Exam|13620,13629|false|false|false|C0945731||Diagnosis
Event|Event|General Exam|13620,13629|false|false|false|||Diagnosis
Finding|Classification|General Exam|13620,13629|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|General Exam|13620,13629|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|General Exam|13620,13629|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Intellectual Product|Principle Diagnosis|13651,13656|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Disorder|Disease or Syndrome|Principle Diagnosis|13651,13702|false|false|false|C2732749|Acute on chronic diastolic heart failure|Acute on chronic diastolic congestive heart failure
Finding|Intellectual Product|Principle Diagnosis|13660,13667|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Principle Diagnosis|13660,13667|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|Principle Diagnosis|13660,13702|false|false|false|C2711480|Chronic diastolic heart failure|chronic diastolic congestive heart failure
Attribute|Clinical Attribute|Principle Diagnosis|13668,13677|false|false|false|C0012000|Diastole|diastolic
Disorder|Disease or Syndrome|Principle Diagnosis|13668,13702|false|false|false|C2183328|diastolic congestive heart failure|diastolic congestive heart failure
Disorder|Disease or Syndrome|Principle Diagnosis|13678,13702|false|false|false|C0018802|Congestive heart failure|congestive heart failure
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|13689,13694|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Principle Diagnosis|13689,13694|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Principle Diagnosis|13689,13694|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|Principle Diagnosis|13689,13702|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Event|Event|Principle Diagnosis|13695,13702|false|false|false|||failure
Finding|Functional Concept|Principle Diagnosis|13695,13702|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|Principle Diagnosis|13695,13702|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|Principle Diagnosis|13695,13702|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Disorder|Neoplastic Process|Principle Diagnosis|13704,13713|false|false|false|C0027627|Neoplasm Metastasis|SECONDARY
Finding|Functional Concept|Principle Diagnosis|13704,13713|false|false|false|C1522484|metastatic qualifier|SECONDARY
Procedure|Diagnostic Procedure|Principle Diagnosis|13714,13723|false|false|false|C0011900|Diagnosis|DIAGNOSES
Disorder|Disease or Syndrome|Principle Diagnosis|13726,13738|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|Principle Diagnosis|13726,13738|false|false|false|||Hypertension
Event|Event|Principle Diagnosis|13741,13748|false|false|false|||History
Finding|Conceptual Entity|Principle Diagnosis|13741,13748|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|Principle Diagnosis|13741,13748|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|Principle Diagnosis|13741,13748|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|Principle Diagnosis|13741,13751|false|false|false|C0262926|Medical History|History of
Anatomy|Body Location or Region|Principle Diagnosis|13758,13761|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Principle Diagnosis|13758,13761|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Principle Diagnosis|13758,13761|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|Principle Diagnosis|13758,13761|false|false|false|||DVT
Disorder|Disease or Syndrome|Principle Diagnosis|13764,13770|false|false|false|C0002871|Anemia|Anemia
Event|Event|Principle Diagnosis|13764,13770|false|false|false|||Anemia
Event|Event|Principle Diagnosis|13772,13775|false|false|false|||NOS
Finding|Intellectual Product|Principle Diagnosis|13778,13785|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|Principle Diagnosis|13778,13785|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Disorder|Disease or Syndrome|Principle Diagnosis|13778,13800|false|false|false|C1561643|Chronic Kidney Diseases|Chronic Kidney Disease
Finding|Classification|Principle Diagnosis|13778,13806|false|false|false|C2074731|chronic kidney disease stage|Chronic Kidney Disease stage
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|13786,13792|false|false|false|C0022646;C0227665|Both kidneys;Kidney|Kidney
Disorder|Neoplastic Process|Principle Diagnosis|13786,13792|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|Kidney
Event|Event|Principle Diagnosis|13786,13792|false|false|false|||Kidney
Finding|Sign or Symptom|Principle Diagnosis|13786,13792|false|false|false|C0812426|Kidney problem|Kidney
Procedure|Diagnostic Procedure|Principle Diagnosis|13786,13792|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|Kidney
Procedure|Therapeutic or Preventive Procedure|Principle Diagnosis|13786,13792|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|Kidney
Disorder|Disease or Syndrome|Principle Diagnosis|13786,13800|false|false|false|C0022658|Kidney Diseases|Kidney Disease
Disorder|Disease or Syndrome|Principle Diagnosis|13793,13800|false|false|false|C0012634|Disease|Disease
Attribute|Clinical Attribute|Principle Diagnosis|13793,13806|false|false|false|C0699749;C3260349|disease stage|Disease stage
Attribute|Clinical Attribute|Principle Diagnosis|13801,13806|false|false|false|C1300072|Tumor stage|stage
Event|Event|Principle Diagnosis|13801,13806|false|false|false|||stage
Finding|Intellectual Product|Principle Diagnosis|13801,13809|false|false|false|C0441772|Stage level 4|stage IV
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|13812,13820|false|false|false|C0018787|Heart|Coronary
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|13812,13827|false|false|false|C0205042|Coronary artery|Coronary Artery
Disorder|Disease or Syndrome|Principle Diagnosis|13812,13835|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|Coronary Artery Disease
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|13821,13827|false|false|false|C0003842;C0226004|Arterial system;Arteries|Artery
Anatomy|Body System|Principle Diagnosis|13821,13827|false|false|false|C0003842;C0226004|Arterial system;Arteries|Artery
Disorder|Disease or Syndrome|Principle Diagnosis|13821,13835|false|false|false|C0852949|Arteriopathic disease|Artery Disease
Disorder|Disease or Syndrome|Principle Diagnosis|13828,13835|false|false|false|C0012634|Disease|Disease
Event|Event|Principle Diagnosis|13828,13835|false|false|false|||Disease
Drug|Pharmacologic Substance|Principle Diagnosis|13840,13844|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|drug
Finding|Finding|Principle Diagnosis|13840,13844|false|false|false|C0740721|Drug problem|drug
Event|Event|Principle Diagnosis|13853,13858|false|false|false|||stent
Disorder|Disease or Syndrome|Principle Diagnosis|13861,13869|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|Diabetes
Disorder|Disease or Syndrome|Principle Diagnosis|13861,13878|false|false|false|C0011849|Diabetes Mellitus|Diabetes Mellitus
Disorder|Disease or Syndrome|Principle Diagnosis|13861,13885|false|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|Diabetes Mellitus Type 2
Finding|Gene or Genome|Principle Diagnosis|13879,13883|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|Type
Finding|Intellectual Product|Principle Diagnosis|13879,13883|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|Type
Finding|Classification|Principle Diagnosis|13879,13885|false|false|false|C0441730|Type 2|Type 2
Event|Event|Principle Diagnosis|13886,13896|false|false|false|||controlled
Finding|Finding|Principle Diagnosis|13886,13896|false|false|false|C2587213;C2911690;C4761797|Control function;Controlled mark;Disease Controlled|controlled
Finding|Functional Concept|Principle Diagnosis|13886,13896|false|false|false|C2587213;C2911690;C4761797|Control function;Controlled mark;Disease Controlled|controlled
Finding|Idea or Concept|Principle Diagnosis|13886,13896|false|false|false|C2587213;C2911690;C4761797|Control function;Controlled mark;Disease Controlled|controlled
Finding|Mental Process|Discharge Condition|13921,13927|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|13921,13934|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|13921,13934|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|13928,13934|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|13928,13934|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|13936,13941|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|13936,13941|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|13946,13954|false|false|false|||coherent
Finding|Finding|Discharge Condition|13946,13954|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|13956,13961|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|13956,13978|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|13956,13978|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|13965,13978|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|13965,13978|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|13965,13978|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|13980,13985|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|13980,13985|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|13980,13985|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|13980,13985|false|false|false|||Alert
Finding|Finding|Discharge Condition|13980,13985|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|13980,13985|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|13980,13985|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|13990,14001|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|13990,14001|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|14003,14011|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|14003,14011|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|14003,14011|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|14012,14018|false|false|false|C5889824||Status
Event|Event|Discharge Condition|14012,14018|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|14012,14018|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|14020,14030|false|false|false|||Ambulatory
Finding|Functional Concept|Discharge Condition|14020,14030|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|14020,14030|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|14020,14030|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|14020,14030|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|14033,14044|false|false|false|||Independent
Finding|Finding|Discharge Condition|14033,14044|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Condition|14033,14044|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Gene or Genome|Discharge Instructions|14073,14077|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|Discharge Instructions|14093,14101|false|false|false|||admitted
Finding|Idea or Concept|Discharge Instructions|14109,14117|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|Discharge Instructions|14123,14132|false|false|false|||shortness
Attribute|Clinical Attribute|Discharge Instructions|14123,14142|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|Discharge Instructions|14123,14142|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|Discharge Instructions|14136,14142|false|false|false|C0225386|Breath|breath
Attribute|Clinical Attribute|Discharge Instructions|14148,14154|false|false|false|C0944911||weight
Event|Event|Discharge Instructions|14148,14154|false|false|false|||weight
Finding|Finding|Discharge Instructions|14148,14154|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|Discharge Instructions|14148,14154|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|Discharge Instructions|14148,14154|false|false|false|C1305866|Weighing patient|weight
Finding|Finding|Discharge Instructions|14148,14159|false|false|false|C0043094;C3814804|Gaining Weight question;Weight Gain|weight gain
Finding|Intellectual Product|Discharge Instructions|14148,14159|false|false|false|C0043094;C3814804|Gaining Weight question;Weight Gain|weight gain
Event|Event|Discharge Instructions|14155,14159|false|false|false|||gain
Finding|Finding|Discharge Instructions|14171,14177|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Discharge Instructions|14171,14177|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|Discharge Instructions|14178,14184|false|false|false|||caused
Event|Event|Discharge Instructions|14191,14203|false|false|false|||exacerbation
Finding|Finding|Discharge Instructions|14191,14203|false|false|false|C4086268|Exacerbation|exacerbation
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|14213,14218|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|14213,14218|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Discharge Instructions|14213,14218|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|Discharge Instructions|14213,14226|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Event|Event|Discharge Instructions|14219,14226|false|false|false|||failure
Finding|Functional Concept|Discharge Instructions|14219,14226|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|Discharge Instructions|14219,14226|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|Discharge Instructions|14219,14226|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Finding|Discharge Instructions|14227,14235|false|false|false|C0332149|Possible|possibly
Drug|Food|Discharge Instructions|14247,14252|false|false|false|C0016452|Food|foods
Event|Event|Discharge Instructions|14247,14252|false|false|false|||foods
Event|Event|Discharge Instructions|14262,14269|false|false|false|||holiday
Event|Event|Discharge Instructions|14262,14269|false|false|false|C0019843|Holidays|holiday
Finding|Idea or Concept|Discharge Instructions|14295,14303|false|false|false|C1547192|Organization unit type - Hospital|hospital
Drug|Pharmacologic Substance|Discharge Instructions|14322,14331|false|false|false|C0012798|Diuretics|diuretics
Event|Event|Discharge Instructions|14322,14331|false|false|false|||diuretics
Event|Event|Discharge Instructions|14335,14339|false|false|false|||help
Event|Event|Discharge Instructions|14340,14346|false|false|false|||remove
Drug|Substance|Discharge Instructions|14353,14358|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|Discharge Instructions|14353,14358|false|false|false|||fluid
Finding|Intellectual Product|Discharge Instructions|14353,14358|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|Discharge Instructions|14364,14371|false|false|false|||checked
Disorder|Disease or Syndrome|Discharge Instructions|14376,14385|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|Discharge Instructions|14376,14385|false|false|false|||pneumonia
Anatomy|Body Location or Region|Discharge Instructions|14393,14398|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Discharge Instructions|14393,14398|true|false|false|C0741025|Chest problem|chest
Procedure|Diagnostic Procedure|Discharge Instructions|14393,14404|true|false|false|C0039985|Plain chest X-ray|chest x-ray
Event|Event|Discharge Instructions|14399,14404|true|false|false|||x-ray
Finding|Functional Concept|Discharge Instructions|14399,14404|true|false|false|C0034571;C3244296|ActClaimAttachmentCategoryCode - x-ray;roentgenographic|x-ray
Finding|Intellectual Product|Discharge Instructions|14399,14404|true|false|false|C0034571;C3244296|ActClaimAttachmentCategoryCode - x-ray;roentgenographic|x-ray
Phenomenon|Natural Phenomenon or Process|Discharge Instructions|14399,14404|true|false|false|C0043309|Roentgen Rays|x-ray
Procedure|Diagnostic Procedure|Discharge Instructions|14399,14404|true|false|false|C0043299;C1306645;C1962945|Diagnostic radiologic examination;Plain x-ray;Radiographic imaging procedure|x-ray
Event|Event|Discharge Instructions|14419,14423|true|false|false|||sign
Finding|Finding|Discharge Instructions|14419,14423|true|false|false|C0311392;C1547188|Language Ability - Sign;Physical findings|sign
Finding|Idea or Concept|Discharge Instructions|14419,14423|true|false|false|C0311392;C1547188|Language Ability - Sign;Physical findings|sign
Disorder|Disease or Syndrome|Discharge Instructions|14430,14439|true|false|false|C0032285|Pneumonia|pneumonia
Event|Event|Discharge Instructions|14430,14439|true|false|false|||pneumonia
Event|Event|Discharge Instructions|14445,14452|false|false|false|||checked
Event|Event|Discharge Instructions|14457,14462|false|false|false|||signs
Finding|Finding|Discharge Instructions|14457,14462|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Discharge Instructions|14457,14462|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Finding|Discharge Instructions|14466,14469|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Discharge Instructions|14466,14469|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Event|Event|Discharge Instructions|14470,14475|true|false|false|||clots
Finding|Pathologic Function|Discharge Instructions|14470,14475|true|false|false|C0302148|Blood Clot|clots
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|14484,14488|true|false|false|C1140621|Leg|legs
Attribute|Clinical Attribute|Discharge Instructions|14484,14488|true|false|false|C5781420||legs
Finding|Finding|Discharge Instructions|14504,14507|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Discharge Instructions|14504,14507|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Drug|Organic Chemical|Discharge Instructions|14508,14512|true|false|false|C0009074|clotrimazole|clot
Drug|Pharmacologic Substance|Discharge Instructions|14508,14512|true|false|false|C0009074|clotrimazole|clot
Event|Event|Discharge Instructions|14508,14512|true|false|false|||clot
Finding|Pathologic Function|Discharge Instructions|14508,14512|true|false|false|C0302148|Blood Clot|clot
Event|Event|Discharge Instructions|14537,14541|false|false|false|||home
Finding|Idea or Concept|Discharge Instructions|14537,14541|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Discharge Instructions|14537,14541|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Discharge Instructions|14537,14541|false|false|false|C1553498|home health encounter|home
Event|Event|Discharge Instructions|14545,14553|false|false|false|||continue
Finding|Idea or Concept|Discharge Instructions|14545,14553|false|false|false|C0549178|Continuous|continue
Event|Event|Discharge Instructions|14557,14561|false|false|false|||take
Attribute|Clinical Attribute|Discharge Instructions|14574,14585|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|14574,14585|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|14574,14585|false|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|14574,14585|false|false|false|C4284232|Medications|medications
Event|Event|Discharge Instructions|14589,14599|false|false|false|||prescribed
Event|Event|Discharge Instructions|14602,14609|false|false|false|||monitor
Drug|Chemical Viewed Structurally|Discharge Instructions|14615,14619|true|false|false|C0036140;C0037494;C0206136|Salts;Sodium Chloride, Dietary;sodium chloride|salt
Drug|Food|Discharge Instructions|14615,14619|true|false|false|C0036140;C0037494;C0206136|Salts;Sodium Chloride, Dietary;sodium chloride|salt
Drug|Inorganic Chemical|Discharge Instructions|14615,14619|true|false|false|C0036140;C0037494;C0206136|Salts;Sodium Chloride, Dietary;sodium chloride|salt
Event|Event|Discharge Instructions|14620,14626|true|false|false|||intake
Finding|Functional Concept|Discharge Instructions|14620,14626|true|false|false|C1512806|Intake|intake
Procedure|Health Care Activity|Discharge Instructions|14620,14626|true|false|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|intake
Finding|Idea or Concept|Discharge Instructions|14671,14674|true|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Discharge Instructions|14671,14674|true|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Discharge Instructions|14676,14679|false|false|false|||ask
Event|Event|Discharge Instructions|14685,14692|false|false|false|||doctors
Event|Event|Discharge Instructions|14697,14701|false|false|false|||help
Finding|Intellectual Product|Discharge Instructions|14697,14701|false|false|false|C1552861|Help document|help
Event|Event|Discharge Instructions|14727,14731|true|false|false|||know
Event|Event|Discharge Instructions|14739,14743|false|false|false|||keep
Drug|Chemical Viewed Structurally|Discharge Instructions|14758,14762|false|false|false|C0036140;C0037494;C0206136|Salts;Sodium Chloride, Dietary;sodium chloride|salt
Drug|Food|Discharge Instructions|14758,14762|false|false|false|C0036140;C0037494;C0206136|Salts;Sodium Chloride, Dietary;sodium chloride|salt
Drug|Inorganic Chemical|Discharge Instructions|14758,14762|false|false|false|C0036140;C0037494;C0206136|Salts;Sodium Chloride, Dietary;sodium chloride|salt
Event|Event|Discharge Instructions|14758,14762|false|false|false|||salt
Event|Event|Discharge Instructions|14765,14773|false|false|false|||continue
Finding|Idea or Concept|Discharge Instructions|14765,14773|false|false|false|C0549178|Continuous|continue
Event|Event|Discharge Instructions|14777,14782|false|false|false|||weigh
Event|Event|Discharge Instructions|14807,14811|false|false|false|||call
Finding|Intellectual Product|Discharge Instructions|14817,14823|false|false|false|C2348314|Doctor - Title|doctor
Attribute|Clinical Attribute|Discharge Instructions|14828,14834|false|false|false|C0944911||weight
Event|Event|Discharge Instructions|14828,14834|false|false|false|||weight
Finding|Finding|Discharge Instructions|14828,14834|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|Discharge Instructions|14828,14834|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|Discharge Instructions|14828,14834|false|false|false|C1305866|Weighing patient|weight
Event|Event|Discharge Instructions|14835,14839|false|false|false|||goes
Event|Event|Discharge Instructions|14855,14858|false|false|false|||lbs
Procedure|Laboratory Procedure|Discharge Instructions|14855,14858|false|false|false|C3161851|liquid-based cytology (procedure)|lbs
Event|Event|Discharge Instructions|14862,14868|false|false|false|||follow
Finding|Functional Concept|Discharge Instructions|14862,14868|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|Discharge Instructions|14862,14868|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|Discharge Instructions|14862,14871|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|Discharge Instructions|14862,14871|false|false|false|C1522577|follow-up|follow-up
Finding|Intellectual Product|Discharge Instructions|14882,14894|false|false|false|C1547426|Location Service Code - Primary Care|primary care
Procedure|Health Care Activity|Discharge Instructions|14882,14894|false|false|false|C0033137|Primary Health Care|primary care
Event|Activity|Discharge Instructions|14890,14894|false|false|false|C1947933|care activity|care
Event|Event|Discharge Instructions|14890,14894|false|false|false|||care
Finding|Finding|Discharge Instructions|14890,14894|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|14890,14894|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|14895,14901|false|false|false|C2348314|Doctor - Title|doctor
Disorder|Disease or Syndrome|Discharge Instructions|14917,14922|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Discharge Instructions|14917,14922|false|false|false|||blood
Finding|Body Substance|Discharge Instructions|14917,14922|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Event|Discharge Instructions|14924,14932|false|false|false|||pressure
Finding|Finding|Discharge Instructions|14924,14932|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|Discharge Instructions|14924,14932|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|Discharge Instructions|14924,14932|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|Discharge Instructions|14924,14932|false|false|false|C0033095||pressure
Disorder|Disease or Syndrome|Discharge Instructions|14937,14942|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Discharge Instructions|14937,14942|false|false|false|||blood
Finding|Body Substance|Discharge Instructions|14937,14942|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Organic Chemical|Discharge Instructions|14937,14948|false|false|false|C0005802|Blood Glucose|blood sugar
Procedure|Laboratory Procedure|Discharge Instructions|14937,14948|false|false|false|C0392201|Blood glucose measurement|blood sugar
Drug|Biomedical or Dental Material|Discharge Instructions|14943,14948|false|false|false|C0007004;C0242209;C3665462|Carbohydrates;Sugars;raw sugar|sugar
Drug|Organic Chemical|Discharge Instructions|14943,14948|false|false|false|C0007004;C0242209;C3665462|Carbohydrates;Sugars;raw sugar|sugar
Drug|Pharmacologic Substance|Discharge Instructions|14943,14948|false|false|false|C0007004;C0242209;C3665462|Carbohydrates;Sugars;raw sugar|sugar
Drug|Organic Chemical|Discharge Instructions|14949,14956|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|Discharge Instructions|14949,14956|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|Discharge Instructions|14949,14956|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Event|Event|Discharge Instructions|14949,14956|false|false|false|||control
Finding|Conceptual Entity|Discharge Instructions|14949,14956|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|Discharge Instructions|14949,14956|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|Discharge Instructions|14949,14956|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Event|Event|Discharge Instructions|14967,14975|false|false|false|||pleasure
Finding|Intellectual Product|Discharge Instructions|14967,14975|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|Discharge Instructions|14967,14975|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|Discharge Instructions|14983,14987|false|false|false|C1947933|care activity|care
Event|Event|Discharge Instructions|14983,14987|false|false|false|||care
Finding|Finding|Discharge Instructions|14983,14987|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|14983,14987|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|14983,14990|false|false|false|C1555558|care of - AddressPartType|care of
Event|Event|Discharge Instructions|15006,15015|false|false|false|||Inpatient
Finding|Idea or Concept|Discharge Instructions|15006,15015|false|false|false|C1548438;C1549404|Patient Class - Inpatient;Referral category - Inpatient|Inpatient
Procedure|Health Care Activity|Discharge Instructions|15006,15015|false|false|false|C1555324|inpatient encounter|Inpatient
Procedure|Health Care Activity|Discharge Instructions|15006,15020|false|false|false|C0019993|Hospitalization|Inpatient Care
Event|Activity|Discharge Instructions|15016,15020|false|false|false|C1947933|care activity|Care
Finding|Finding|Discharge Instructions|15016,15020|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Discharge Instructions|15016,15020|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Attribute|Clinical Attribute|Discharge Instructions|15016,15025|false|false|false|C4321316||Care Team
Finding|Finding|Discharge Instructions|15016,15025|false|false|false|C4321315|Care team|Care Team
Procedure|Health Care Activity|Discharge Instructions|15028,15036|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|15037,15049|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|15037,15049|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|15037,15049|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

