 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|49,58|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|49,58|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|49,63|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|83,92|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|83,92|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|83,92|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|83,92|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|83,92|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|83,97|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|115,120|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|115,120|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|115,120|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|139,142|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|139,142|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|139,142|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|139,142|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|139,142|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|150,157|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|150,157|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|SIMPLE_SEGMENT|159,166|false|false|false|||SURGERY
Finding|Finding|SIMPLE_SEGMENT|159,166|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Finding|Functional Concept|SIMPLE_SEGMENT|159,166|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Finding|Idea or Concept|SIMPLE_SEGMENT|159,166|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|159,166|false|false|false|C0543467|Operative Surgical Procedures|SURGERY
Attribute|Clinical Attribute|SIMPLE_SEGMENT|169,178|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|169,178|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|169,178|false|false|false|C0020517|Hypersensitivity|Allergies
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|184,187|false|false|false|C0013343|Dyes|Dye
Event|Event|SIMPLE_SEGMENT|184,187|false|false|false|||Dye
Drug|Biologically Active Substance|SIMPLE_SEGMENT|189,195|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|189,195|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|189,195|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Event|Activity|SIMPLE_SEGMENT|196,206|false|false|false|C2700400|Contain (action)|Containing
Event|Event|SIMPLE_SEGMENT|196,206|false|false|false|||Containing
Finding|Functional Concept|SIMPLE_SEGMENT|196,206|false|false|false|C0332256|Containing (qualifier value)|Containing
Event|Event|SIMPLE_SEGMENT|209,218|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|209,218|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|227,242|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|233,242|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|233,242|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|233,242|false|false|false|C5441521|Complaint (finding)|Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|244,250|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|244,250|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|244,250|false|false|false|C0027497|Nausea|nausea
Event|Event|SIMPLE_SEGMENT|252,260|false|false|false|||vomiting
Finding|Sign or Symptom|SIMPLE_SEGMENT|252,260|false|false|false|C0042963|Vomiting|vomiting
Finding|Idea or Concept|SIMPLE_SEGMENT|265,268|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|265,268|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Classification|SIMPLE_SEGMENT|271,276|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|277,285|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|277,285|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|289,307|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|298,307|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|298,307|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|298,307|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|298,307|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|298,307|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|SIMPLE_SEGMENT|316,323|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|316,323|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|316,323|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|316,323|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|316,326|false|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|316,342|false|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|316,342|false|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|327,334|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|327,334|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|327,342|false|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|335,342|false|false|false|C0221423|Illness (finding)|Illness
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|352,359|false|false|false|C0227391|Sigmoid colon|sigmoid
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|352,369|false|false|false|C0192866|Sigmoid colectomy|sigmoid colectomy
Event|Event|SIMPLE_SEGMENT|360,369|false|false|false|||colectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|360,369|false|false|false|C0009274|Colectomy|colectomy
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|384,398|false|false|false|C0012813|Diverticulitis|diverticulitis
Event|Event|SIMPLE_SEGMENT|384,398|false|false|false|||diverticulitis
Event|Event|SIMPLE_SEGMENT|407,417|false|false|false|||discharged
Event|Event|SIMPLE_SEGMENT|418,422|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|418,422|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|418,422|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|418,422|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|436,446|false|false|false|||tolerating
Finding|Finding|SIMPLE_SEGMENT|449,452|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|SIMPLE_SEGMENT|449,452|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|449,465|false|false|false|C0425404|Low residue diet|low residue diet
Finding|Conceptual Entity|SIMPLE_SEGMENT|453,460|false|false|false|C1709915|Residue|residue
Drug|Food|SIMPLE_SEGMENT|461,465|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|SIMPLE_SEGMENT|461,465|false|false|false|||diet
Finding|Functional Concept|SIMPLE_SEGMENT|461,465|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|SIMPLE_SEGMENT|461,465|false|false|false|C0012159|Diet therapy|diet
Drug|Antibiotic|SIMPLE_SEGMENT|474,485|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|SIMPLE_SEGMENT|474,485|false|false|false|||antibiotics
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|492,497|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Event|Event|SIMPLE_SEGMENT|492,497|false|false|false|||wound
Finding|Body Substance|SIMPLE_SEGMENT|492,497|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|SIMPLE_SEGMENT|492,497|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|SIMPLE_SEGMENT|492,497|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Pathologic Function|SIMPLE_SEGMENT|492,507|false|false|false|C0043241|Wound Infection|wound infection
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|498,507|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|498,507|false|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|498,507|false|false|false|C3714514|Infection|infection
Event|Event|SIMPLE_SEGMENT|514,522|false|false|false|||returned
Finding|Intellectual Product|SIMPLE_SEGMENT|527,531|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|SIMPLE_SEGMENT|539,548|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|539,548|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|539,548|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|539,548|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|539,548|false|false|false|C0030685|Patient Discharge|discharge
Finding|Idea or Concept|SIMPLE_SEGMENT|556,559|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|556,559|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Attribute|Clinical Attribute|SIMPLE_SEGMENT|571,577|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|571,577|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|571,577|false|false|false|C0027497|Nausea|nausea
Event|Event|SIMPLE_SEGMENT|582,588|false|false|false|||emesis
Finding|Body Substance|SIMPLE_SEGMENT|582,588|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Physiologic Function|SIMPLE_SEGMENT|582,588|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Sign or Symptom|SIMPLE_SEGMENT|582,588|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|622,628|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|622,628|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|622,628|false|false|false|C0027497|Nausea|nausea
Event|Event|SIMPLE_SEGMENT|632,642|false|false|false|||associated
Finding|Finding|SIMPLE_SEGMENT|651,657|false|false|false|C5202796|Intensity and Distress 1|slight
Event|Event|SIMPLE_SEGMENT|658,666|false|false|false|||increase
Finding|Functional Concept|SIMPLE_SEGMENT|658,666|false|false|false|C0442805|Increase|increase
Anatomy|Body Location or Region|SIMPLE_SEGMENT|670,680|false|false|false|C0521440|Epigastric|epigastric
Finding|Sign or Symptom|SIMPLE_SEGMENT|670,695|false|false|false|C0232493|Epigastric pain|epigastric abdominal pain
Anatomy|Body Location or Region|SIMPLE_SEGMENT|681,690|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|SIMPLE_SEGMENT|681,695|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|691,695|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|691,695|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|691,695|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|691,695|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Idea or Concept|SIMPLE_SEGMENT|709,720|false|false|false|C0750502|Significant|significant
Event|Event|SIMPLE_SEGMENT|721,731|false|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|721,731|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|721,731|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Event|SIMPLE_SEGMENT|735,739|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|735,739|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|735,739|false|false|false|C0582103|Medical Examination|exam
Finding|Finding|SIMPLE_SEGMENT|744,764|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|749,756|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|749,756|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|749,756|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|749,756|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|749,756|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|749,764|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|757,764|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|757,764|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|757,764|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|766,780|false|false|false|C0012813|Diverticulitis|diverticulitis
Event|Event|SIMPLE_SEGMENT|766,780|false|false|false|||diverticulitis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|785,788|false|false|false|C0396060|Congenital laryngeal adductor palsy|lap
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|785,788|false|false|false|C1870042|ACP2 protein, human|lap
Drug|Enzyme|SIMPLE_SEGMENT|785,788|false|false|false|C1870042|ACP2 protein, human|lap
Event|Event|SIMPLE_SEGMENT|785,788|false|false|false|||lap
Finding|Finding|SIMPLE_SEGMENT|785,788|false|false|false|C0456170;C1412132;C1413323;C1423544;C1424863;C1425522;C2827449;C3540509;C5575443;C5890955|ACP2 gene;ACP2 wt Allele;CEBPB gene;CEBPB wt Allele;CENPJ gene;LAP3 gene;LAP3 wt Allele;Left atrial pressure;PICALM gene;PICALM wt Allele|lap
Finding|Gene or Genome|SIMPLE_SEGMENT|785,788|false|false|false|C0456170;C1412132;C1413323;C1423544;C1424863;C1425522;C2827449;C3540509;C5575443;C5890955|ACP2 gene;ACP2 wt Allele;CEBPB gene;CEBPB wt Allele;CENPJ gene;LAP3 gene;LAP3 wt Allele;Left atrial pressure;PICALM gene;PICALM wt Allele|lap
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|785,788|false|false|false|C0031150|Laparoscopy|lap
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|789,796|false|false|false|C0227391|Sigmoid colon|sigmoid
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|789,806|false|false|false|C0192866|Sigmoid colectomy|sigmoid colectomy
Event|Event|SIMPLE_SEGMENT|797,806|false|false|false|||colectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|797,806|false|false|false|C0009274|Colectomy|colectomy
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|811,816|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Finding|Body Substance|SIMPLE_SEGMENT|811,816|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|SIMPLE_SEGMENT|811,816|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|SIMPLE_SEGMENT|811,816|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Pathologic Function|SIMPLE_SEGMENT|811,826|false|false|false|C0043241|Wound Infection|wound infection
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|817,826|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|817,826|false|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|817,826|false|false|false|C3714514|Infection|infection
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|828,837|false|false|false|C0149931|Migraine Disorders|Migraines
Event|Event|SIMPLE_SEGMENT|828,837|false|false|false|||Migraines
Finding|Functional Concept|SIMPLE_SEGMENT|838,842|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|843,849|false|false|false|C0016129;C0851278;C4299059|Fingers;Fingers not including thumb;Upper extremity>Finger|finger
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|850,860|false|false|false|C0007642|Cellulitis|cellulitis
Event|Event|SIMPLE_SEGMENT|850,860|false|false|false|||cellulitis
Finding|Finding|SIMPLE_SEGMENT|850,860|false|false|false|C2025995|cellulitis on exam (physical finding)|cellulitis
Finding|Functional Concept|SIMPLE_SEGMENT|863,869|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|863,877|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|870,877|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|870,877|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|870,877|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|870,877|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|883,889|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|883,889|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|883,889|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|883,889|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|883,897|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|890,897|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|890,897|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|890,897|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|890,897|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Event|Event|SIMPLE_SEGMENT|899,905|false|false|false|||father
Finding|Conceptual Entity|SIMPLE_SEGMENT|899,905|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Finding|Idea or Concept|SIMPLE_SEGMENT|899,905|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|915,922|false|true|false|C0009319|Colitis|colitis
Event|Event|SIMPLE_SEGMENT|915,922|false|false|false|||colitis
Event|Event|SIMPLE_SEGMENT|925,933|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|925,933|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|925,933|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|925,933|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|925,938|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|925,938|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|934,938|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|934,938|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|934,938|false|false|false|C0582103|Medical Examination|Exam
Event|Event|SIMPLE_SEGMENT|940,948|false|false|false|||afebrile
Finding|Finding|SIMPLE_SEGMENT|940,948|false|false|false|C0277797|Apyrexial|afebrile
Drug|Food|SIMPLE_SEGMENT|950,955|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|vital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|950,961|false|false|false|C0488614;C0518766|Vital signs|vital signs
Procedure|Health Care Activity|SIMPLE_SEGMENT|950,961|false|false|false|C0150404|Taking vital signs|vital signs
Event|Event|SIMPLE_SEGMENT|956,961|false|false|false|||signs
Finding|Finding|SIMPLE_SEGMENT|956,961|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|956,961|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Finding|SIMPLE_SEGMENT|962,982|false|false|false|C0442816||within normal limits
Event|Event|SIMPLE_SEGMENT|976,982|false|false|false|||limits
Finding|Functional Concept|SIMPLE_SEGMENT|976,982|false|false|false|C0439801|Limited (extensiveness)|limits
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|983,986|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|983,986|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|983,986|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|983,986|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|983,986|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|983,986|false|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|983,986|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Event|Event|SIMPLE_SEGMENT|988,997|false|false|false|||talkative
Finding|Individual Behavior|SIMPLE_SEGMENT|988,997|false|false|false|C0241331|talkative|talkative
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|998,1001|false|false|false|C0028863|Muscle of orbit|EOM
Finding|Functional Concept|SIMPLE_SEGMENT|998,1001|false|false|false|C0241886|Extraocular|EOM
Event|Event|SIMPLE_SEGMENT|1002,1006|false|false|false|||full
Event|Event|SIMPLE_SEGMENT|1008,1013|false|false|false|||PERRL
Finding|Finding|SIMPLE_SEGMENT|1008,1013|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Finding|Finding|SIMPLE_SEGMENT|1015,1024|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1025,1031|false|false|false|C0036410|Sclera|sclera
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1025,1031|false|false|false|C0036412|Scleral Diseases|sclera
Event|Event|SIMPLE_SEGMENT|1025,1031|false|false|false|||sclera
Procedure|Health Care Activity|SIMPLE_SEGMENT|1025,1031|false|false|false|C2228481|examination of sclera|sclera
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1032,1037|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|SIMPLE_SEGMENT|1032,1037|false|false|false|C0741025|Chest problem|Chest
Finding|Finding|SIMPLE_SEGMENT|1032,1043|false|false|false|C0578395|chest clear|Chest clear
Event|Event|SIMPLE_SEGMENT|1038,1043|false|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|1038,1043|false|false|false|C1550016|Remote control command - Clear|clear
Event|Event|SIMPLE_SEGMENT|1044,1047|false|false|false|||RRR
Event|Event|SIMPLE_SEGMENT|1052,1059|false|false|false|||murmurs
Finding|Finding|SIMPLE_SEGMENT|1052,1059|true|false|false|C0018808|Heart murmur|murmurs
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1060,1067|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1060,1067|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Finding|Finding|SIMPLE_SEGMENT|1060,1067|false|false|false|C0941288|Abdomen problem|Abdomen
Finding|Finding|SIMPLE_SEGMENT|1060,1072|false|false|false|C0426663|Abdomen soft|Abdomen soft
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1068,1072|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|SIMPLE_SEGMENT|1068,1072|false|false|false|||soft
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1125,1144|false|false|false|C1261209|Transverse incision|transverse incision
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1136,1144|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|1136,1144|false|false|false|C0332803|Surgical wound|incision
Event|Event|SIMPLE_SEGMENT|1136,1144|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1136,1144|false|false|false|C0184898|Surgical incisions|incision
Anatomy|Tissue|SIMPLE_SEGMENT|1157,1165|false|false|false|C0222331;C0278403|Subcutaneous Fat;Subcutaneous Tissue|subcutis
Finding|Finding|SIMPLE_SEGMENT|1171,1177|false|false|false|C1554187|Gender Status - Intact|intact
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1178,1182|false|false|false|C4318566|Deep Resection Margin|deep
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1184,1190|false|false|false|C0015641|Fascia|fascia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1195,1203|true|false|false|C0041834|Erythema|erythema
Event|Event|SIMPLE_SEGMENT|1195,1203|false|false|false|||erythema
Event|Event|SIMPLE_SEGMENT|1207,1217|false|false|false|||induration
Finding|Pathologic Function|SIMPLE_SEGMENT|1207,1217|true|false|false|C0332534|Induration|induration
Event|Event|SIMPLE_SEGMENT|1234,1240|false|false|false|||output
Finding|Conceptual Entity|SIMPLE_SEGMENT|1234,1240|false|false|false|C1709366|system output|output
Procedure|Health Care Activity|SIMPLE_SEGMENT|1234,1240|false|false|false|C3251815|Measurement of fluid output|output
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1256,1261|true|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|1256,1261|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|1256,1261|true|false|false|C0013604|Edema|edema
Drug|Food|SIMPLE_SEGMENT|1269,1275|false|false|false|C5890763||pulses
Event|Event|SIMPLE_SEGMENT|1269,1275|false|false|false|||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|1269,1275|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|1269,1275|false|false|false|C0034107|Pulse taking|pulses
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1297,1307|false|false|false|C1644645||CT ABDOMEN
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1297,1307|false|false|false|C0412620|CT of abdomen|CT ABDOMEN
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1297,1320|false|false|false|C0202838|Computed tomography, abdomen; without contrast material|CT ABDOMEN W/O CONTRAST
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1300,1307|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1300,1307|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|SIMPLE_SEGMENT|1300,1307|false|false|false|||ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|1300,1307|false|false|false|C0941288|Abdomen problem|ABDOMEN
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|1312,1320|false|false|false|C0009924|Contrast Media|CONTRAST
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|1342,1350|false|true|false|C0009924|Contrast Media|CONTRAST
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1352,1361|false|false|false|C0882057||CT PELVIS
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1352,1361|false|false|false|C0412628|Computed tomography of pelvis|CT PELVIS
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1355,1361|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|PELVIS
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|1355,1361|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|PELVIS
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1355,1361|false|false|false|C0153663|Malignant neoplasm of pelvis|PELVIS
Event|Event|SIMPLE_SEGMENT|1355,1361|false|false|false|||PELVIS
Finding|Finding|SIMPLE_SEGMENT|1355,1361|false|false|false|C0812455|Pelvis problem|PELVIS
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|1366,1374|false|false|false|C0009924|Contrast Media|CONTRAST
Event|Event|SIMPLE_SEGMENT|1376,1382|false|false|false|||Reason
Finding|Idea or Concept|SIMPLE_SEGMENT|1376,1382|false|false|false|C0392360|Indication of (contextual qualifier)|Reason
Event|Event|SIMPLE_SEGMENT|1384,1385|false|false|false|||r
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1388,1395|false|true|false|C0000833|Abscess|abscess
Event|Event|SIMPLE_SEGMENT|1388,1395|false|false|false|||abscess
Finding|Intellectual Product|SIMPLE_SEGMENT|1388,1395|false|true|false|C1546533||abscess
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|1399,1410|true|false|false|C4072741|IV contrast|IV contrast
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|1402,1410|true|false|false|C0009924|Contrast Media|contrast
Event|Event|SIMPLE_SEGMENT|1402,1410|false|false|false|||contrast
Event|Event|SIMPLE_SEGMENT|1421,1426|false|false|false|||Field
Finding|Conceptual Entity|SIMPLE_SEGMENT|1421,1426|false|false|false|C1521738;C2346620;C2349184|Field;Force Field;Knowledge Field|Field
Procedure|Health Care Activity|SIMPLE_SEGMENT|1421,1426|false|false|false|C1553496|field - patient encounter|Field
Event|Event|SIMPLE_SEGMENT|1451,1458|false|false|false|||MEDICAL
Finding|Functional Concept|SIMPLE_SEGMENT|1451,1458|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|MEDICAL
Finding|Idea or Concept|SIMPLE_SEGMENT|1451,1458|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|MEDICAL
Finding|Intellectual Product|SIMPLE_SEGMENT|1451,1458|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|MEDICAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|1451,1458|false|false|false|C0199168|Medical service|MEDICAL
Finding|Finding|SIMPLE_SEGMENT|1451,1468|false|false|false|C4745084|Medical Condition|MEDICAL CONDITION
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1459,1468|false|false|false|C3864998||CONDITION
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1459,1468|false|false|false|C0012634|Disease|CONDITION
Event|Event|SIMPLE_SEGMENT|1459,1468|false|false|false|||CONDITION
Finding|Conceptual Entity|SIMPLE_SEGMENT|1459,1468|false|false|false|C1705253|Logical Condition|CONDITION
Finding|Idea or Concept|SIMPLE_SEGMENT|1474,1478|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|SIMPLE_SEGMENT|1474,1478|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|SIMPLE_SEGMENT|1479,1482|false|false|false|||old
Event|Event|SIMPLE_SEGMENT|1483,1488|false|false|false|||woman
Event|Event|SIMPLE_SEGMENT|1511,1520|false|false|false|||colectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1511,1520|false|false|false|C0009274|Colectomy|colectomy
Anatomy|Cell|SIMPLE_SEGMENT|1541,1544|false|false|false|C0023516|Leukocytes|WBC
Event|Event|SIMPLE_SEGMENT|1541,1544|false|false|false|||WBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1549,1555|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|1549,1555|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1549,1555|false|false|false|C0027497|Nausea|nausea
Event|Event|SIMPLE_SEGMENT|1557,1563|false|false|false|||REASON
Finding|Idea or Concept|SIMPLE_SEGMENT|1557,1563|false|false|false|C0392360|Indication of (contextual qualifier)|REASON
Finding|Idea or Concept|SIMPLE_SEGMENT|1557,1567|false|false|false|C0392360|Indication of (contextual qualifier)|REASON FOR
Event|Activity|SIMPLE_SEGMENT|1573,1584|false|false|false|C4321457|Examination|EXAMINATION
Event|Event|SIMPLE_SEGMENT|1573,1584|false|false|false|||EXAMINATION
Procedure|Health Care Activity|SIMPLE_SEGMENT|1573,1584|false|false|false|C0031809;C0582103|Medical Examination;Physical Examination|EXAMINATION
Event|Event|SIMPLE_SEGMENT|1586,1587|false|false|false|||r
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1590,1597|false|true|false|C0000833|Abscess|abscess
Event|Event|SIMPLE_SEGMENT|1590,1597|false|false|false|||abscess
Finding|Intellectual Product|SIMPLE_SEGMENT|1590,1597|false|true|false|C1546533||abscess
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|1601,1612|true|false|false|C4072741|IV contrast|IV contrast
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|1604,1612|true|false|false|C0009924|Contrast Media|contrast
Event|Event|SIMPLE_SEGMENT|1604,1612|false|false|false|||contrast
Event|Event|SIMPLE_SEGMENT|1623,1640|false|false|false|||CONTRAINDICATIONS
Finding|Finding|SIMPLE_SEGMENT|1623,1640|false|false|false|C1301624|Medical contraindication|CONTRAINDICATIONS
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|1645,1656|false|false|false|C4072741|IV contrast|IV CONTRAST
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|1648,1656|false|false|false|C0009924|Contrast Media|CONTRAST
Event|Event|SIMPLE_SEGMENT|1648,1656|false|false|false|||CONTRAST
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1662,1672|false|false|false|C5890010||INDICATION
Event|Event|SIMPLE_SEGMENT|1662,1672|false|false|false|||INDICATION
Finding|Idea or Concept|SIMPLE_SEGMENT|1662,1672|false|false|false|C0392360;C3146298|Indication;Indication of (contextual qualifier)|INDICATION
Anatomy|Cell|SIMPLE_SEGMENT|1698,1714|false|false|false|C0023516|Leukocytes|white blood cell
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1704,1709|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|1704,1709|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|1704,1709|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Anatomy|Cell|SIMPLE_SEGMENT|1704,1714|false|false|false|C0005773|Blood Cells|blood cell
Anatomy|Cell|SIMPLE_SEGMENT|1710,1714|false|false|false|C0007634|Cells|cell
Finding|Gene or Genome|SIMPLE_SEGMENT|1710,1714|false|false|false|C1413336;C1413337|CEL gene;CELP gene|cell
Event|Event|SIMPLE_SEGMENT|1716,1721|false|false|false|||count
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1726,1732|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|1726,1732|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1726,1732|false|false|false|C0027497|Nausea|nausea
Event|Event|SIMPLE_SEGMENT|1734,1741|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|1734,1741|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|1734,1741|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|1734,1741|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|1734,1744|false|false|false|C0262926|Medical History|history of
Event|Event|SIMPLE_SEGMENT|1752,1761|false|false|false|||colectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1752,1761|false|false|false|C0009274|Colectomy|colectomy
Event|Event|SIMPLE_SEGMENT|1766,1775|false|false|false|||recurrent
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1777,1791|false|false|false|C0012813|Diverticulitis|diverticulitis
Event|Event|SIMPLE_SEGMENT|1777,1791|false|false|false|||diverticulitis
Event|Activity|SIMPLE_SEGMENT|1794,1804|false|false|false|C1707455|Comparison|COMPARISON
Event|Event|SIMPLE_SEGMENT|1794,1804|false|false|false|||COMPARISON
Event|Event|SIMPLE_SEGMENT|1806,1808|false|false|false|||CT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1806,1816|false|false|false|C1644645||CT abdomen
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1806,1816|false|false|false|C0412620|CT of abdomen|CT abdomen
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1806,1827|false|false|false|C1715387||CT abdomen and pelvis
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1809,1816|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1809,1816|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Event|Event|SIMPLE_SEGMENT|1809,1816|false|false|false|||abdomen
Finding|Finding|SIMPLE_SEGMENT|1809,1816|false|false|false|C0941288|Abdomen problem|abdomen
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1809,1820|false|false|false|C0000726|Abdomen|abdomen and
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1809,1827|false|false|false|C1508499|Abdominopelvic structure|abdomen and pelvis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1821,1827|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|1821,1827|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1821,1827|false|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Event|Event|SIMPLE_SEGMENT|1821,1827|false|false|false|||pelvis
Finding|Finding|SIMPLE_SEGMENT|1821,1827|false|false|false|C0812455|Pelvis problem|pelvis
Finding|Functional Concept|SIMPLE_SEGMENT|1837,1846|false|false|false|C0449851|Techniques|TECHNIQUE
Event|Event|SIMPLE_SEGMENT|1848,1852|false|false|false|||MDCT
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1848,1852|false|false|false|C3179130|Multidetector Computed Tomography|MDCT
Finding|Intellectual Product|SIMPLE_SEGMENT|1853,1861|false|false|false|C3245488|Acquired Name|acquired
Event|Event|SIMPLE_SEGMENT|1868,1874|false|false|false|||images
Event|Event|SIMPLE_SEGMENT|1880,1888|false|false|false|||obtained
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1902,1909|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1902,1909|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Event|Event|SIMPLE_SEGMENT|1902,1909|false|false|false|||abdomen
Finding|Finding|SIMPLE_SEGMENT|1902,1909|false|false|false|C0941288|Abdomen problem|abdomen
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1902,1913|false|false|false|C0000726|Abdomen|abdomen and
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1902,1920|false|false|false|C1508499|Abdominopelvic structure|abdomen and pelvis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1914,1920|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|1914,1920|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1914,1920|false|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Event|Event|SIMPLE_SEGMENT|1914,1920|false|false|false|||pelvis
Finding|Finding|SIMPLE_SEGMENT|1914,1920|false|false|false|C0812455|Pelvis problem|pelvis
Event|Event|SIMPLE_SEGMENT|1931,1945|false|false|false|||administration
Event|Occupational Activity|SIMPLE_SEGMENT|1931,1945|false|false|false|C0001554|Administration occupational activities|administration
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1931,1945|false|false|false|C1533734|Administration (procedure)|administration
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|1949,1953|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1949,1953|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|1949,1953|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|1949,1953|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|1954,1962|false|false|false|C0009924|Contrast Media|contrast
Event|Event|SIMPLE_SEGMENT|1954,1962|false|false|false|||contrast
Finding|Functional Concept|SIMPLE_SEGMENT|1968,1979|false|false|false|C1522726|Intravenous Route of Administration|intravenous
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|1968,1988|false|false|false|C4072741|IV contrast|intravenous contrast
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|1980,1988|false|false|false|C0009924|Contrast Media|contrast
Event|Event|SIMPLE_SEGMENT|1980,1988|false|false|false|||contrast
Event|Event|SIMPLE_SEGMENT|1993,2005|false|false|false|||administered
Event|Event|SIMPLE_SEGMENT|2019,2030|false|false|false|||reformatted
Event|Event|SIMPLE_SEGMENT|2032,2038|false|false|false|||images
Event|Event|SIMPLE_SEGMENT|2049,2057|false|false|false|||obtained
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2060,2068|false|false|false|C2926606||FINDINGS
Event|Event|SIMPLE_SEGMENT|2060,2068|false|false|false|||FINDINGS
Finding|Functional Concept|SIMPLE_SEGMENT|2060,2068|false|false|false|C2607943|findings aspects|FINDINGS
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2076,2080|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2076,2080|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2076,2080|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|2076,2080|false|false|false|C0740941|Lung Problem|lung
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|2081,2086|false|false|false|C0178499|Base|bases
Event|Event|SIMPLE_SEGMENT|2081,2086|false|false|false|||bases
Event|Event|SIMPLE_SEGMENT|2091,2096|false|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|2091,2096|false|false|false|C1550016|Remote control command - Clear|clear
Finding|Pathologic Function|SIMPLE_SEGMENT|2105,2124|false|false|false|C0333404|Calcified granuloma|calcified granuloma
Event|Event|SIMPLE_SEGMENT|2115,2124|false|false|false|||granuloma
Finding|Intellectual Product|SIMPLE_SEGMENT|2115,2124|false|false|false|C0018188;C1546654|Granuloma|granuloma
Finding|Pathologic Function|SIMPLE_SEGMENT|2115,2124|false|false|false|C0018188;C1546654|Granuloma|granuloma
Finding|Functional Concept|SIMPLE_SEGMENT|2133,2138|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2133,2143|false|false|false|C0225706|Right lung|right lung
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2133,2148|false|false|false|C0225708|Structure of base of right lung|right lung base
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2139,2143|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2139,2143|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2139,2143|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|2139,2143|false|false|false|C0740941|Lung Problem|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2139,2148|false|false|false|C0225704|Basal segment of lung|lung base
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2144,2148|false|false|false|C2987514|Anatomical base|base
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2144,2148|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|2144,2148|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|2144,2148|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Event|Event|SIMPLE_SEGMENT|2144,2148|false|false|false|||base
Finding|Gene or Genome|SIMPLE_SEGMENT|2144,2148|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Finding|Idea or Concept|SIMPLE_SEGMENT|2144,2148|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Event|Event|SIMPLE_SEGMENT|2152,2161|false|false|false|||unchanged
Finding|Finding|SIMPLE_SEGMENT|2152,2161|false|false|false|C0442739||unchanged
Finding|Functional Concept|SIMPLE_SEGMENT|2163,2170|false|false|false|C0439801;C3542948|Limited (extensiveness);Limited component (foundation metadata concept)|Limited
Finding|Intellectual Product|SIMPLE_SEGMENT|2163,2170|false|false|false|C0439801;C3542948|Limited (extensiveness);Limited component (foundation metadata concept)|Limited
Event|Event|SIMPLE_SEGMENT|2171,2177|false|false|false|||images
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2185,2190|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2185,2190|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|2185,2190|false|false|false|C0795691|HEART PROBLEM|heart
Event|Event|SIMPLE_SEGMENT|2196,2208|false|false|false|||unremarkable
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2222,2233|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2222,2233|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2222,2242|true|false|false|C0031039|Pericardial effusion|pericardial effusion
Finding|Body Substance|SIMPLE_SEGMENT|2222,2242|true|false|false|C1253937|Pericardial effusion body substance|pericardial effusion
Event|Event|SIMPLE_SEGMENT|2234,2242|false|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|2234,2242|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|2234,2242|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|2234,2242|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2252,2259|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2252,2259|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Finding|Finding|SIMPLE_SEGMENT|2252,2259|false|false|false|C0941288|Abdomen problem|abdomen
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2265,2270|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2265,2270|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2265,2270|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|SIMPLE_SEGMENT|2265,2270|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2265,2270|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|SIMPLE_SEGMENT|2265,2270|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|SIMPLE_SEGMENT|2265,2270|false|false|false|||liver
Finding|Finding|SIMPLE_SEGMENT|2265,2270|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|SIMPLE_SEGMENT|2265,2270|false|false|false|C0872387|Procedures on liver|liver
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2272,2283|false|false|false|C0016976;C1524055;C4071903|Abdomen>Gallbladder;Gallbladder;Gallbladder (MMHCC)|gallbladder
Anatomy|Tissue|SIMPLE_SEGMENT|2272,2283|false|false|false|C0016976;C1524055;C4071903|Abdomen>Gallbladder;Gallbladder;Gallbladder (MMHCC)|gallbladder
Event|Event|SIMPLE_SEGMENT|2272,2283|false|false|false|||gallbladder
Procedure|Health Care Activity|SIMPLE_SEGMENT|2272,2283|false|false|false|C2032932|examination of gallbladder|gallbladder
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2285,2291|false|false|false|C0037993;C4037984|Abdomen>Spleen;Spleen|spleen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2285,2291|false|false|false|C0153470|Malignant neoplasm of spleen|spleen
Event|Event|SIMPLE_SEGMENT|2285,2291|false|false|false|||spleen
Finding|Finding|SIMPLE_SEGMENT|2285,2291|false|false|false|C0812414|Spleen problem|spleen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2285,2291|false|false|false|C0869677|Procedures on Spleen|spleen
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2293,2300|false|false|false|C0022646;C0227665|Both kidneys;Kidney|kidneys
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2302,2309|false|false|false|C0001625|Adrenal Glands|adrenal
Finding|Finding|SIMPLE_SEGMENT|2302,2309|false|false|false|C0521428|Adrenal|adrenal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2311,2317|false|false|false|C1285092|Gland|glands
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2319,2327|false|false|false|C0030274;C4037927|Abdomen>Pancreas;Pancreas|pancreas
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2319,2327|false|false|false|C0030286;C0347284|Benign tumor of pancreas;Pancreatic Diseases|pancreas
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2319,2327|false|false|false|C0030286;C0347284|Benign tumor of pancreas;Pancreatic Diseases|pancreas
Drug|Organic Chemical|SIMPLE_SEGMENT|2319,2327|false|false|false|C0771711|pancreas extract|pancreas
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2319,2327|false|false|false|C0771711|pancreas extract|pancreas
Event|Event|SIMPLE_SEGMENT|2319,2327|false|false|false|||pancreas
Finding|Finding|SIMPLE_SEGMENT|2319,2327|false|false|false|C0813176|Pancreas problem|pancreas
Procedure|Health Care Activity|SIMPLE_SEGMENT|2319,2327|false|false|false|C0869826|Procedures on Pancreas|pancreas
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2329,2336|false|false|false|C0038351;C3714551;C4266636|Abdomen>Stomach;Stomach;Stomach structure|stomach
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2329,2336|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2329,2336|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Event|Event|SIMPLE_SEGMENT|2329,2336|false|false|false|||stomach
Finding|Finding|SIMPLE_SEGMENT|2329,2336|false|false|false|C0577027|Stomach problem|stomach
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2329,2336|false|false|false|C0872393|Procedure on stomach|stomach
Finding|Functional Concept|SIMPLE_SEGMENT|2342,2357|false|false|false|C1512911|Intraabdominal Route of Administration|intra-abdominal
Event|Event|SIMPLE_SEGMENT|2358,2363|false|false|false|||loops
Finding|Gene or Genome|SIMPLE_SEGMENT|2378,2383|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2378,2389|false|false|false|C0021851|Large Intestine|large bowel
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2384,2389|false|false|false|C0021853|Intestines|bowel
Event|Event|SIMPLE_SEGMENT|2394,2406|false|false|false|||unremarkable
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2420,2430|false|false|false|C0025474|Mesentery|mesenteric
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2432,2447|false|false|false|C0497156|Lymphadenopathy|lymphadenopathy
Event|Event|SIMPLE_SEGMENT|2432,2447|false|false|false|||lymphadenopathy
Finding|Sign or Symptom|SIMPLE_SEGMENT|2432,2447|false|false|false|C4282165|Swollen Lymph Node|lymphadenopathy
Finding|Functional Concept|SIMPLE_SEGMENT|2461,2465|true|false|false|C0332296|Free of (attribute)|free
Finding|Pathologic Function|SIMPLE_SEGMENT|2461,2471|true|false|false|C0013687|effusion|free fluid
Drug|Substance|SIMPLE_SEGMENT|2466,2471|true|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|2466,2471|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|2466,2471|true|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|2475,2479|false|false|false|||free
Finding|Functional Concept|SIMPLE_SEGMENT|2475,2479|true|false|false|C0332296|Free of (attribute)|free
Drug|Inorganic Chemical|SIMPLE_SEGMENT|2480,2483|true|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2480,2483|true|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|SIMPLE_SEGMENT|2480,2483|true|false|false|C0001861;C3536832|Air (substance);air|air
Event|Event|SIMPLE_SEGMENT|2480,2483|false|false|false|||air
Finding|Finding|SIMPLE_SEGMENT|2480,2483|true|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|SIMPLE_SEGMENT|2480,2483|true|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|SIMPLE_SEGMENT|2480,2483|true|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2492,2499|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2492,2499|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Event|Event|SIMPLE_SEGMENT|2492,2499|false|false|false|||abdomen
Finding|Finding|SIMPLE_SEGMENT|2492,2499|false|false|false|C0941288|Abdomen problem|abdomen
Event|Event|SIMPLE_SEGMENT|2513,2521|false|false|false|||adjacent
Finding|Functional Concept|SIMPLE_SEGMENT|2529,2533|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2529,2553|false|false|false|C0226363|Structure of left common iliac artery|left common iliac artery
Finding|Functional Concept|SIMPLE_SEGMENT|2534,2540|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Finding|Intellectual Product|SIMPLE_SEGMENT|2534,2540|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2534,2553|false|false|false|C1261084|Common iliac artery structure|common iliac artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2541,2546|false|false|false|C0020889|Bone structure of ilium|iliac
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2541,2553|false|false|false|C0020887|Structure of iliac artery|iliac artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2547,2553|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|2547,2553|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Event|Event|SIMPLE_SEGMENT|2568,2573|false|false|false|||focus
Finding|Functional Concept|SIMPLE_SEGMENT|2568,2573|false|false|false|C1285542|Has focus|focus
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2577,2582|false|false|false|C0424295|Hyperactive behavior|hyper
Drug|Substance|SIMPLE_SEGMENT|2595,2603|false|false|false|C0520510|Materials|material
Event|Event|SIMPLE_SEGMENT|2595,2603|false|false|false|||material
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2615,2625|false|false|false|C0550215||appearance
Event|Event|SIMPLE_SEGMENT|2615,2625|false|false|false|||appearance
Procedure|Health Care Activity|SIMPLE_SEGMENT|2615,2625|false|false|false|C2051406|patient appearance regarding mental status exam|appearance
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|2629,2635|false|false|false|C0502420|Suture Joint|suture
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2629,2635|false|false|false|C1706068|Suture Dosage Form|suture
Finding|Intellectual Product|SIMPLE_SEGMENT|2629,2635|false|false|false|C1546803||suture
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2629,2635|false|false|false|C0009068|Closure by suture|suture
Drug|Substance|SIMPLE_SEGMENT|2636,2644|false|false|false|C0520510|Materials|material
Event|Event|SIMPLE_SEGMENT|2636,2644|false|false|false|||material
Event|Event|SIMPLE_SEGMENT|2654,2663|false|false|false|||unchanged
Finding|Finding|SIMPLE_SEGMENT|2654,2663|false|false|false|C0442739||unchanged
Event|Activity|SIMPLE_SEGMENT|2680,2691|false|false|false|C4321457|Examination|examination
Event|Event|SIMPLE_SEGMENT|2680,2691|false|false|false|||examination
Procedure|Health Care Activity|SIMPLE_SEGMENT|2680,2691|false|false|false|C0031809;C0582103|Medical Examination;Physical Examination|examination
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2701,2707|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|2701,2707|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2701,2707|true|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Finding|Finding|SIMPLE_SEGMENT|2701,2707|true|false|false|C0812455|Pelvis problem|pelvis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|2709,2715|false|false|false|C0502420|Suture Joint|suture
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2709,2715|false|false|false|C1706068|Suture Dosage Form|suture
Finding|Intellectual Product|SIMPLE_SEGMENT|2709,2715|false|false|false|C1546803||suture
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2709,2715|false|false|false|C0009068|Closure by suture|suture
Drug|Substance|SIMPLE_SEGMENT|2716,2724|false|false|false|C0520510|Materials|material
Event|Event|SIMPLE_SEGMENT|2716,2724|false|false|false|||material
Event|Event|SIMPLE_SEGMENT|2728,2732|false|false|false|||seen
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2740,2746|false|false|false|C4522154|Distal Resection Margin|distal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2747,2754|false|false|false|C0227391|Sigmoid colon|sigmoid
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2756,2761|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2756,2761|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2756,2761|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Event|Event|SIMPLE_SEGMENT|2756,2761|false|false|false|||colon
Finding|Finding|SIMPLE_SEGMENT|2756,2761|false|false|false|C0750873|COLON PROBLEM|colon
Event|Event|SIMPLE_SEGMENT|2763,2772|false|false|false|||unchanged
Finding|Finding|SIMPLE_SEGMENT|2763,2772|false|false|false|C0442739||unchanged
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2776,2786|false|false|false|C0550215||appearance
Event|Event|SIMPLE_SEGMENT|2776,2786|false|false|false|||appearance
Procedure|Health Care Activity|SIMPLE_SEGMENT|2776,2786|false|false|false|C2051406|patient appearance regarding mental status exam|appearance
Event|Activity|SIMPLE_SEGMENT|2798,2809|false|false|false|C4321457|Examination|examination
Event|Event|SIMPLE_SEGMENT|2798,2809|false|false|false|||examination
Procedure|Health Care Activity|SIMPLE_SEGMENT|2798,2809|false|false|false|C0031809;C0582103|Medical Examination;Physical Examination|examination
Event|Event|SIMPLE_SEGMENT|2815,2825|false|false|false|||consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|2815,2825|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|2815,2830|false|false|false|C0332290|Consistent with|consistent with
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2831,2838|false|false|false|C0009368|Colon structure (body structure)|colonic
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2831,2850|false|false|false|C0852681|Large intestine anastomosis|colonic anastomosis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|2839,2850|false|false|false|C0500470|Anatomical anastomosis|anastomosis
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|2839,2850|false|false|false|C0332853|Anastomosis|anastomosis
Event|Event|SIMPLE_SEGMENT|2839,2850|false|false|false|||anastomosis
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2839,2850|false|false|false|C0677554||anastomosis
Event|Event|SIMPLE_SEGMENT|2864,2872|false|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|2864,2872|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|2864,2875|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Event|Event|SIMPLE_SEGMENT|2877,2886|false|false|false|||stricture
Finding|Pathologic Function|SIMPLE_SEGMENT|2877,2886|false|false|false|C1261287|Stenosis|stricture
Event|Event|SIMPLE_SEGMENT|2890,2901|false|false|false|||obstruction
Finding|Finding|SIMPLE_SEGMENT|2890,2901|true|false|false|C0028778|Obstruction|obstruction
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2910,2914|false|false|false|C1515974|Anatomic Site|site
Finding|Intellectual Product|SIMPLE_SEGMENT|2910,2914|false|false|false|C1546778||site
Finding|Idea or Concept|SIMPLE_SEGMENT|2928,2933|true|false|false|C1550012|Local Remote Control State - Local|local
Drug|Substance|SIMPLE_SEGMENT|2934,2939|true|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|2934,2939|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|2934,2939|true|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|2941,2951|false|false|false|||collection
Finding|Conceptual Entity|SIMPLE_SEGMENT|2941,2951|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|2941,2951|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|2941,2951|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|2941,2951|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Event|Event|SIMPLE_SEGMENT|2955,2963|false|false|false|||indicate
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2964,2971|false|false|false|C0000833|Abscess|abscess
Event|Event|SIMPLE_SEGMENT|2964,2971|false|false|false|||abscess
Finding|Intellectual Product|SIMPLE_SEGMENT|2964,2971|false|false|false|C1546533||abscess
Event|Event|SIMPLE_SEGMENT|2986,2991|false|false|false|||signs
Finding|Finding|SIMPLE_SEGMENT|2986,2991|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|2986,2991|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Event|Event|SIMPLE_SEGMENT|2996,3008|false|false|false|||inflammation
Finding|Pathologic Function|SIMPLE_SEGMENT|2996,3008|false|false|false|C0021368|Inflammation|inflammation
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|3014,3025|false|false|false|C0559769|Pelvic cavity structure|intrapelvic
Event|Event|SIMPLE_SEGMENT|3026,3031|false|false|false|||loops
Finding|Gene or Genome|SIMPLE_SEGMENT|3045,3050|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3045,3056|false|false|false|C0021851|Large Intestine|large bowel
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3051,3056|false|false|false|C0021853|Intestines|bowel
Event|Event|SIMPLE_SEGMENT|3062,3074|false|false|false|||unremarkable
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3087,3090|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3087,3090|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|SIMPLE_SEGMENT|3087,3090|false|false|false|C0001861;C3536832|Air (substance);air|air
Event|Event|SIMPLE_SEGMENT|3087,3090|false|false|false|||air
Finding|Finding|SIMPLE_SEGMENT|3087,3090|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|SIMPLE_SEGMENT|3087,3090|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|SIMPLE_SEGMENT|3087,3090|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Event|Event|SIMPLE_SEGMENT|3095,3100|false|false|false|||stool
Finding|Body Substance|SIMPLE_SEGMENT|3095,3100|false|false|false|C0015733|Feces|stool
Event|Event|SIMPLE_SEGMENT|3113,3120|false|false|false|||pattern
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3130,3135|false|false|false|C0021853|Intestines|bowel
Event|Event|SIMPLE_SEGMENT|3136,3146|false|false|false|||dilatation
Finding|Finding|SIMPLE_SEGMENT|3136,3146|true|false|false|C0012359;C0700124|Dilated;Pathological Dilatation|dilatation
Finding|Pathologic Function|SIMPLE_SEGMENT|3136,3146|true|false|false|C0012359;C0700124|Dilated;Pathological Dilatation|dilatation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3136,3146|true|false|false|C1322279|Dilate procedure|dilatation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3152,3160|false|false|false|C0003617;C4037994|Abdomen+Pelvis>Appendix;Appendix|appendix
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3152,3160|false|false|false|C0348899;C0496779;C0496860|Benign neoplasm of appendix;Malignant neoplasm of appendix;Neoplasm of uncertain or unknown behavior of appendix|appendix
Event|Event|SIMPLE_SEGMENT|3152,3160|false|false|false|||appendix
Finding|Intellectual Product|SIMPLE_SEGMENT|3152,3160|false|false|false|C1552860|appendix - HTML link|appendix
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3152,3160|false|false|false|C0869813|Procedure on appendix|appendix
Event|Event|SIMPLE_SEGMENT|3164,3174|false|false|false|||visualized
Event|Event|SIMPLE_SEGMENT|3183,3189|false|false|false|||normal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3195,3202|false|false|false|C0042027|Urinary tract|urinary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3195,3210|false|false|false|C0005682;C4037992|Abdomen+Pelvis>Urinary bladder;Urinary Bladder|urinary bladder
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3203,3210|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3203,3210|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Event|Event|SIMPLE_SEGMENT|3203,3210|false|false|false|||bladder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3203,3210|false|false|false|C0872388|Procedures on bladder|bladder
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3212,3218|false|false|false|C0042149;C1519876;C4266525|Mouse Uterus;Pelvis>Uterus;Uterus|uterus
Anatomy|Tissue|SIMPLE_SEGMENT|3212,3218|false|false|false|C0042149;C1519876;C4266525|Mouse Uterus;Pelvis>Uterus;Uterus|uterus
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3212,3218|false|false|false|C0042131;C0496919|Neoplasm of uncertain or unknown behavior of uterus;Uterine Diseases|uterus
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3212,3218|false|false|false|C0042131;C0496919|Neoplasm of uncertain or unknown behavior of uterus;Uterine Diseases|uterus
Event|Event|SIMPLE_SEGMENT|3212,3218|false|false|false|||uterus
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3212,3218|false|false|false|C0869889|examination of uterus|uterus
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3224,3230|false|false|false|C0001575;C0229243;C4522151|Adnexa;Ocular adnexa structure;Uterine adnexae structure|adnexa
Event|Event|SIMPLE_SEGMENT|3236,3248|false|false|false|||unremarkable
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3274,3282|false|false|false|C1293134|Enlargement procedure|enlarged
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3274,3294|true|false|false|C0497156|Lymphadenopathy|enlarged lymph nodes
Finding|Sign or Symptom|SIMPLE_SEGMENT|3274,3294|true|false|false|C4282165|Swollen Lymph Node|enlarged lymph nodes
Finding|Body Substance|SIMPLE_SEGMENT|3283,3288|false|false|false|C0024202|Lymph|lymph
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3283,3294|false|false|false|C0024204|lymph nodes|lymph nodes
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3283,3294|true|false|false|C0154054|benign neoplasm of lymph nodes|lymph nodes
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3303,3309|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|3303,3309|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3303,3309|false|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Event|Event|SIMPLE_SEGMENT|3303,3309|false|false|false|||pelvis
Finding|Finding|SIMPLE_SEGMENT|3303,3309|false|false|false|C0812455|Pelvis problem|pelvis
Anatomy|Tissue|SIMPLE_SEGMENT|3313,3316|false|false|false|C0001527|Adipose tissue|fat
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3313,3316|false|false|false|C0015677;C1435181;C3887682|FAT1 protein, human;Fatty acid glycerol esters;Platelet Glycoprotein 4, human|fat
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3313,3316|false|false|false|C0015677;C1435181;C3887682|FAT1 protein, human;Fatty acid glycerol esters;Platelet Glycoprotein 4, human|fat
Drug|Organic Chemical|SIMPLE_SEGMENT|3313,3316|false|false|false|C0015677;C1435181;C3887682|FAT1 protein, human;Fatty acid glycerol esters;Platelet Glycoprotein 4, human|fat
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3313,3316|false|false|false|C0015677;C1435181;C3887682|FAT1 protein, human;Fatty acid glycerol esters;Platelet Glycoprotein 4, human|fat
Finding|Gene or Genome|SIMPLE_SEGMENT|3313,3316|false|false|false|C0812278;C1366645;C1705088;C1708004;C3887682|CD36 gene;CD36 wt Allele;FAT1 gene;FAT1 wt Allele;Platelet Glycoprotein 4, human|fat
Finding|Receptor|SIMPLE_SEGMENT|3313,3316|false|false|false|C0812278;C1366645;C1705088;C1708004;C3887682|CD36 gene;CD36 wt Allele;FAT1 gene;FAT1 wt Allele;Platelet Glycoprotein 4, human|fat
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3313,3316|false|false|false|C0279453|doxorubicin/fluorouracil/triazinate protocol|fat
Finding|Functional Concept|SIMPLE_SEGMENT|3328,3332|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|3328,3348|false|false|false|C0262537|Left inguinal hernia|left inguinal hernia
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3333,3341|false|false|false|C0018246|Inguinal region|inguinal
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|3333,3348|false|false|false|C0019294|Hernia, Inguinal|inguinal hernia
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|3342,3348|false|false|false|C0019270|Hernia|hernia
Event|Event|SIMPLE_SEGMENT|3342,3348|false|false|false|||hernia
Event|Event|SIMPLE_SEGMENT|3352,3361|false|false|false|||unchanged
Finding|Finding|SIMPLE_SEGMENT|3352,3361|false|false|false|C0442739||unchanged
Event|Activity|SIMPLE_SEGMENT|3364,3375|false|false|false|C4321457|Examination|Examination
Event|Event|SIMPLE_SEGMENT|3364,3375|false|false|false|||Examination
Procedure|Health Care Activity|SIMPLE_SEGMENT|3364,3375|false|false|false|C0031809;C0582103|Medical Examination;Physical Examination|Examination
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3379,3383|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Anatomy|Tissue|SIMPLE_SEGMENT|3379,3391|false|false|false|C0225317|soft tissue|soft tissues
Anatomy|Tissue|SIMPLE_SEGMENT|3384,3391|false|false|false|C0040300|Body tissue|tissues
Event|Event|SIMPLE_SEGMENT|3392,3399|false|false|false|||reveals
Event|Event|SIMPLE_SEGMENT|3400,3409|false|false|false|||stranding
Event|Event|SIMPLE_SEGMENT|3414,3426|false|false|false|||subcutaneous
Finding|Functional Concept|SIMPLE_SEGMENT|3414,3426|false|false|false|C1522438|Subcutaneous Route of Administration|subcutaneous
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3428,3431|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3428,3431|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|SIMPLE_SEGMENT|3428,3431|false|false|false|C0001861;C3536832|Air (substance);air|air
Event|Event|SIMPLE_SEGMENT|3428,3431|false|false|false|||air
Finding|Finding|SIMPLE_SEGMENT|3428,3431|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|SIMPLE_SEGMENT|3428,3431|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|SIMPLE_SEGMENT|3428,3431|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3439,3443|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Anatomy|Tissue|SIMPLE_SEGMENT|3439,3451|false|false|false|C0225317|soft tissue|soft tissues
Anatomy|Tissue|SIMPLE_SEGMENT|3444,3451|false|false|false|C0040300|Body tissue|tissues
Anatomy|Cell Component|SIMPLE_SEGMENT|3462,3469|false|false|false|C1660780|midline cell component|midline
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3470,3475|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|3470,3475|false|false|false|C2003888|Lower (action)|lower
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3476,3484|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Event|Event|SIMPLE_SEGMENT|3476,3484|false|false|false|||anterior
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3486,3495|false|false|false|C0000726|Abdomen|abdominal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3486,3500|false|false|false|C0836916|Abdominal wall structure|abdominal wall
Event|Event|SIMPLE_SEGMENT|3511,3517|false|false|false|||larger
Event|Activity|SIMPLE_SEGMENT|3545,3556|false|false|false|C4321457|Examination|examination
Event|Event|SIMPLE_SEGMENT|3545,3556|false|false|false|||examination
Procedure|Health Care Activity|SIMPLE_SEGMENT|3545,3556|false|false|false|C0031809;C0582103|Medical Examination;Physical Examination|examination
Finding|Gene or Genome|SIMPLE_SEGMENT|3582,3585|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|SIMPLE_SEGMENT|3610,3615|false|false|false|||focus
Finding|Functional Concept|SIMPLE_SEGMENT|3610,3615|false|false|false|C1285542|Has focus|focus
Drug|Substance|SIMPLE_SEGMENT|3619,3624|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|3619,3624|false|false|false|C1546638|Fluid Specimen Code|fluid
Drug|Substance|SIMPLE_SEGMENT|3637,3645|false|false|false|C0520510|Materials|material
Event|Event|SIMPLE_SEGMENT|3637,3645|false|false|false|||material
Event|Event|SIMPLE_SEGMENT|3650,3657|false|false|false|||extends
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3668,3677|false|false|false|C0000726|Abdomen|abdominal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3668,3682|false|false|false|C0836916|Abdominal wall structure|abdominal wall
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3683,3694|false|false|false|C1995013|Set of muscles|musculature
Finding|Functional Concept|SIMPLE_SEGMENT|3707,3719|false|false|false|C1522438|Subcutaneous Route of Administration|subcutaneous
Anatomy|Tissue|SIMPLE_SEGMENT|3707,3727|false|false|false|C0278403|Subcutaneous Tissue|subcutaneous tissues
Anatomy|Tissue|SIMPLE_SEGMENT|3720,3727|false|false|false|C0040300|Body tissue|tissues
Event|Event|SIMPLE_SEGMENT|3745,3750|false|false|false|||drain
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3759,3767|false|false|false|C1548801|Body Site Modifier - External|external
Finding|Functional Concept|SIMPLE_SEGMENT|3759,3767|false|false|false|C0521134|External route|external
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|3768,3778|false|false|false|C0424290|Compulsive hoarding|collecting
Event|Event|SIMPLE_SEGMENT|3768,3778|false|false|false|||collecting
Finding|Functional Concept|SIMPLE_SEGMENT|3768,3778|false|false|false|C1516698|Collection (action)|collecting
Event|Event|SIMPLE_SEGMENT|3779,3785|false|false|false|||device
Finding|Functional Concept|SIMPLE_SEGMENT|3779,3785|false|false|false|C1550509|Participation Type - device|device
Drug|Substance|SIMPLE_SEGMENT|3800,3805|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|3800,3805|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|3800,3805|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|3806,3816|false|false|false|||collection
Finding|Conceptual Entity|SIMPLE_SEGMENT|3806,3816|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|3806,3816|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|3806,3816|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|3806,3816|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Event|Event|SIMPLE_SEGMENT|3820,3830|false|false|false|||identified
Event|Event|SIMPLE_SEGMENT|3834,3842|false|false|false|||indicate
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3843,3850|false|false|false|C0000833|Abscess|abscess
Finding|Intellectual Product|SIMPLE_SEGMENT|3843,3850|false|false|false|C1546533||abscess
Finding|Finding|SIMPLE_SEGMENT|3843,3860|false|false|false|C4014106|Abscess formation|abscess formation
Event|Event|SIMPLE_SEGMENT|3851,3860|false|false|false|||formation
Finding|Functional Concept|SIMPLE_SEGMENT|3851,3860|false|false|false|C1522492|Formation|formation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|3851,3860|false|false|false|C0220781|Anabolism|formation
Event|Event|SIMPLE_SEGMENT|3880,3888|false|false|false|||amenable
Event|Event|SIMPLE_SEGMENT|3892,3900|false|false|false|||drainage
Finding|Body Substance|SIMPLE_SEGMENT|3892,3900|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|SIMPLE_SEGMENT|3892,3900|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3892,3900|false|false|false|C0013103|Drainage procedure|drainage
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3916,3926|false|false|false|C0550215||appearance
Event|Event|SIMPLE_SEGMENT|3916,3926|false|false|false|||appearance
Procedure|Health Care Activity|SIMPLE_SEGMENT|3916,3926|false|false|false|C2051406|patient appearance regarding mental status exam|appearance
Event|Event|SIMPLE_SEGMENT|3928,3936|false|false|false|||suggests
Finding|Idea or Concept|SIMPLE_SEGMENT|3937,3946|false|false|false|C0549178|Continuous|continued
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3947,3957|false|false|false|C0007642|Cellulitis|cellulitis
Event|Event|SIMPLE_SEGMENT|3947,3957|false|false|false|||cellulitis
Finding|Finding|SIMPLE_SEGMENT|3947,3957|false|false|false|C2025995|cellulitis on exam (physical finding)|cellulitis
Event|Activity|SIMPLE_SEGMENT|3960,3971|false|false|false|C4321457|Examination|Examination
Event|Event|SIMPLE_SEGMENT|3960,3971|false|false|false|||Examination
Procedure|Health Care Activity|SIMPLE_SEGMENT|3960,3971|false|false|false|C0031809;C0582103|Medical Examination;Physical Examination|Examination
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3975,3982|false|false|false|C0262950;C4520924|Bone Tissue, Human;Skeletal bone|osseous
Anatomy|Tissue|SIMPLE_SEGMENT|3975,3982|false|false|false|C0262950;C4520924|Bone Tissue, Human;Skeletal bone|osseous
Event|Event|SIMPLE_SEGMENT|3994,4001|false|false|false|||reveals
Finding|Intellectual Product|SIMPLE_SEGMENT|4002,4006|false|false|false|C1547225|Mild Severity of Illness Code|mild
Event|Event|SIMPLE_SEGMENT|4007,4019|false|false|false|||degenerative
Finding|Functional Concept|SIMPLE_SEGMENT|4007,4019|false|false|false|C0011164;C1880269|Abnormal degeneration;biologic degeneration|degenerative
Finding|Pathologic Function|SIMPLE_SEGMENT|4007,4019|false|false|false|C0011164;C1880269|Abnormal degeneration;biologic degeneration|degenerative
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4021,4028|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|4021,4028|false|false|false|||disease
Event|Event|SIMPLE_SEGMENT|4056,4068|false|false|false|||unremarkable
Event|Event|SIMPLE_SEGMENT|4071,4081|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|4071,4081|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|4071,4081|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|4086,4092|false|false|false|C1547311|Patient Condition Code - Stable|Stable
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4093,4103|false|false|false|C0550215||appearance
Event|Event|SIMPLE_SEGMENT|4093,4103|false|false|false|||appearance
Procedure|Health Care Activity|SIMPLE_SEGMENT|4093,4103|false|false|false|C2051406|patient appearance regarding mental status exam|appearance
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4107,4114|false|false|false|C0227391|Sigmoid colon|sigmoid
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4107,4120|false|false|false|C0227391|Sigmoid colon|sigmoid colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4107,4120|false|false|false|C0153436;C0496864|Benign neoplasm of sigmoid colon;Malignant neoplasm of sigmoid colon|sigmoid colon
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4115,4120|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4115,4120|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4115,4120|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Finding|Finding|SIMPLE_SEGMENT|4115,4120|false|false|false|C0750873|COLON PROBLEM|colon
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4115,4132|false|false|false|C0852681|Large intestine anastomosis|colon anastomosis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4121,4132|false|false|false|C0500470|Anatomical anastomosis|anastomosis
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|4121,4132|false|false|false|C0332853|Anastomosis|anastomosis
Event|Event|SIMPLE_SEGMENT|4121,4132|false|false|false|||anastomosis
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4121,4132|false|false|false|C0677554||anastomosis
Event|Event|SIMPLE_SEGMENT|4142,4153|false|false|false|||obstruction
Finding|Finding|SIMPLE_SEGMENT|4142,4153|false|false|false|C0028778|Obstruction|obstruction
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4157,4164|false|false|false|C0000833|Abscess|abscess
Event|Event|SIMPLE_SEGMENT|4157,4164|false|false|false|||abscess
Finding|Intellectual Product|SIMPLE_SEGMENT|4157,4164|false|false|false|C1546533||abscess
Finding|Finding|SIMPLE_SEGMENT|4157,4174|false|false|false|C4014106|Abscess formation|abscess formation
Event|Event|SIMPLE_SEGMENT|4165,4174|false|false|false|||formation
Finding|Functional Concept|SIMPLE_SEGMENT|4165,4174|false|false|false|C1522492|Formation|formation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|4165,4174|false|false|false|C0220781|Anabolism|formation
Event|Event|SIMPLE_SEGMENT|4179,4188|false|false|false|||Stranding
Finding|Functional Concept|SIMPLE_SEGMENT|4193,4205|false|false|false|C1522438|Subcutaneous Route of Administration|subcutaneous
Finding|Finding|SIMPLE_SEGMENT|4193,4209|false|false|false|C3842127|Subcutaneous air|subcutaneous air
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4206,4209|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4206,4209|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|SIMPLE_SEGMENT|4206,4209|false|false|false|C0001861;C3536832|Air (substance);air|air
Event|Event|SIMPLE_SEGMENT|4206,4209|false|false|false|||air
Finding|Finding|SIMPLE_SEGMENT|4206,4209|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|SIMPLE_SEGMENT|4206,4209|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|SIMPLE_SEGMENT|4206,4209|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4220,4225|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|4220,4225|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4226,4235|false|false|false|C0000726|Abdomen|abdominal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4226,4240|false|false|false|C0836916|Abdominal wall structure|abdominal wall
Anatomy|Cell Component|SIMPLE_SEGMENT|4249,4256|false|false|false|C1660780|midline cell component|midline
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4269,4279|false|false|false|C0007642|Cellulitis|cellulitis
Event|Event|SIMPLE_SEGMENT|4269,4279|false|false|false|||cellulitis
Finding|Finding|SIMPLE_SEGMENT|4269,4279|false|false|false|C2025995|cellulitis on exam (physical finding)|cellulitis
Event|Event|SIMPLE_SEGMENT|4293,4301|false|false|false|||discrete
Drug|Substance|SIMPLE_SEGMENT|4316,4321|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|4316,4321|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|4316,4321|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|4322,4332|false|false|false|||collection
Finding|Conceptual Entity|SIMPLE_SEGMENT|4322,4332|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|4322,4332|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|4322,4332|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|4322,4332|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Event|Event|SIMPLE_SEGMENT|4338,4343|false|false|false|||study
Finding|Intellectual Product|SIMPLE_SEGMENT|4338,4343|false|false|false|C1705923|Study Object|study
Procedure|Research Activity|SIMPLE_SEGMENT|4338,4343|false|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|study
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4352,4358|false|false|false|C4255046||report
Event|Event|SIMPLE_SEGMENT|4352,4358|false|false|false|||report
Finding|Intellectual Product|SIMPLE_SEGMENT|4352,4358|false|false|false|C0684224|Report (document)|report
Procedure|Health Care Activity|SIMPLE_SEGMENT|4352,4358|false|false|false|C0700287|Reporting|report
Event|Event|SIMPLE_SEGMENT|4364,4372|false|false|false|||reviewed
Finding|Finding|SIMPLE_SEGMENT|4380,4385|false|false|false|C1551040|Encounter Special Courtesy - staff|staff
Event|Event|SIMPLE_SEGMENT|4386,4397|false|false|false|||radiologist
Finding|Intellectual Product|SIMPLE_SEGMENT|4386,4397|false|false|false|C1549438|Procedure Practitioner Identifier Code Type - Radiologist|radiologist
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|4427,4430|false|false|false|C0038817|Sunlight|SUN
Finding|Body Substance|SIMPLE_SEGMENT|4501,4506|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|4501,4506|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|4501,4506|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Finding|SIMPLE_SEGMENT|4501,4513|false|false|false|C0278030|Color of urine|URINE  COLOR
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4508,4513|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|COLOR
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|4508,4513|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|COLOR
Event|Event|SIMPLE_SEGMENT|4508,4513|false|false|false|||COLOR
Drug|Organic Chemical|SIMPLE_SEGMENT|4514,4519|false|false|false|C4047917|Cereal plant straw|Straw
Event|Event|SIMPLE_SEGMENT|4527,4532|false|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|4527,4532|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Body Substance|SIMPLE_SEGMENT|4552,4557|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|4552,4557|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|4552,4557|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4552,4564|false|false|false|C0018965|Hematuria|URINE  BLOOD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4559,4564|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4559,4564|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4559,4564|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Event|SIMPLE_SEGMENT|4565,4568|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|4565,4568|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4569,4576|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4569,4576|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4569,4576|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Finding|Finding|SIMPLE_SEGMENT|4577,4580|false|false|false|C5848551|Neg - answer|NEG
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4581,4588|false|false|false|C0033684|Proteins|PROTEIN
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4581,4588|false|false|false|C0033684|Proteins|PROTEIN
Event|Event|SIMPLE_SEGMENT|4581,4588|false|false|false|||PROTEIN
Finding|Conceptual Entity|SIMPLE_SEGMENT|4581,4588|false|false|false|C1521746|Protein Info|PROTEIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4581,4588|false|false|false|C0202202|Protein measurement|PROTEIN
Event|Event|SIMPLE_SEGMENT|4589,4592|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|4589,4592|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4594,4601|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|SIMPLE_SEGMENT|4594,4601|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4594,4601|false|false|false|C0017725|glucose|GLUCOSE
Event|Event|SIMPLE_SEGMENT|4594,4601|false|false|false|||GLUCOSE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4594,4601|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4594,4601|false|false|false|C0337438|Glucose measurement|GLUCOSE
Event|Event|SIMPLE_SEGMENT|4602,4605|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|4602,4605|false|false|false|C5848551|Neg - answer|NEG
Drug|Organic Chemical|SIMPLE_SEGMENT|4606,4612|false|false|false|C0022634|Ketones|KETONE
Event|Event|SIMPLE_SEGMENT|4613,4616|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|4613,4616|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4617,4626|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Drug|Organic Chemical|SIMPLE_SEGMENT|4617,4626|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4617,4626|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4617,4626|false|false|false|C0201913;C0863174|Bilirubin, total measurement;blood bilirubin level test|BILIRUBIN
Event|Event|SIMPLE_SEGMENT|4627,4630|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|4627,4630|false|false|false|C5848551|Neg - answer|NEG
Event|Event|SIMPLE_SEGMENT|4641,4644|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|4641,4644|false|false|false|C5848551|Neg - answer|NEG
Event|Event|SIMPLE_SEGMENT|4658,4661|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|4658,4661|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4676,4683|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|SIMPLE_SEGMENT|4676,4683|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4676,4683|false|false|false|C0017725|glucose|GLUCOSE
Event|Event|SIMPLE_SEGMENT|4676,4683|false|false|false|||GLUCOSE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4676,4683|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4676,4683|false|false|false|C0337438|Glucose measurement|GLUCOSE
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4689,4693|false|false|false|C0041942|urea|UREA
Drug|Organic Chemical|SIMPLE_SEGMENT|4689,4693|false|false|false|C0041942|urea|UREA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4689,4693|false|false|false|C0041942|urea|UREA
Event|Event|SIMPLE_SEGMENT|4689,4693|false|false|false|||UREA
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4689,4693|false|false|false|C0523961|Urea measurement|UREA
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4710,4716|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4710,4716|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4710,4716|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Event|Event|SIMPLE_SEGMENT|4710,4716|false|false|false|||SODIUM
Finding|Physiologic Function|SIMPLE_SEGMENT|4710,4716|false|false|false|C4553025|Sodium metabolic function|SODIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4710,4716|false|false|false|C0337443|Sodium measurement|SODIUM
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4722,4731|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4722,4731|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Food|SIMPLE_SEGMENT|4722,4731|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4722,4731|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4722,4731|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Event|Event|SIMPLE_SEGMENT|4722,4731|false|false|false|||POTASSIUM
Finding|Physiologic Function|SIMPLE_SEGMENT|4722,4731|false|false|false|C4553027|Potassium metabolic function|POTASSIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4722,4731|false|false|false|C0202194|Potassium measurement|POTASSIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4736,4744|false|false|false|C0008203;C0596019|Chlorides;chloride ion|CHLORIDE
Event|Event|SIMPLE_SEGMENT|4736,4744|false|false|false|||CHLORIDE
Finding|Physiologic Function|SIMPLE_SEGMENT|4736,4744|false|false|false|C4553021|Chloride metabolic function|CHLORIDE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4736,4744|false|false|false|C0201952|Chloride measurement|CHLORIDE
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4754,4757|false|false|false|C0007012|carbon dioxide|CO2
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4754,4757|false|false|false|C0007012|carbon dioxide|CO2
Event|Event|SIMPLE_SEGMENT|4754,4757|false|false|false|||CO2
Finding|Finding|SIMPLE_SEGMENT|4754,4757|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Finding|Gene or Genome|SIMPLE_SEGMENT|4754,4757|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4761,4766|false|false|false|C0003075|Anions|ANION
Event|Event|SIMPLE_SEGMENT|4761,4766|false|false|false|||ANION
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4761,4770|false|false|false|C0003074|Anion Gap|ANION GAP
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4761,4770|false|false|false|C1509129|Anion gap result|ANION GAP
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4761,4770|false|false|false|C0201889;C2189246|Anion gap measurement;blood anion gap (lab test)|ANION GAP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4767,4770|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4767,4770|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Event|Event|SIMPLE_SEGMENT|4767,4770|false|false|false|||GAP
Finding|Gene or Genome|SIMPLE_SEGMENT|4767,4770|false|false|false|C1419277;C2984552|RASA1 gene;RASA1 wt Allele|GAP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4820,4823|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4820,4823|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|4820,4823|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|4820,4823|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|4820,4823|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|4820,4823|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|4820,4823|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4820,4823|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4824,4828|false|false|false|C0376147|SGPT - Glutamate pyruvate transaminase|SGPT
Drug|Enzyme|SIMPLE_SEGMENT|4824,4828|false|false|false|C0376147|SGPT - Glutamate pyruvate transaminase|SGPT
Event|Event|SIMPLE_SEGMENT|4824,4828|false|false|false|||SGPT
Finding|Gene or Genome|SIMPLE_SEGMENT|4824,4828|false|false|false|C1415274|GPT gene|SGPT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4824,4828|false|false|false|C0036828|Serum Alanine Transaminase Test|SGPT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4833,4836|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4833,4836|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4833,4836|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4833,4836|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|4833,4836|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|4833,4836|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|4833,4836|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4837,4841|false|false|false|C0242192|SGOT - Glutamate oxaloacetate transaminase|SGOT
Drug|Enzyme|SIMPLE_SEGMENT|4837,4841|false|false|false|C0242192|SGOT - Glutamate oxaloacetate transaminase|SGOT
Event|Event|SIMPLE_SEGMENT|4837,4841|false|false|false|||SGOT
Finding|Gene or Genome|SIMPLE_SEGMENT|4837,4841|false|false|false|C1415181|GOT1 gene|SGOT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4837,4841|false|false|false|C0201899|Aspartate aminotransferase measurement|SGOT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4846,4849|false|false|false|C1663627|ALK protein, human|ALK
Drug|Enzyme|SIMPLE_SEGMENT|4846,4849|false|false|false|C1663627|ALK protein, human|ALK
Event|Event|SIMPLE_SEGMENT|4846,4849|false|false|false|||ALK
Finding|Gene or Genome|SIMPLE_SEGMENT|4846,4849|false|false|false|C1332080;C1663627;C1704943|ALK gene;ALK protein, human;ALK wt Allele|ALK
Finding|Receptor|SIMPLE_SEGMENT|4846,4849|false|false|false|C1332080;C1663627;C1704943|ALK gene;ALK protein, human;ALK wt Allele|ALK
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4846,4854|false|false|false|C0002059|Alkaline Phosphatase|ALK PHOS
Drug|Enzyme|SIMPLE_SEGMENT|4846,4854|false|false|false|C0002059|Alkaline Phosphatase|ALK PHOS
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4846,4854|false|false|false|C0201850|Alkaline phosphatase measurement|ALK PHOS
Event|Event|SIMPLE_SEGMENT|4850,4854|false|false|false|||PHOS
Event|Event|SIMPLE_SEGMENT|4859,4862|false|false|false|||TOT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4887,4893|false|false|false|C0023764|lipase|LIPASE
Drug|Enzyme|SIMPLE_SEGMENT|4887,4893|false|false|false|C0023764|lipase|LIPASE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4887,4893|false|false|false|C0023764|lipase|LIPASE
Event|Event|SIMPLE_SEGMENT|4887,4893|false|false|false|||LIPASE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4887,4893|false|false|false|C0373670|Lipase measurement|LIPASE
Anatomy|Cell|SIMPLE_SEGMENT|4912,4915|false|false|false|C0023516|Leukocytes|WBC
Event|Event|SIMPLE_SEGMENT|4912,4915|false|false|false|||WBC
Anatomy|Cell|SIMPLE_SEGMENT|4923,4926|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4923,4926|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4923,4926|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4933,4936|false|false|false|C0019046|Hemoglobin|HGB
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4933,4936|false|false|false|C0019046|Hemoglobin|HGB
Finding|Gene or Genome|SIMPLE_SEGMENT|4933,4936|false|false|false|C1424337|CYGB gene|HGB
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4933,4936|false|false|false|C0019029|Hemoglobin concentration|HGB
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4942,4945|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4942,4945|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Disorder|Virus|SIMPLE_SEGMENT|4953,4956|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|4953,4956|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4953,4956|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4953,4956|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4953,4956|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|4960,4963|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4960,4963|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|4960,4963|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|4960,4963|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|4960,4963|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4960,4963|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|4969,4973|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4969,4973|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Event|Event|SIMPLE_SEGMENT|5002,5007|false|false|false|||NEUTS
Finding|Body Substance|SIMPLE_SEGMENT|5014,5020|false|false|false|C0024202|Lymph|LYMPHS
Drug|Antibiotic|SIMPLE_SEGMENT|5027,5032|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5027,5032|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Organic Chemical|SIMPLE_SEGMENT|5027,5032|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5037,5040|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|EOS
Event|Event|SIMPLE_SEGMENT|5037,5040|false|false|false|||EOS
Finding|Gene or Genome|SIMPLE_SEGMENT|5037,5040|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|EOS
Event|Event|SIMPLE_SEGMENT|5070,5073|false|false|false|||PLT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5070,5073|false|false|false|C0201617|Primed lymphocyte test|PLT
Finding|Intellectual Product|SIMPLE_SEGMENT|5088,5093|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|5094,5102|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5094,5109|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|5094,5109|false|false|false|C0489547|Hospital course|Hospital Course
Event|Event|SIMPLE_SEGMENT|5115,5123|false|false|false|||Admitted
Procedure|Health Care Activity|SIMPLE_SEGMENT|5115,5123|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admitted
Event|Event|SIMPLE_SEGMENT|5164,5167|false|false|false|||NPO
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5164,5167|false|false|false|C0419179|NPO - Nothing by mouth|NPO
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5174,5177|false|false|false|C0016520|Structure of interventricular foramen|IVF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5174,5177|false|false|false|C2751898|Ventricular Fibrillation, Paroxysmal Familial, 1|IVF
Event|Event|SIMPLE_SEGMENT|5174,5177|false|false|false|||IVF
Finding|Gene or Genome|SIMPLE_SEGMENT|5174,5177|false|false|false|C1419864;C4321334|SCN5A gene;SCN5A wt Allele|IVF
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5174,5177|false|false|false|C0015915;C0872104|Assisted Reproductive Technologies;Fertilization in Vitro|IVF
Event|Event|SIMPLE_SEGMENT|5178,5191|false|false|false|||resuscitation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5178,5191|false|false|false|C0035273|Resuscitation (procedure)|resuscitation
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5196,5205|false|false|false|C0000726|Abdomen|abdominal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5206,5212|false|false|false|C0030797|Pelvis|pelvic
Event|Event|SIMPLE_SEGMENT|5213,5215|false|false|false|||CT
Event|Event|SIMPLE_SEGMENT|5230,5242|false|false|false|||demonstrated
Finding|Intellectual Product|SIMPLE_SEGMENT|5245,5251|false|false|false|C1547311|Patient Condition Code - Stable|stable
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5252,5259|false|false|false|C0227391|Sigmoid colon|sigmoid
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5260,5271|false|false|false|C0500470|Anatomical anastomosis|anastomosis
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|5260,5271|false|false|false|C0332853|Anastomosis|anastomosis
Event|Event|SIMPLE_SEGMENT|5260,5271|false|false|false|||anastomosis
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5260,5271|false|false|false|C0677554||anastomosis
Drug|Substance|SIMPLE_SEGMENT|5284,5289|true|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|5284,5289|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|5284,5289|true|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|5291,5302|false|false|false|||collections
Event|Event|SIMPLE_SEGMENT|5306,5310|false|false|false|||free
Finding|Functional Concept|SIMPLE_SEGMENT|5306,5310|false|false|false|C0332296|Free of (attribute)|free
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5311,5314|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5311,5314|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|SIMPLE_SEGMENT|5311,5314|false|false|false|C0001861;C3536832|Air (substance);air|air
Event|Event|SIMPLE_SEGMENT|5311,5314|false|false|false|||air
Finding|Finding|SIMPLE_SEGMENT|5311,5314|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|SIMPLE_SEGMENT|5311,5314|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|SIMPLE_SEGMENT|5311,5314|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Body Substance|SIMPLE_SEGMENT|5342,5347|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|SIMPLE_SEGMENT|5342,5347|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|SIMPLE_SEGMENT|5342,5347|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5342,5354|false|false|false|C0232856;C0489132||urine output
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5342,5354|false|false|false|C2094175|monitoring of urine output for fluid balance|urine output
Event|Event|SIMPLE_SEGMENT|5348,5354|false|false|false|||output
Finding|Conceptual Entity|SIMPLE_SEGMENT|5348,5354|false|false|false|C1709366|system output|output
Procedure|Health Care Activity|SIMPLE_SEGMENT|5348,5354|false|false|false|C3251815|Measurement of fluid output|output
Event|Event|SIMPLE_SEGMENT|5356,5365|false|false|false|||increased
Event|Event|SIMPLE_SEGMENT|5372,5377|false|false|false|||foley
Event|Event|SIMPLE_SEGMENT|5386,5392|false|false|false|||placed
Finding|Intellectual Product|SIMPLE_SEGMENT|5406,5414|false|false|false|C1720529|Constant - dosing instruction fragment|constant
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5422,5428|false|false|false|C0489144||stools
Event|Event|SIMPLE_SEGMENT|5422,5428|false|false|false|||stools
Finding|Body Substance|SIMPLE_SEGMENT|5422,5428|false|false|false|C0015733|Feces|stools
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5430,5435|false|false|false|C0040549|Toxin|toxin
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|5430,5435|false|false|false|C0040549|Toxin|toxin
Event|Event|SIMPLE_SEGMENT|5436,5443|false|false|false|||screens
Event|Event|SIMPLE_SEGMENT|5459,5463|false|false|false|||sent
Event|Event|SIMPLE_SEGMENT|5468,5476|false|false|false|||returned
Event|Event|SIMPLE_SEGMENT|5477,5485|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|5477,5485|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|5477,5485|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5477,5485|false|false|false|C5237010|Expression Negative|negative
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5492,5495|false|false|false|C2713652|HDAC2 protein, human|HD2
Drug|Enzyme|SIMPLE_SEGMENT|5492,5495|false|false|false|C2713652|HDAC2 protein, human|HD2
Event|Event|SIMPLE_SEGMENT|5492,5495|false|false|false|||HD2
Finding|Gene or Genome|SIMPLE_SEGMENT|5492,5495|false|false|false|C1706172|HDAC2 wt Allele|HD2
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5501,5507|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|5501,5507|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|5501,5507|false|false|false|C0027497|Nausea|nausea
Event|Event|SIMPLE_SEGMENT|5508,5517|false|false|false|||persisted
Procedure|Health Care Activity|SIMPLE_SEGMENT|5523,5533|false|false|false|C0744396|GI CONSULT|GI consult
Event|Event|SIMPLE_SEGMENT|5526,5533|false|false|false|||consult
Procedure|Health Care Activity|SIMPLE_SEGMENT|5526,5533|false|false|false|C0009818|Consultation|consult
Event|Event|SIMPLE_SEGMENT|5538,5546|false|false|false|||obtained
Event|Occupational Activity|SIMPLE_SEGMENT|5557,5564|false|false|false|C0557854|Services|service
Finding|Idea or Concept|SIMPLE_SEGMENT|5557,5564|false|false|false|C3245478|ActInformationPrivacyReason - service|service
Event|Event|SIMPLE_SEGMENT|5565,5573|false|false|false|||believed
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5578,5584|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|5578,5584|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|5578,5584|false|false|false|C0027497|Nausea|nausea
Drug|Organic Chemical|SIMPLE_SEGMENT|5591,5598|false|false|false|C0163712|Relate - vinyl resin|related
Event|Event|SIMPLE_SEGMENT|5591,5598|false|false|false|||related
Finding|Finding|SIMPLE_SEGMENT|5591,5598|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|SIMPLE_SEGMENT|5591,5598|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5602,5610|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|SIMPLE_SEGMENT|5602,5610|false|false|false|||baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|5602,5610|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|SIMPLE_SEGMENT|5611,5617|false|false|false|||reflux
Finding|Pathologic Function|SIMPLE_SEGMENT|5611,5617|false|false|false|C0232483|Reflux|reflux
Event|Event|SIMPLE_SEGMENT|5619,5630|false|false|false|||exacerbated
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|5665,5670|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Event|Event|SIMPLE_SEGMENT|5665,5670|false|false|false|||wound
Finding|Body Substance|SIMPLE_SEGMENT|5665,5670|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|SIMPLE_SEGMENT|5665,5670|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|SIMPLE_SEGMENT|5665,5670|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Pathologic Function|SIMPLE_SEGMENT|5665,5680|false|false|false|C0043241|Wound Infection|wound infection
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5671,5680|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|5671,5680|false|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|5671,5680|false|false|false|C3714514|Infection|infection
Event|Event|SIMPLE_SEGMENT|5694,5709|false|false|false|||recommendations
Finding|Idea or Concept|SIMPLE_SEGMENT|5694,5709|false|false|false|C0034866|Recommendation|recommendations
Event|Event|SIMPLE_SEGMENT|5719,5726|false|false|false|||started
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5733,5740|false|false|false|C0003138;C0003216|Antacids;Anti-Ulcer Agent|antacid
Event|Event|SIMPLE_SEGMENT|5733,5740|false|false|false|||antacid
Finding|Physiologic Function|SIMPLE_SEGMENT|5733,5740|false|false|false|C1383090|Antacid [PE]|antacid
Event|Event|SIMPLE_SEGMENT|5751,5760|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|5751,5760|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|5751,5760|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|5751,5760|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|5751,5760|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|5770,5776|false|false|false|||follow
Event|Event|SIMPLE_SEGMENT|5810,5819|false|false|false|||determine
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5833,5839|false|false|false|C5889824||status
Event|Event|SIMPLE_SEGMENT|5833,5839|false|false|false|||status
Finding|Idea or Concept|SIMPLE_SEGMENT|5833,5839|false|false|false|C1546481|What subject filter - Status|status
Event|Event|SIMPLE_SEGMENT|5852,5861|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|5852,5861|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|5852,5861|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|5852,5861|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|5852,5861|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|5872,5882|false|false|false|||tolerating
Finding|Finding|SIMPLE_SEGMENT|5885,5888|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|SIMPLE_SEGMENT|5885,5888|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5885,5901|false|false|false|C0425404|Low residue diet|low residue diet
Finding|Conceptual Entity|SIMPLE_SEGMENT|5889,5896|false|false|false|C1709915|Residue|residue
Drug|Food|SIMPLE_SEGMENT|5897,5901|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|SIMPLE_SEGMENT|5897,5901|false|false|false|||diet
Finding|Functional Concept|SIMPLE_SEGMENT|5897,5901|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|SIMPLE_SEGMENT|5897,5901|false|false|false|C0012159|Diet therapy|diet
Event|Event|SIMPLE_SEGMENT|5906,5910|false|false|false|||able
Finding|Finding|SIMPLE_SEGMENT|5906,5910|false|false|false|C1299581|Able (qualifier value)|able
Event|Event|SIMPLE_SEGMENT|5914,5921|false|false|false|||hydrate
Event|Event|SIMPLE_SEGMENT|5935,5944|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|5935,5944|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|5935,5944|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|5935,5944|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|5935,5944|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|5935,5956|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5945,5956|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5945,5956|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|5945,5956|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|5945,5956|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|5961,5973|false|false|false|C1099456|escitalopram|Escitalopram
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5961,5973|false|false|false|C1099456|escitalopram|Escitalopram
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5980,5986|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6000,6006|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|6000,6006|false|false|false|||Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6034,6040|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|SIMPLE_SEGMENT|6045,6052|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|6060,6072|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6060,6072|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6079,6085|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|6079,6085|false|false|false|||Tablet
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6087,6094|false|false|false|C1545665|Views delayed|Delayed
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6087,6102|false|false|false|C1707664|Delayed Release Dosage Form|Delayed Release
Event|Event|SIMPLE_SEGMENT|6095,6102|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|6095,6102|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|6095,6102|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6095,6102|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Event|Event|SIMPLE_SEGMENT|6110,6113|false|false|false|||Sig
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6124,6130|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|6124,6130|false|false|false|||Tablet
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6132,6139|false|false|false|C1545665|Views delayed|Delayed
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6132,6147|false|false|false|C1707664|Delayed Release Dosage Form|Delayed Release
Event|Event|SIMPLE_SEGMENT|6140,6147|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|6140,6147|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|6140,6147|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6140,6147|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6190,6196|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|6190,6196|false|false|false|||Tablet
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6198,6205|false|false|false|C1545665|Views delayed|Delayed
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6198,6213|false|false|false|C1707664|Delayed Release Dosage Form|Delayed Release
Event|Event|SIMPLE_SEGMENT|6206,6213|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|6206,6213|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|6206,6213|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6206,6213|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Finding|Idea or Concept|SIMPLE_SEGMENT|6225,6232|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|6240,6250|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6240,6250|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Organic Chemical|SIMPLE_SEGMENT|6240,6254|false|false|false|C0700466|ranitidine hydrochloride|Ranitidine HCl
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6240,6254|false|false|false|C0700466|ranitidine hydrochloride|Ranitidine HCl
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6251,6254|false|false|false|C0023443|Hairy Cell Leukemia|HCl
Drug|Immunologic Factor|SIMPLE_SEGMENT|6251,6254|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Inorganic Chemical|SIMPLE_SEGMENT|6251,6254|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6251,6254|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Event|Event|SIMPLE_SEGMENT|6251,6254|false|false|false|||HCl
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6262,6268|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6282,6288|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|6282,6288|false|false|false|||Tablet
Event|Event|SIMPLE_SEGMENT|6300,6307|false|false|false|||bedtime
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6319,6325|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|SIMPLE_SEGMENT|6330,6337|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|6345,6356|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6345,6356|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|SIMPLE_SEGMENT|6345,6356|false|false|false|||Fluticasone
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6374,6379|false|false|false|C1154182|Spray Dosage Form|Spray
Event|Activity|SIMPLE_SEGMENT|6374,6379|false|false|false|C2003858|Spray (action)|Spray
Event|Event|SIMPLE_SEGMENT|6374,6379|false|false|false|||Spray
Finding|Functional Concept|SIMPLE_SEGMENT|6374,6379|false|false|false|C4521772|Spray (administration method)|Spray
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6374,6391|false|false|false|C1710170|SPRAY, SUSPENSION|Spray, Suspension
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6381,6391|false|false|false|C0038960;C1382107|Suspension substance;Suspensions|Suspension
Drug|Substance|SIMPLE_SEGMENT|6381,6391|false|false|false|C0038960;C1382107|Suspension substance;Suspensions|Suspension
Event|Event|SIMPLE_SEGMENT|6381,6391|false|false|false|||Suspension
Finding|Functional Concept|SIMPLE_SEGMENT|6381,6391|false|false|false|C1705537|Suspension (action)|Suspension
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6406,6411|false|false|false|C1154182|Spray Dosage Form|Spray
Event|Activity|SIMPLE_SEGMENT|6406,6411|false|false|false|C2003858|Spray (action)|Spray
Event|Event|SIMPLE_SEGMENT|6406,6411|false|false|false|||Spray
Finding|Functional Concept|SIMPLE_SEGMENT|6406,6411|false|false|false|C4521772|Spray (administration method)|Spray
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6412,6417|false|false|false|C0028429||Nasal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6412,6417|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Organic Chemical|SIMPLE_SEGMENT|6412,6417|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6412,6417|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Finding|Finding|SIMPLE_SEGMENT|6412,6417|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Functional Concept|SIMPLE_SEGMENT|6412,6417|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Event|Event|SIMPLE_SEGMENT|6418,6423|false|false|false|||DAILY
Finding|Idea or Concept|SIMPLE_SEGMENT|6443,6450|false|false|false|C0807726|refill|Refills
Event|Event|SIMPLE_SEGMENT|6458,6467|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|6458,6467|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6458,6467|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6458,6467|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6458,6467|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6458,6479|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|6458,6479|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6468,6479|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|6468,6479|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|6468,6479|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|SIMPLE_SEGMENT|6481,6485|false|false|false|||Home
Finding|Idea or Concept|SIMPLE_SEGMENT|6481,6485|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|6481,6485|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|6481,6485|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|SIMPLE_SEGMENT|6491,6498|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|6491,6498|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|SIMPLE_SEGMENT|6501,6509|false|false|false|||Facility
Finding|Intellectual Product|SIMPLE_SEGMENT|6501,6509|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|SIMPLE_SEGMENT|6517,6526|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|6517,6526|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6517,6526|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6517,6526|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6517,6526|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|6517,6536|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6527,6536|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|6527,6536|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|6527,6536|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|6527,6536|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6527,6536|false|false|false|C0011900|Diagnosis|Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6538,6544|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|6538,6544|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|6538,6544|false|false|false|C0027497|Nausea|nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|6538,6557|false|false|false|C0027498|Nausea and vomiting|nausea and vomiting
Event|Event|SIMPLE_SEGMENT|6549,6557|false|false|false|||vomiting
Finding|Sign or Symptom|SIMPLE_SEGMENT|6549,6557|false|false|false|C0042963|Vomiting|vomiting
Event|Event|SIMPLE_SEGMENT|6561,6570|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|6561,6570|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6561,6570|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6561,6570|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6561,6570|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6571,6580|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6571,6580|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|6571,6580|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|6571,6580|false|false|false|C1705253|Logical Condition|Condition
Procedure|Health Care Activity|SIMPLE_SEGMENT|6582,6590|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6591,6603|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|6591,6603|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|6591,6603|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

