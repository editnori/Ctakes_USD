 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|25,29
No|30,32
:|32,33
_|36,37
_|37,38
_|38,39
<EOL>|39,40
<EOL>|41,42
Admission|42,51
Date|52,56
:|56,57
_|59,60
_|60,61
_|61,62
Discharge|76,85
Date|86,90
:|90,91
_|94,95
_|95,96
_|96,97
<EOL>|97,98
<EOL>|99,100
Date|100,104
of|105,107
Birth|108,113
:|113,114
_|116,117
_|117,118
_|118,119
Sex|132,135
:|135,136
F|139,140
<EOL>|140,141
<EOL>|142,143
Service|143,150
:|150,151
MEDICINE|152,160
<EOL>|160,161
<EOL>|162,163
Allergies|163,172
:|172,173
<EOL>|174,175
IV|175,177
Dye|178,181
,|181,182
Iodine|183,189
Containing|190,200
Contrast|201,209
Media|210,215
/|216,217
Oxycodone|218,227
/|228,229
<EOL>|230,231
cilostazol|231,241
/|242,243
Varenicline|244,255
<EOL>|255,256
<EOL>|257,258
Attending|258,267
:|267,268
_|269,270
_|270,271
_|271,272
.|272,273
<EOL>|273,274
<EOL>|275,276
Chief|276,281
Complaint|282,291
:|291,292
<EOL>|292,293
Dyspnea|293,300
<EOL>|301,302
<EOL>|303,304
Major|304,309
Surgical|310,318
or|319,321
Invasive|322,330
Procedure|331,340
:|340,341
<EOL>|341,342
None|342,346
.|346,347
<EOL>|347,348
<EOL>|348,349
<EOL>|350,351
History|351,358
of|359,361
Present|362,369
Illness|370,377
:|377,378
<EOL>|378,379
_|379,380
_|380,381
_|381,382
y|383,384
/|384,385
o|385,386
F|387,388
with|389,393
asthma|394,400
,|400,401
CAD|402,405
s|406,407
/|407,408
p|408,409
stents|410,416
(|417,418
reported|418,426
by|427,429
patient|430,437
)|437,438
,|438,439
<EOL>|440,441
COPD|441,445
,|445,446
PAD|447,450
,|450,451
HTN|452,455
,|455,456
who|457,460
presents|461,469
with|470,474
shortness|475,484
of|485,487
breath|488,494
.|494,495
The|496,499
<EOL>|500,501
patient|501,508
was|509,512
sitting|513,520
at|521,523
home|524,528
ewhen|529,534
she|535,538
suddenly|539,547
felt|548,552
short|553,558
of|559,561
<EOL>|562,563
breath|563,569
.|569,570
She|571,574
drank|575,580
some|581,585
water|586,591
and|592,595
took|596,600
nebulizers|601,611
which|612,617
she|618,621
felt|622,626
<EOL>|627,628
helped|628,634
some|635,639
.|639,640
She|641,644
also|645,649
has|650,653
noticed|654,661
hoarseness|662,672
of|673,675
her|676,679
voice|680,685
.|685,686
<EOL>|688,689
She|689,692
presented|693,702
because|703,710
her|711,714
symptoms|715,723
have|724,728
gotten|729,735
worse|736,741
throughout|742,752
<EOL>|753,754
the|754,757
day|758,761
.|761,762
Denies|763,769
fever|770,775
/|775,776
chills|776,782
,|782,783
sore|784,788
throat|789,795
.|795,796
Says|797,801
she|802,805
does|806,810
have|811,815
a|816,817
<EOL>|818,819
cough|819,824
from|825,829
asthma|830,836
and|837,840
noticed|841,848
increased|849,858
wheezing|859,867
.|867,868
She|869,872
had|873,876
an|877,879
<EOL>|880,881
episode|881,888
of|889,891
substernal|892,902
chest|903,908
pain|909,913
this|914,918
morning|919,926
that|927,931
lasted|932,938
_|939,940
_|940,941
_|941,942
<EOL>|943,944
minutes|944,951
that|952,956
was|957,960
nonextertional|961,975
.|975,976
No|977,979
radiation|980,989
to|990,992
jaw|993,996
,|996,997
arm|998,1001
,|1001,1002
or|1003,1005
<EOL>|1006,1007
back|1007,1011
.|1011,1012
It|1013,1015
resolved|1016,1024
without|1025,1032
any|1033,1036
intervention|1037,1049
.|1049,1050
She|1051,1054
reported|1055,1063
some|1064,1068
<EOL>|1069,1070
leg|1070,1073
swelling|1074,1082
but|1083,1086
says|1087,1091
that|1092,1096
has|1097,1100
resolved|1101,1109
.|1109,1110
She|1111,1114
denies|1115,1121
PND|1122,1125
,|1125,1126
<EOL>|1127,1128
orthopnea|1128,1137
.|1137,1138
<EOL>|1140,1141
<EOL>|1141,1142
In|1142,1144
the|1145,1148
ED|1149,1151
,|1151,1152
initial|1153,1160
vitals|1161,1167
were|1168,1172
:|1172,1173
<EOL>|1173,1174
96.5|1174,1178
77|1179,1181
143|1182,1185
/|1185,1186
68|1186,1188
22|1189,1191
97|1192,1194
%|1194,1195
RA|1196,1198
<EOL>|1200,1201
<EOL>|1201,1202
Labs|1202,1206
were|1207,1211
notable|1212,1219
for|1220,1223
:|1223,1224
<EOL>|1225,1226
-|1226,1227
Labs|1228,1232
were|1233,1237
significant|1238,1249
for|1250,1253
neg|1254,1257
trop|1258,1262
x1|1263,1265
,|1265,1266
normal|1267,1273
CBC|1274,1277
,|1277,1278
normal|1279,1285
<EOL>|1286,1287
chemistry|1287,1296
panel|1297,1302
.|1302,1303
<EOL>|1305,1306
-|1306,1307
CXR|1308,1311
was|1312,1315
negative|1316,1324
.|1324,1325
EKG|1326,1329
shows|1330,1335
LBBB|1336,1340
consistent|1341,1351
with|1352,1356
prior|1357,1362
.|1362,1363
<EOL>|1365,1366
<EOL>|1366,1367
Patient|1367,1374
was|1375,1378
given|1379,1384
:|1384,1385
<EOL>|1385,1386
The|1386,1389
patient|1390,1397
was|1398,1401
given|1402,1407
albuterol|1408,1417
/|1417,1418
ipra|1418,1422
nebs|1423,1427
,|1427,1428
prednisone|1429,1439
60|1440,1442
mg|1443,1445
x|1446,1447
1|1448,1449
.|1449,1450
<EOL>|1450,1451
<EOL>|1451,1452
Consults|1452,1460
:|1460,1461
<EOL>|1461,1462
ED|1462,1464
spoke|1465,1470
with|1471,1475
Dr.|1476,1479
_|1480,1481
_|1481,1482
_|1482,1483
wanted|1484,1490
admission|1491,1500
for|1501,1504
stress|1505,1511
test|1512,1516
<EOL>|1517,1518
in|1518,1520
morning|1521,1528
.|1528,1529
ED|1530,1532
did|1533,1536
not|1537,1540
feel|1541,1545
she|1546,1549
is|1550,1552
CDU|1553,1556
candidate|1557,1566
given|1567,1572
she|1573,1576
is|1577,1579
on|1580,1582
<EOL>|1583,1584
theophylline|1584,1596
and|1597,1600
would|1601,1606
require|1607,1614
more|1615,1619
than|1620,1624
one|1625,1628
day|1629,1632
in|1633,1635
hospital|1636,1644
.|1644,1645
<EOL>|1647,1648
<EOL>|1648,1649
Vitals|1649,1655
prior|1656,1661
to|1662,1664
transfer|1665,1673
were|1674,1678
:|1678,1679
71|1680,1682
149|1683,1686
/|1686,1687
73|1687,1689
20|1690,1692
94|1693,1695
%|1695,1696
RA|1697,1699
<EOL>|1701,1702
On|1702,1704
arrival|1705,1712
to|1713,1715
floor|1716,1721
,|1721,1722
she|1723,1726
denies|1727,1733
chest|1734,1739
pain|1740,1744
.|1744,1745
Shortness|1746,1755
of|1756,1758
breath|1759,1765
<EOL>|1766,1767
has|1767,1770
improved|1771,1779
after|1780,1785
receiving|1786,1795
inhalers|1796,1804
.|1804,1805
<EOL>|1805,1806
<EOL>|1807,1808
Past|1808,1812
Medical|1813,1820
History|1821,1828
:|1828,1829
<EOL>|1829,1830
ASTHMA|1830,1836
/|1836,1837
COPD|1837,1841
/|1841,1842
Tobacco|1842,1849
use|1850,1853
,|1853,1854
Peripheral|1855,1865
Arterial|1866,1874
disease|1875,1882
s|1883,1884
/|1884,1885
p|1885,1886
recent|1887,1893
<EOL>|1894,1895
common|1895,1901
iliac|1902,1907
stenting|1908,1916
,|1916,1917
ATRIAL|1918,1924
TACHYCARDIA|1925,1936
,|1936,1937
ATYPICAL|1938,1946
CHEST|1947,1952
PAIN|1953,1957
,|1957,1958
<EOL>|1959,1960
CERVICAL|1960,1968
RADICULITIS|1969,1980
,|1980,1981
CERVICAL|1982,1990
SPONDYLOSIS|1991,2002
,|2002,2003
CORONARY|2004,2012
ARTERY|2013,2019
<EOL>|2020,2021
DISEASE|2021,2028
<EOL>|2030,2031
HEADACHE|2031,2039
,|2039,2040
HIP|2041,2044
REPLACEMENT|2045,2056
,|2056,2057
HYPERLIPIDEMIA|2058,2072
,|2072,2073
HYPERTENSION|2074,2086
,|2086,2087
<EOL>|2088,2089
OSTEOARTHRITIS|2089,2103
,|2103,2104
HERPES|2105,2111
ZOSTER|2112,2118
,|2118,2119
TOBACCO|2120,2127
ABUSE|2128,2133
,|2133,2134
ATRIAL|2135,2141
<EOL>|2142,2143
FIBRILLATION|2143,2155
<EOL>|2157,2158
ANXIETY|2158,2165
,|2165,2166
GASTROINTESTINAL|2166,2182
BLEEDING|2183,2191
,|2191,2192
OSTEOARTHRITIS|2193,2207
,|2207,2208
<EOL>|2209,2210
ATHEROSCLEROTIC|2210,2225
CARDIOVASCULAR|2226,2240
DISEASE|2241,2248
,|2248,2249
PERIPHERAL|2250,2260
VASCULAR|2261,2269
<EOL>|2270,2271
DISEASE|2271,2278
,|2278,2279
CATARACT|2280,2288
SURGERY|2289,2296
_|2297,2298
_|2298,2299
_|2299,2300
<EOL>|2302,2303
Surgery|2303,2310
:|2310,2311
<EOL>|2313,2314
BILATERAL|2314,2323
COMMON|2324,2330
ILIAC|2331,2336
ARTERY|2337,2343
STENTING|2344,2352
_|2353,2354
_|2354,2355
_|2355,2356
<EOL>|2358,2359
BUNIONECTOMY|2359,2371
<EOL>|2373,2374
HIP|2374,2377
REPLACEMENT|2378,2389
<EOL>|2391,2392
PRIOR|2392,2397
CESAREAN|2398,2406
SECTION|2407,2414
<EOL>|2416,2417
GANGLION|2417,2425
CYST|2426,2430
<EOL>|2430,2431
<EOL>|2432,2433
Social|2433,2439
History|2440,2447
:|2447,2448
<EOL>|2448,2449
_|2449,2450
_|2450,2451
_|2451,2452
<EOL>|2452,2453
Family|2453,2459
History|2460,2467
:|2467,2468
<EOL>|2468,2469
Mother|2469,2475
:|2475,2476
_|2477,2478
_|2478,2479
_|2479,2480
,|2480,2481
HTN|2482,2485
<EOL>|2487,2488
Father|2488,2494
:|2494,2495
_|2496,2497
_|2497,2498
_|2498,2499
CA|2500,2502
<EOL>|2504,2505
Brother|2505,2512
:|2512,2513
CA|2514,2516
?|2516,2517
<EOL>|2519,2520
Brother|2520,2527
:|2527,2528
_|2529,2530
_|2530,2531
_|2531,2532
<EOL>|2533,2534
<EOL>|2535,2536
Physical|2536,2544
_|2545,2546
_|2546,2547
_|2547,2548
:|2548,2549
<EOL>|2549,2550
=|2550,2551
=|2551,2552
=|2552,2553
=|2553,2554
=|2554,2555
=|2555,2556
=|2556,2557
=|2557,2558
=|2558,2559
=|2559,2560
=|2560,2561
=|2561,2562
=|2562,2563
=|2563,2564
=|2564,2565
=|2565,2566
=|2566,2567
=|2567,2568
=|2568,2569
<EOL>|2569,2570
ADMISSION|2570,2579
PHYSICAL|2580,2588
<EOL>|2588,2589
=|2589,2590
=|2590,2591
=|2591,2592
=|2592,2593
=|2593,2594
=|2594,2595
=|2595,2596
=|2596,2597
=|2597,2598
=|2598,2599
=|2599,2600
=|2600,2601
=|2601,2602
=|2602,2603
=|2603,2604
=|2604,2605
=|2605,2606
=|2606,2607
=|2607,2608
<EOL>|2608,2609
Vitals|2609,2615
:|2615,2616
98.9|2617,2621
_|2622,2623
_|2623,2624
_|2624,2625
74|2626,2628
18|2629,2631
96|2632,2634
%|2634,2635
RA|2636,2638
<EOL>|2640,2641
General|2641,2648
:|2648,2649
Alert|2650,2655
,|2655,2656
oriented|2657,2665
,|2665,2666
no|2667,2669
acute|2670,2675
distress|2676,2684
,|2684,2685
breathing|2686,2695
<EOL>|2696,2697
comfortably|2697,2708
<EOL>|2710,2711
HEENT|2711,2716
:|2716,2717
Sclera|2718,2724
anicteric|2725,2734
,|2734,2735
MMM|2736,2739
,|2739,2740
oropharynx|2741,2751
clear|2752,2757
,|2757,2758
EOMI|2759,2763
,|2763,2764
PERRL|2765,2770
<EOL>|2772,2773
Neck|2773,2777
:|2777,2778
Supple|2779,2785
,|2785,2786
JVP|2787,2790
not|2791,2794
elevated|2795,2803
,|2803,2804
no|2805,2807
LAD|2808,2811
<EOL>|2813,2814
CV|2814,2816
:|2816,2817
Regular|2818,2825
rate|2826,2830
and|2831,2834
rhythm|2835,2841
,|2841,2842
normal|2843,2849
S1|2850,2852
+|2853,2854
S2|2855,2857
,|2857,2858
no|2859,2861
murmurs|2862,2869
,|2869,2870
rubs|2871,2875
,|2875,2876
<EOL>|2877,2878
gallops|2878,2885
<EOL>|2887,2888
Lungs|2888,2893
:|2893,2894
Scattered|2895,2904
wheezes|2905,2912
throughout|2913,2923
,|2923,2924
bibasilar|2925,2934
crackles|2935,2943
,|2943,2944
<EOL>|2945,2946
moderate|2946,2954
air|2955,2958
movement|2959,2967
.|2967,2968
<EOL>|2970,2971
Abdomen|2971,2978
:|2978,2979
Soft|2980,2984
,|2984,2985
non-tender|2986,2996
,|2996,2997
non-distended|2998,3011
,|3011,3012
bowel|3013,3018
sounds|3019,3025
present|3026,3033
,|3033,3034
<EOL>|3035,3036
no|3036,3038
organomegaly|3039,3051
,|3051,3052
no|3053,3055
rebound|3056,3063
or|3064,3066
guarding|3067,3075
<EOL>|3077,3078
GU|3078,3080
:|3080,3081
No|3082,3084
foley|3085,3090
<EOL>|3092,3093
Ext|3093,3096
:|3096,3097
Warm|3098,3102
,|3102,3103
well|3104,3108
perfused|3109,3117
,|3117,3118
2|3119,3120
+|3120,3121
pulses|3122,3128
,|3128,3129
no|3130,3132
clubbing|3133,3141
,|3141,3142
cyanosis|3143,3151
or|3152,3154
<EOL>|3155,3156
edema|3156,3161
<EOL>|3163,3164
Neuro|3164,3169
:|3169,3170
Moves|3171,3176
all|3177,3180
extremities|3181,3192
well|3193,3197
<EOL>|3199,3200
<EOL>|3200,3201
=|3201,3202
=|3202,3203
=|3203,3204
=|3204,3205
=|3205,3206
=|3206,3207
=|3207,3208
=|3208,3209
=|3209,3210
=|3210,3211
=|3211,3212
=|3212,3213
=|3213,3214
=|3214,3215
=|3215,3216
=|3216,3217
=|3217,3218
=|3218,3219
<EOL>|3219,3220
DISCHARGE|3220,3229
PHYSICAL|3230,3238
<EOL>|3238,3239
=|3239,3240
=|3240,3241
=|3241,3242
=|3242,3243
=|3243,3244
=|3244,3245
=|3245,3246
=|3246,3247
=|3247,3248
=|3248,3249
=|3249,3250
=|3250,3251
=|3251,3252
=|3252,3253
=|3253,3254
=|3254,3255
=|3255,3256
=|3256,3257
<EOL>|3257,3258
Vitals|3258,3264
:|3264,3265
T|3266,3267
:|3267,3268
98.3|3269,3273
BP|3274,3276
:|3276,3277
149|3278,3281
/|3281,3282
87|3282,3284
P|3285,3286
:|3286,3287
83|3288,3290
R|3291,3292
:|3292,3293
18|3293,3295
O2|3296,3298
:|3298,3299
98|3300,3302
%|3302,3303
ra|3304,3306
<EOL>|3306,3307
General|3307,3314
:|3314,3315
NAD|3316,3319
<EOL>|3319,3320
Lungs|3320,3325
:|3325,3326
Diffuse|3327,3334
end|3335,3338
expiratory|3339,3349
wheezing|3350,3358
.|3358,3359
No|3360,3362
crackles|3363,3371
or|3372,3374
rhonchi|3375,3382
<EOL>|3382,3383
CV|3383,3385
:|3385,3386
RRR|3387,3390
.|3390,3391
no|3392,3394
M|3395,3396
/|3396,3397
R|3397,3398
/|3398,3399
G|3399,3400
<EOL>|3400,3401
Abdomen|3401,3408
:|3408,3409
NTND|3410,3414
<EOL>|3415,3416
Ext|3416,3419
:|3419,3420
No|3421,3423
edema|3424,3429
<EOL>|3430,3431
<EOL>|3432,3433
Pertinent|3433,3442
Results|3443,3450
:|3450,3451
<EOL>|3451,3452
=|3452,3453
=|3453,3454
=|3454,3455
=|3455,3456
=|3456,3457
=|3457,3458
=|3458,3459
=|3459,3460
=|3460,3461
=|3461,3462
=|3462,3463
=|3463,3464
=|3464,3465
=|3465,3466
=|3466,3467
=|3467,3468
=|3468,3469
=|3469,3470
=|3470,3471
=|3471,3472
=|3472,3473
<EOL>|3473,3474
ADMISSION|3474,3483
LABS|3484,3488
<EOL>|3488,3489
=|3489,3490
=|3490,3491
=|3491,3492
=|3492,3493
=|3493,3494
=|3494,3495
=|3495,3496
=|3496,3497
=|3497,3498
=|3498,3499
=|3499,3500
=|3500,3501
=|3501,3502
=|3502,3503
=|3503,3504
=|3504,3505
=|3505,3506
=|3506,3507
=|3507,3508
=|3508,3509
=|3509,3510
<EOL>|3510,3511
_|3511,3512
_|3512,3513
_|3513,3514
06|3515,3517
:|3517,3518
15PM|3518,3522
BLOOD|3523,3528
WBC|3529,3532
-|3532,3533
5.7|3533,3536
RBC|3537,3540
-|3540,3541
4|3541,3542
.|3542,3543
46|3543,3545
Hgb|3546,3549
-|3549,3550
12.9|3550,3554
Hct|3555,3558
-|3558,3559
40.2|3559,3563
MCV|3564,3567
-|3567,3568
90|3568,3570
<EOL>|3571,3572
MCH|3572,3575
-|3575,3576
28.9|3576,3580
MCHC|3581,3585
-|3585,3586
32.1|3586,3590
RDW|3591,3594
-|3594,3595
14.6|3595,3599
RDWSD|3600,3605
-|3605,3606
48|3606,3608
.|3608,3609
5|3609,3610
*|3610,3611
Plt|3612,3615
_|3616,3617
_|3617,3618
_|3618,3619
<EOL>|3619,3620
_|3620,3621
_|3621,3622
_|3622,3623
06|3624,3626
:|3626,3627
15PM|3627,3631
BLOOD|3632,3637
Neuts|3638,3643
-|3643,3644
62.1|3644,3648
_|3649,3650
_|3650,3651
_|3651,3652
Monos|3653,3658
-|3658,3659
9.4|3659,3662
Eos|3663,3666
-|3666,3667
0|3667,3668
.|3668,3669
3|3669,3670
*|3670,3671
<EOL>|3672,3673
Baso|3673,3677
-|3677,3678
0.3|3678,3681
Im|3682,3684
_|3685,3686
_|3686,3687
_|3687,3688
AbsNeut|3689,3696
-|3696,3697
3|3697,3698
.|3698,3699
55|3699,3701
AbsLymp|3702,3709
-|3709,3710
1|3710,3711
.|3711,3712
59|3712,3714
AbsMono|3715,3722
-|3722,3723
0|3723,3724
.|3724,3725
54|3725,3727
<EOL>|3728,3729
AbsEos|3729,3735
-|3735,3736
0|3736,3737
.|3737,3738
02|3738,3740
*|3740,3741
AbsBaso|3742,3749
-|3749,3750
0|3750,3751
.|3751,3752
02|3752,3754
<EOL>|3754,3755
_|3755,3756
_|3756,3757
_|3757,3758
06|3759,3761
:|3761,3762
15PM|3762,3766
BLOOD|3767,3772
Glucose|3773,3780
-|3780,3781
96|3781,3783
UreaN|3784,3789
-|3789,3790
15|3790,3792
Creat|3793,3798
-|3798,3799
0.9|3799,3802
Na|3803,3805
-|3805,3806
138|3806,3809
<EOL>|3810,3811
K|3811,3812
-|3812,3813
3.8|3813,3816
Cl|3817,3819
-|3819,3820
96|3820,3822
HCO3|3823,3827
-|3827,3828
32|3828,3830
AnGap|3831,3836
-|3836,3837
14|3837,3839
<EOL>|3839,3840
<EOL>|3840,3841
=|3841,3842
=|3842,3843
=|3843,3844
=|3844,3845
=|3845,3846
=|3846,3847
=|3847,3848
=|3848,3849
=|3849,3850
=|3850,3851
=|3851,3852
=|3852,3853
=|3853,3854
=|3854,3855
=|3855,3856
=|3856,3857
=|3857,3858
=|3858,3859
=|3859,3860
=|3860,3861
<EOL>|3861,3862
PERTINENT|3862,3871
LABS|3872,3876
<EOL>|3876,3877
=|3877,3878
=|3878,3879
=|3879,3880
=|3880,3881
=|3881,3882
=|3882,3883
=|3883,3884
=|3884,3885
=|3885,3886
=|3886,3887
=|3887,3888
=|3888,3889
=|3889,3890
=|3890,3891
=|3891,3892
=|3892,3893
=|3893,3894
=|3894,3895
=|3895,3896
=|3896,3897
<EOL>|3897,3898
_|3898,3899
_|3899,3900
_|3900,3901
05|3902,3904
:|3904,3905
55AM|3905,3909
BLOOD|3910,3915
cTropnT|3916,3923
-|3923,3924
<|3924,3925
0|3925,3926
.|3926,3927
01|3927,3929
<EOL>|3929,3930
_|3930,3931
_|3931,3932
_|3932,3933
12|3934,3936
:|3936,3937
16AM|3937,3941
BLOOD|3942,3947
cTropnT|3948,3955
-|3955,3956
<|3956,3957
0|3957,3958
.|3958,3959
01|3959,3961
<EOL>|3961,3962
_|3962,3963
_|3963,3964
_|3964,3965
06|3966,3968
:|3968,3969
15PM|3969,3973
BLOOD|3974,3979
cTropnT|3980,3987
-|3987,3988
<|3988,3989
0|3989,3990
.|3990,3991
01|3991,3993
<EOL>|3993,3994
<EOL>|3994,3995
=|3995,3996
=|3996,3997
=|3997,3998
=|3998,3999
=|3999,4000
=|4000,4001
=|4001,4002
=|4002,4003
=|4003,4004
=|4004,4005
=|4005,4006
=|4006,4007
=|4007,4008
=|4008,4009
=|4009,4010
=|4010,4011
=|4011,4012
=|4012,4013
=|4013,4014
=|4014,4015
<EOL>|4015,4016
DISCHARGE|4016,4025
LABS|4026,4030
<EOL>|4030,4031
=|4031,4032
=|4032,4033
=|4033,4034
=|4034,4035
=|4035,4036
=|4036,4037
=|4037,4038
=|4038,4039
=|4039,4040
=|4040,4041
=|4041,4042
=|4042,4043
=|4043,4044
=|4044,4045
=|4045,4046
=|4046,4047
=|4047,4048
=|4048,4049
=|4049,4050
=|4050,4051
<EOL>|4051,4052
_|4052,4053
_|4053,4054
_|4054,4055
05|4056,4058
:|4058,4059
55AM|4059,4063
BLOOD|4064,4069
WBC|4070,4073
-|4073,4074
4.8|4074,4077
RBC|4078,4081
-|4081,4082
4|4082,4083
.|4083,4084
13|4084,4086
Hgb|4087,4090
-|4090,4091
11.9|4091,4095
Hct|4096,4099
-|4099,4100
37.2|4100,4104
MCV|4105,4108
-|4108,4109
90|4109,4111
<EOL>|4112,4113
MCH|4113,4116
-|4116,4117
28.8|4117,4121
MCHC|4122,4126
-|4126,4127
32.0|4127,4131
RDW|4132,4135
-|4135,4136
14.6|4136,4140
RDWSD|4141,4146
-|4146,4147
47|4147,4149
.|4149,4150
8|4150,4151
*|4151,4152
Plt|4153,4156
_|4157,4158
_|4158,4159
_|4159,4160
<EOL>|4160,4161
_|4161,4162
_|4162,4163
_|4163,4164
05|4165,4167
:|4167,4168
55AM|4168,4172
BLOOD|4173,4178
_|4179,4180
_|4180,4181
_|4181,4182
PTT|4183,4186
-|4186,4187
29.0|4187,4191
_|4192,4193
_|4193,4194
_|4194,4195
<EOL>|4195,4196
_|4196,4197
_|4197,4198
_|4198,4199
05|4200,4202
:|4202,4203
55AM|4203,4207
BLOOD|4208,4213
Glucose|4214,4221
-|4221,4222
149|4222,4225
*|4225,4226
UreaN|4227,4232
-|4232,4233
17|4233,4235
Creat|4236,4241
-|4241,4242
0.8|4242,4245
Na|4246,4248
-|4248,4249
137|4249,4252
<EOL>|4253,4254
K|4254,4255
-|4255,4256
4.5|4256,4259
Cl|4260,4262
-|4262,4263
99|4263,4265
HCO3|4266,4270
-|4270,4271
29|4271,4273
AnGap|4274,4279
-|4279,4280
14|4280,4282
<EOL>|4282,4283
_|4283,4284
_|4284,4285
_|4285,4286
05|4287,4289
:|4289,4290
55AM|4290,4294
BLOOD|4295,4300
Calcium|4301,4308
-|4308,4309
9.6|4309,4312
Phos|4313,4317
-|4317,4318
2.9|4318,4321
Mg|4322,4324
-|4324,4325
2.0|4325,4328
<EOL>|4328,4329
<EOL>|4329,4330
=|4330,4331
=|4331,4332
=|4332,4333
=|4333,4334
=|4334,4335
=|4335,4336
=|4336,4337
=|4337,4338
=|4338,4339
=|4339,4340
=|4340,4341
=|4341,4342
=|4342,4343
=|4343,4344
=|4344,4345
=|4345,4346
=|4346,4347
=|4347,4348
=|4348,4349
=|4349,4350
<EOL>|4350,4351
EKG|4351,4354
<EOL>|4354,4355
=|4355,4356
=|4356,4357
=|4357,4358
=|4358,4359
=|4359,4360
=|4360,4361
=|4361,4362
=|4362,4363
=|4363,4364
=|4364,4365
=|4365,4366
=|4366,4367
=|4367,4368
=|4368,4369
=|4369,4370
=|4370,4371
=|4371,4372
=|4372,4373
=|4373,4374
=|4374,4375
<EOL>|4375,4376
_|4376,4377
_|4377,4378
_|4378,4379
<EOL>|4380,4381
Baseline|4381,4389
artifact|4390,4398
.|4398,4399
Probable|4400,4408
ectopic|4409,4416
atrial|4417,4423
rhythm|4424,4430
with|4431,4435
frequent|4436,4444
<EOL>|4445,4446
premature|4446,4455
<EOL>|4456,4457
atrial|4457,4463
contractions|4464,4476
.|4476,4477
Left|4478,4482
bundle|4483,4489
-|4489,4490
branch|4490,4496
block|4497,4502
.|4502,4503
Compared|4504,4512
to|4513,4515
the|4516,4519
<EOL>|4520,4521
previous|4521,4529
<EOL>|4530,4531
tracing|4531,4538
of|4539,4541
_|4542,4543
_|4543,4544
_|4544,4545
ectopic|4546,4553
atrial|4554,4560
rhythm|4561,4567
is|4568,4570
new|4571,4574
.|4574,4575
<EOL>|4576,4577
<EOL>|4577,4578
=|4578,4579
=|4579,4580
=|4580,4581
=|4581,4582
=|4582,4583
=|4583,4584
=|4584,4585
=|4585,4586
=|4586,4587
=|4587,4588
=|4588,4589
=|4589,4590
=|4590,4591
=|4591,4592
=|4592,4593
=|4593,4594
=|4594,4595
=|4595,4596
=|4596,4597
=|4597,4598
<EOL>|4598,4599
CXR|4599,4602
<EOL>|4602,4603
=|4603,4604
=|4604,4605
=|4605,4606
=|4606,4607
=|4607,4608
=|4608,4609
=|4609,4610
=|4610,4611
=|4611,4612
=|4612,4613
=|4613,4614
=|4614,4615
=|4615,4616
=|4616,4617
=|4617,4618
=|4618,4619
=|4619,4620
=|4620,4621
=|4621,4622
=|4622,4623
<EOL>|4623,4624
_|4624,4625
_|4625,4626
_|4626,4627
<EOL>|4627,4628
IMPRESSION|4628,4638
:|4638,4639
<EOL>|4639,4640
No|4640,4642
acute|4643,4648
cardiopulmonary|4649,4664
process|4665,4672
.|4672,4673
<EOL>|4673,4674
<EOL>|4675,4676
Brief|4676,4681
Hospital|4682,4690
Course|4691,4697
:|4697,4698
<EOL>|4698,4699
_|4699,4700
_|4700,4701
_|4701,4702
y|4703,4704
/|4704,4705
o|4705,4706
F|4707,4708
with|4709,4713
asthma|4714,4720
,|4720,4721
CAD|4722,4725
s|4726,4727
/|4727,4728
p|4728,4729
stents|4730,4736
(|4737,4738
reported|4738,4746
by|4747,4749
patient|4750,4757
)|4757,4758
,|4758,4759
<EOL>|4760,4761
COPD|4761,4765
,|4765,4766
PAD|4767,4770
,|4770,4771
HTN|4772,4775
,|4775,4776
who|4777,4780
presents|4781,4789
with|4790,4794
shortness|4795,4804
of|4805,4807
breath|4808,4814
and|4815,4818
<EOL>|4819,4820
intermittent|4820,4832
episode|4833,4840
of|4841,4843
chest|4844,4849
pain|4850,4854
.|4854,4855
<EOL>|4856,4857
<EOL>|4857,4858
#|4858,4859
Mild|4860,4864
COPD|4865,4869
exacerbation|4870,4882
:|4882,4883
Patient|4884,4891
with|4892,4896
shortness|4897,4906
of|4907,4909
breath|4910,4916
at|4917,4919
<EOL>|4920,4921
rest|4921,4925
,|4925,4926
no|4927,4929
cough|4930,4935
or|4936,4938
increased|4939,4948
sputum|4949,4955
production|4956,4966
.|4966,4967
Exam|4968,4972
with|4973,4977
wheezes|4978,4985
<EOL>|4986,4987
on|4987,4989
examination|4990,5001
and|5002,5005
some|5006,5010
improvement|5011,5022
with|5023,5027
nebs|5028,5032
/|5032,5033
pred|5033,5037
.|5037,5038
Lower|5039,5044
<EOL>|5045,5046
suspicion|5046,5055
for|5056,5059
PNA|5060,5063
given|5064,5069
normal|5070,5076
WBC|5077,5080
and|5081,5084
lack|5085,5089
of|5090,5092
fevers|5093,5099
.|5099,5100
Also|5101,5105
no|5106,5108
<EOL>|5109,5110
evidence|5110,5118
of|5119,5121
volume|5122,5128
overload|5129,5137
on|5138,5140
examination|5141,5152
.|5152,5153
Since|5154,5159
patient|5160,5167
only|5168,5172
<EOL>|5173,5174
has|5174,5177
a|5178,5179
mild|5180,5184
exacerbation|5185,5197
she|5198,5201
will|5202,5206
not|5207,5210
require|5211,5218
antibiotics|5219,5230
.|5230,5231
<EOL>|5232,5233
Paitent|5233,5240
will|5241,5245
recieve|5246,5253
5|5254,5255
days|5256,5260
of|5261,5263
predinose|5264,5273
(|5274,5275
last|5275,5279
day|5280,5283
_|5284,5285
_|5285,5286
_|5286,5287
in|5288,5290
<EOL>|5291,5292
addition|5292,5300
to|5301,5303
taking|5304,5310
her|5311,5314
home|5315,5319
albuterol|5320,5329
,|5329,5330
fluticasone|5331,5342
and|5343,5346
<EOL>|5347,5348
tiotropoium|5348,5359
inhalers|5360,5368
.|5368,5369
<EOL>|5369,5370
<EOL>|5370,5371
#|5371,5372
Episode|5373,5380
of|5381,5383
chest|5384,5389
pain|5390,5394
:|5394,5395
There|5396,5401
was|5402,5405
a|5406,5407
concern|5408,5415
for|5416,5419
ACS|5420,5423
given|5424,5429
<EOL>|5430,5431
cardiac|5431,5438
history|5439,5446
but|5447,5450
trops|5451,5456
x|5457,5458
2|5459,5460
negative|5461,5469
.|5469,5470
EKG|5471,5474
with|5475,5479
no|5480,5482
significant|5483,5494
<EOL>|5495,5496
changes|5496,5503
from|5504,5508
prior|5509,5514
.|5514,5515
The|5516,5519
chest|5520,5525
pain|5526,5530
was|5531,5534
non-exertional|5535,5549
,|5549,5550
resolved|5551,5559
<EOL>|5560,5561
without|5561,5568
intervention|5569,5581
prior|5582,5587
to|5588,5590
arriving|5591,5599
at|5600,5602
the|5603,5606
hospital|5607,5615
,|5615,5616
likely|5617,5623
<EOL>|5624,5625
related|5625,5632
to|5633,5635
her|5636,5639
COPD|5640,5644
exacerbation|5645,5657
.|5657,5658
<EOL>|5658,5659
<EOL>|5659,5660
TRANSITIONAL|5660,5672
ISSUES|5673,5679
:|5679,5680
<EOL>|5680,5681
[|5681,5682
]|5683,5684
Please|5685,5691
confirm|5692,5699
patient|5700,5707
completed|5708,5717
course|5718,5724
of|5725,5727
prednisone|5728,5738
(|5739,5740
last|5740,5744
<EOL>|5745,5746
day|5746,5749
_|5750,5751
_|5751,5752
_|5752,5753
with|5754,5758
resolution|5759,5769
of|5770,5772
symptoms|5773,5781
<EOL>|5781,5782
[|5782,5783
]|5784,5785
Consider|5786,5794
outpatient|5795,5805
stress|5806,5812
testing|5813,5820
if|5821,5823
chest|5824,5829
pain|5830,5834
returns|5835,5842
<EOL>|5842,5843
<EOL>|5844,5845
Medications|5845,5856
on|5857,5859
Admission|5860,5869
:|5869,5870
<EOL>|5870,5871
The|5871,5874
Preadmission|5875,5887
Medication|5888,5898
list|5899,5903
is|5904,5906
accurate|5907,5915
and|5916,5919
complete|5920,5928
.|5928,5929
<EOL>|5929,5930
1.|5930,5932
Acetaminophen|5933,5946
325|5947,5950
mg|5951,5953
PO|5954,5956
Q4H|5957,5960
:|5960,5961
PRN|5961,5964
pain|5965,5969
<EOL>|5970,5971
2.|5971,5973
Albuterol|5974,5983
0.083|5984,5989
%|5989,5990
Neb|5991,5994
Soln|5995,5999
1|6000,6001
NEB|6002,6005
IH|6006,6008
Q6H|6009,6012
:|6012,6013
PRN|6013,6016
shortness|6017,6026
of|6027,6029
<EOL>|6030,6031
breath|6031,6037
<EOL>|6038,6039
3.|6039,6041
Aspirin|6042,6049
81|6050,6052
mg|6053,6055
PO|6056,6058
DAILY|6059,6064
<EOL>|6065,6066
4.|6066,6068
Clopidogrel|6069,6080
75|6081,6083
mg|6084,6086
PO|6087,6089
DAILY|6090,6095
<EOL>|6096,6097
5.|6097,6099
Diltiazem|6100,6109
Extended|6110,6118
-|6118,6119
Release|6119,6126
180|6127,6130
mg|6131,6133
PO|6134,6136
DAILY|6137,6142
<EOL>|6143,6144
6.|6144,6146
Fluticasone|6147,6158
Propionate|6159,6169
NASAL|6170,6175
2|6176,6177
SPRY|6178,6182
NU|6183,6185
DAILY|6186,6191
:|6191,6192
PRN|6192,6195
nasal|6196,6201
<EOL>|6202,6203
congestion|6203,6213
<EOL>|6214,6215
7.|6215,6217
Hydrochlorothiazide|6218,6237
50|6238,6240
mg|6241,6243
PO|6244,6246
DAILY|6247,6252
<EOL>|6253,6254
8.|6254,6256
Isosorbide|6257,6267
Mononitrate|6268,6279
(|6280,6281
Extended|6281,6289
Release|6290,6297
)|6297,6298
120|6299,6302
mg|6303,6305
PO|6306,6308
DAILY|6309,6314
<EOL>|6315,6316
9.|6316,6318
Latanoprost|6319,6330
0.005|6331,6336
%|6336,6337
Ophth|6338,6343
.|6343,6344
Soln.|6345,6350
1|6351,6352
DROP|6353,6357
LEFT|6358,6362
EYE|6363,6366
HS|6367,6369
<EOL>|6370,6371
10.|6371,6374
Multivitamins|6375,6388
W|6389,6390
/|6390,6391
minerals|6391,6399
1|6400,6401
TAB|6402,6405
PO|6406,6408
DAILY|6409,6414
<EOL>|6415,6416
11.|6416,6419
Theophylline|6420,6432
ER|6433,6435
300|6436,6439
mg|6440,6442
PO|6443,6445
BID|6446,6449
<EOL>|6450,6451
12.|6451,6454
Tiotropium|6455,6465
Bromide|6466,6473
1|6474,6475
CAP|6476,6479
IH|6480,6482
DAILY|6483,6488
<EOL>|6489,6490
13.|6490,6493
Albuterol|6494,6503
Inhaler|6504,6511
2|6512,6513
PUFF|6514,6518
IH|6519,6521
Q4H|6522,6525
:|6525,6526
PRN|6526,6529
shortness|6530,6539
of|6540,6542
breath|6543,6549
<EOL>|6550,6551
14.|6551,6554
Calcarb|6555,6562
600|6563,6566
With|6567,6571
Vitamin|6572,6579
D|6580,6581
(|6582,6583
calcium|6583,6590
carbonate|6591,6600
-|6600,6601
vitamin|6601,6608
D3|6609,6611
)|6611,6612
<EOL>|6613,6614
315|6614,6617
/|6617,6618
200|6618,6621
mg|6622,6624
oral|6625,6629
daily|6630,6635
<EOL>|6636,6637
15.|6637,6640
cod|6641,6644
liver|6645,6650
oil|6651,6654
1,250|6655,6660
-|6660,6661
135|6661,6664
unit|6665,6669
oral|6670,6674
BID|6675,6678
<EOL>|6679,6680
16|6680,6682
.|6682,6683
Atorvastatin|6684,6696
10|6697,6699
mg|6700,6702
PO|6703,6705
QPM|6706,6709
<EOL>|6710,6711
17.|6711,6714
Fluticasone|6715,6726
-|6726,6727
Salmeterol|6727,6737
Diskus|6738,6744
(|6745,6746
250|6746,6749
/|6749,6750
50|6750,6752
)|6752,6753
1|6755,6756
INH|6757,6760
IH|6761,6763
BID|6764,6767
<EOL>|6768,6769
18.|6769,6772
Guaifenesin|6773,6784
-|6784,6785
CODEINE|6785,6792
Phosphate|6793,6802
5|6803,6804
mL|6805,6807
PO|6808,6810
Q6H|6811,6814
:|6814,6815
PRN|6815,6818
cough|6819,6824
<EOL>|6825,6826
19|6826,6828
.|6828,6829
TraMADOL|6830,6838
(|6839,6840
Ultram|6840,6846
)|6846,6847
50|6848,6850
mg|6851,6853
PO|6854,6856
Q6H|6857,6860
:|6860,6861
PRN|6861,6864
pain|6865,6869
<EOL>|6870,6871
20|6871,6873
.|6873,6874
Ranitidine|6875,6885
150|6886,6889
mg|6890,6892
PO|6893,6895
BID|6896,6899
<EOL>|6900,6901
21|6901,6903
.|6903,6904
Lorazepam|6905,6914
0.5|6915,6918
mg|6919,6921
PO|6922,6924
QHS|6925,6928
:|6928,6929
PRN|6929,6932
insomnia|6933,6941
<EOL>|6942,6943
<EOL>|6943,6944
<EOL>|6945,6946
Discharge|6946,6955
Medications|6956,6967
:|6967,6968
<EOL>|6968,6969
1.|6969,6971
Acetaminophen|6972,6985
325|6986,6989
mg|6990,6992
PO|6993,6995
Q4H|6996,6999
:|6999,7000
PRN|7000,7003
pain|7004,7008
<EOL>|7009,7010
2.|7010,7012
Albuterol|7013,7022
0.083|7023,7028
%|7028,7029
Neb|7030,7033
Soln|7034,7038
1|7039,7040
NEB|7041,7044
IH|7045,7047
Q6H|7048,7051
:|7051,7052
PRN|7052,7055
shortness|7056,7065
of|7066,7068
<EOL>|7069,7070
breath|7070,7076
<EOL>|7077,7078
3.|7078,7080
Aspirin|7081,7088
81|7089,7091
mg|7092,7094
PO|7095,7097
DAILY|7098,7103
<EOL>|7104,7105
4.|7105,7107
Atorvastatin|7108,7120
10|7121,7123
mg|7124,7126
PO|7127,7129
QPM|7130,7133
<EOL>|7134,7135
5.|7135,7137
Clopidogrel|7138,7149
75|7150,7152
mg|7153,7155
PO|7156,7158
DAILY|7159,7164
<EOL>|7165,7166
6.|7166,7168
Diltiazem|7169,7178
Extended|7179,7187
-|7187,7188
Release|7188,7195
180|7196,7199
mg|7200,7202
PO|7203,7205
DAILY|7206,7211
<EOL>|7212,7213
7.|7213,7215
Fluticasone|7216,7227
Propionate|7228,7238
NASAL|7239,7244
2|7245,7246
SPRY|7247,7251
NU|7252,7254
DAILY|7255,7260
:|7260,7261
PRN|7261,7264
nasal|7265,7270
<EOL>|7271,7272
congestion|7272,7282
<EOL>|7283,7284
8.|7284,7286
Fluticasone|7287,7298
-|7298,7299
Salmeterol|7299,7309
Diskus|7310,7316
(|7317,7318
250|7318,7321
/|7321,7322
50|7322,7324
)|7324,7325
1|7327,7328
INH|7329,7332
IH|7333,7335
BID|7336,7339
<EOL>|7340,7341
9.|7341,7343
Hydrochlorothiazide|7344,7363
50|7364,7366
mg|7367,7369
PO|7370,7372
DAILY|7373,7378
<EOL>|7379,7380
10.|7380,7383
Isosorbide|7384,7394
Mononitrate|7395,7406
(|7407,7408
Extended|7408,7416
Release|7417,7424
)|7424,7425
120|7426,7429
mg|7430,7432
PO|7433,7435
DAILY|7436,7441
<EOL>|7442,7443
11.|7443,7446
Latanoprost|7447,7458
0.005|7459,7464
%|7464,7465
Ophth|7466,7471
.|7471,7472
Soln.|7473,7478
1|7479,7480
DROP|7481,7485
LEFT|7486,7490
EYE|7491,7494
HS|7495,7497
<EOL>|7498,7499
12.|7499,7502
Lorazepam|7503,7512
0.5|7513,7516
mg|7517,7519
PO|7520,7522
QHS|7523,7526
:|7526,7527
PRN|7527,7530
insomnia|7531,7539
<EOL>|7540,7541
13.|7541,7544
Multivitamins|7545,7558
W|7559,7560
/|7560,7561
minerals|7561,7569
1|7570,7571
TAB|7572,7575
PO|7576,7578
DAILY|7579,7584
<EOL>|7585,7586
14.|7586,7589
Ranitidine|7590,7600
150|7601,7604
mg|7605,7607
PO|7608,7610
BID|7611,7614
<EOL>|7615,7616
15.|7616,7619
TraMADOL|7620,7628
(|7629,7630
Ultram|7630,7636
)|7636,7637
50|7638,7640
mg|7641,7643
PO|7644,7646
Q6H|7647,7650
:|7650,7651
PRN|7651,7654
pain|7655,7659
<EOL>|7660,7661
16|7661,7663
.|7663,7664
PredniSONE|7665,7675
40|7676,7678
mg|7679,7681
PO|7682,7684
DAILY|7685,7690
Duration|7691,7699
:|7699,7700
4|7701,7702
Days|7703,7707
<EOL>|7708,7709
RX|7709,7711
*|7712,7713
prednisone|7713,7723
20|7724,7726
mg|7727,7729
2|7730,7731
tablet|7732,7738
(|7738,7739
s|7739,7740
)|7740,7741
by|7742,7744
mouth|7745,7750
once|7751,7755
a|7756,7757
day|7758,7761
Disp|7762,7766
#|7767,7768
*|7768,7769
6|7769,7770
<EOL>|7771,7772
Tablet|7772,7778
Refills|7779,7786
:|7786,7787
*|7787,7788
0|7788,7789
<EOL>|7789,7790
17.|7790,7793
Theophylline|7794,7806
ER|7807,7809
300|7810,7813
mg|7814,7816
PO|7817,7819
BID|7820,7823
<EOL>|7824,7825
18.|7825,7828
Tiotropium|7829,7839
Bromide|7840,7847
1|7848,7849
CAP|7850,7853
IH|7854,7856
DAILY|7857,7862
<EOL>|7863,7864
19|7864,7866
.|7866,7867
Guaifenesin|7868,7879
-|7879,7880
CODEINE|7880,7887
Phosphate|7888,7897
5|7898,7899
mL|7900,7902
PO|7903,7905
Q6H|7906,7909
:|7909,7910
PRN|7910,7913
cough|7914,7919
<EOL>|7920,7921
20|7921,7923
.|7923,7924
cod|7925,7928
liver|7929,7934
oil|7935,7938
1,250|7939,7944
-|7944,7945
135|7945,7948
unit|7949,7953
oral|7954,7958
BID|7959,7962
<EOL>|7963,7964
21|7964,7966
.|7966,7967
Calcarb|7968,7975
600|7976,7979
With|7980,7984
Vitamin|7985,7992
D|7993,7994
(|7995,7996
calcium|7996,8003
carbonate|8004,8013
-|8013,8014
vitamin|8014,8021
D3|8022,8024
)|8024,8025
<EOL>|8026,8027
315|8027,8030
/|8030,8031
200|8031,8034
mg|8035,8037
oral|8038,8042
daily|8043,8048
<EOL>|8049,8050
<EOL>|8050,8051
<EOL>|8052,8053
Discharge|8053,8062
Disposition|8063,8074
:|8074,8075
<EOL>|8075,8076
Home|8076,8080
<EOL>|8080,8081
<EOL>|8082,8083
Discharge|8083,8092
Diagnosis|8093,8102
:|8102,8103
<EOL>|8103,8104
Primary|8104,8111
Diagnosis|8112,8121
:|8121,8122
<EOL>|8122,8123
COPD|8123,8127
exacerbation|8128,8140
<EOL>|8140,8141
<EOL>|8141,8142
<EOL>|8143,8144
Discharge|8144,8153
Condition|8154,8163
:|8163,8164
<EOL>|8164,8165
Mental|8165,8171
Status|8172,8178
:|8178,8179
Clear|8180,8185
and|8186,8189
coherent|8190,8198
.|8198,8199
<EOL>|8199,8200
Level|8200,8205
of|8206,8208
Consciousness|8209,8222
:|8222,8223
Alert|8224,8229
and|8230,8233
interactive|8234,8245
.|8245,8246
<EOL>|8246,8247
Activity|8247,8255
Status|8256,8262
:|8262,8263
Ambulatory|8264,8274
-|8275,8276
Independent|8277,8288
.|8288,8289
<EOL>|8289,8290
<EOL>|8290,8291
<EOL>|8292,8293
Discharge|8293,8302
Instructions|8303,8315
:|8315,8316
<EOL>|8316,8317
Dear|8317,8321
Ms.|8322,8325
_|8326,8327
_|8327,8328
_|8328,8329
,|8329,8330
<EOL>|8330,8331
<EOL>|8331,8332
You|8332,8335
were|8336,8340
admitted|8341,8349
to|8350,8352
the|8353,8356
hospital|8357,8365
for|8366,8369
shortness|8370,8379
of|8380,8382
breath|8383,8389
and|8390,8393
<EOL>|8394,8395
mild|8395,8399
chest|8400,8405
pain|8406,8410
.|8410,8411
While|8412,8417
in|8418,8420
the|8421,8424
hospital|8425,8433
we|8434,8436
received|8437,8445
an|8446,8448
EKG|8449,8452
and|8453,8456
<EOL>|8457,8458
blood|8458,8463
work|8464,8468
which|8469,8474
suggested|8475,8484
that|8485,8489
your|8490,8494
pain|8495,8499
was|8500,8503
not|8504,8507
coming|8508,8514
from|8515,8519
<EOL>|8520,8521
your|8521,8525
heart|8526,8531
.|8531,8532
Your|8533,8537
shortness|8538,8547
of|8548,8550
breath|8551,8557
is|8558,8560
likely|8561,8567
from|8568,8572
a|8573,8574
COPD|8575,8579
<EOL>|8580,8581
attack|8581,8587
and|8588,8591
we|8592,8594
gave|8595,8599
you|8600,8603
steroids|8604,8612
and|8613,8616
breathing|8617,8626
treatments|8627,8637
for|8638,8641
<EOL>|8642,8643
your|8643,8647
symptoms|8648,8656
.|8656,8657
<EOL>|8658,8659
<EOL>|8659,8660
You|8660,8663
have|8664,8668
a|8669,8670
follow|8671,8677
up|8678,8680
appointment|8681,8692
with|8693,8697
Dr.|8698,8701
_|8702,8703
_|8703,8704
_|8704,8705
as|8706,8708
detailed|8709,8717
<EOL>|8718,8719
below|8719,8724
.|8724,8725
We|8726,8728
are|8729,8732
also|8733,8737
sending|8738,8745
you|8746,8749
home|8750,8754
with|8755,8759
a|8760,8761
short|8762,8767
course|8768,8774
of|8775,8777
<EOL>|8778,8779
steroids|8779,8787
for|8788,8791
your|8792,8796
COPD|8797,8801
.|8801,8802
Your|8803,8807
other|8808,8813
medications|8814,8825
are|8826,8829
detailed|8830,8838
in|8839,8841
<EOL>|8842,8843
your|8843,8847
discharge|8848,8857
medication|8858,8868
list|8869,8873
.|8873,8874
<EOL>|8874,8875
<EOL>|8875,8876
It|8876,8878
was|8879,8882
a|8883,8884
pleasure|8885,8893
taking|8894,8900
care|8901,8905
of|8906,8908
you|8909,8912
at|8913,8915
_|8916,8917
_|8917,8918
_|8918,8919
.|8919,8920
<EOL>|8920,8921
<EOL>|8921,8922
Sincerely|8922,8931
,|8931,8932
<EOL>|8932,8933
Your|8933,8937
_|8938,8939
_|8939,8940
_|8940,8941
Care|8942,8946
Team|8947,8951
<EOL>|8951,8952
<EOL>|8953,8954
Followup|8954,8962
Instructions|8963,8975
:|8975,8976
<EOL>|8976,8977
_|8977,8978
_|8978,8979
_|8979,8980
<EOL>|8980,8981

