 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Procedure|Health Care Activity|SIMPLE_SEGMENT|46,55|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|46,60|false|false|false|C2598112||Admission Date
Finding|Body Substance|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|80,89|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|80,94|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|136,139|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|147,154|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|147,154|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|156,164|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Drug|Amino Acid, Peptide, or Protein|Allergies|179,189|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|Allergies|179,189|false|false|false|C0065374|lisinopril|lisinopril
Finding|Functional Concept|Allergies|192,201|false|false|false|C1999232|Attending (action)|Attending
Anatomy|Body Location or Region|Chief Complaint|227,232|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|Chief Complaint|227,232|false|false|false|C0741025|Chest problem|Chest
Attribute|Clinical Attribute|Chief Complaint|227,237|false|false|false|C2926613||Chest Pain
Finding|Sign or Symptom|Chief Complaint|227,237|false|false|false|C0008031|Chest Pain|Chest Pain
Attribute|Clinical Attribute|Chief Complaint|233,237|false|true|false|C2598155||Pain
Finding|Functional Concept|Chief Complaint|233,237|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Chief Complaint|233,237|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Classification|Chief Complaint|240,245|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|246,254|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|246,254|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|258,276|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|267,276|false|false|false|C0945766||Procedure
Event|Occupational Activity|Chief Complaint|267,276|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|267,276|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|267,276|false|false|false|C0184661|Interventional procedure|Procedure
Finding|Daily or Recreational Activity|Chief Complaint|278,286|false|false|false|C0015259|Exercise|Exercise
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|278,286|false|false|false|C1522704|Exercise Pain Management|Exercise
Procedure|Diagnostic Procedure|Chief Complaint|287,303|false|false|false|C0013516;C2729489|Echocardiography;echocardiography service|Echocardiography
Procedure|Health Care Activity|Chief Complaint|287,303|false|false|false|C0013516;C2729489|Echocardiography;echocardiography service|Echocardiography
Finding|Finding|History of Present Illness|339,342|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|pmh
Finding|Finding|History of Present Illness|343,349|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|History of Present Illness|343,349|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|History of Present Illness|356,359|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|356,359|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|History of Present Illness|356,359|false|false|false|C1504769|DFFB protein, human|CAD
Finding|Gene or Genome|History of Present Illness|356,359|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|History of Present Illness|356,359|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|History of Present Illness|356,359|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|356,359|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|364,368|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Finding|Intellectual Product|History of Present Illness|394,401|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|History of Present Illness|394,401|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Event|Occupational Activity|History of Present Illness|411,418|false|false|false|C1273870|Management procedure|managed
Attribute|Clinical Attribute|History of Present Illness|419,425|false|false|false|C2926611||angina
Finding|Finding|History of Present Illness|419,425|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Finding|Sign or Symptom|History of Present Illness|419,425|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Disorder|Disease or Syndrome|History of Present Illness|432,435|false|false|false|C0020538|Hypertensive disease|HTN
Finding|Finding|History of Present Illness|459,467|false|false|false|C0741302|atypia morphology|atypical
Finding|Sign or Symptom|History of Present Illness|459,478|false|false|false|C0262384|Atypical chest pain|atypical chest pain
Anatomy|Body Location or Region|History of Present Illness|468,473|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|468,473|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|468,478|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|468,478|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|474,478|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|474,478|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|474,478|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Body Substance|History of Present Illness|486,493|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|486,493|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|486,493|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Functional Concept|History of Present Illness|486,497|false|false|false|C0332310|Has patient|Patient has
Finding|Conceptual Entity|History of Present Illness|498,505|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|498,505|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|498,505|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|498,508|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|History of Present Illness|509,512|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|509,512|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|History of Present Illness|509,512|false|false|false|C1504769|DFFB protein, human|CAD
Finding|Gene or Genome|History of Present Illness|509,512|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|History of Present Illness|509,512|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|History of Present Illness|509,512|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|509,512|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Anatomy|Body Location or Region|History of Present Illness|526,532|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|526,532|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|533,537|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|544,547|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|History of Present Illness|544,547|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|History of Present Illness|544,547|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Disorder|Disease or Syndrome|History of Present Illness|619,625|false|false|false|C4255010||NSTEMI
Finding|Finding|History of Present Illness|619,625|false|false|false|C3537184||NSTEMI
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|634,638|false|false|false|C0007430|Catheterization|cath
Finding|Finding|History of Present Illness|653,661|false|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Finding|Functional Concept|History of Present Illness|653,661|false|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Anatomy|Tissue|History of Present Illness|662,667|false|false|false|C0332835|Transplanted tissue|graft
Drug|Biomedical or Dental Material|History of Present Illness|662,667|false|false|false|C0181074;C1705210|Graft Dosage Form;Graft material|graft
Finding|Intellectual Product|History of Present Illness|662,667|false|false|false|C1546653|Graft - Specimen Source Codes|graft
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|662,667|false|false|false|C1961139;C3683798|Graft Procedures on the Head;Grafting procedure|graft
Drug|Chemical Viewed Structurally|History of Present Illness|688,694|false|false|false|C1881507|Macromolecular Branch|branch
Finding|Finding|History of Present Illness|699,703|false|false|false|C5575035|Well (answer to question)|well
Finding|Pathologic Function|History of Present Illness|714,722|false|false|false|C1261287|Stenosis|stenosis
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|730,733|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|History of Present Illness|730,733|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|History of Present Illness|730,733|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Finding|Pathologic Function|History of Present Illness|753,761|false|false|false|C1261287|Stenosis|stenosis
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|769,772|false|false|false|C2987138|Methylcytosine Dioxygenase TET1|LCx
Drug|Enzyme|History of Present Illness|769,772|false|false|false|C2987138|Methylcytosine Dioxygenase TET1|LCx
Finding|Gene or Genome|History of Present Illness|769,772|false|false|false|C1428863;C2987137|TET1 gene;TET1 wt Allele|LCx
Finding|Classification|History of Present Illness|774,780|false|false|false|C0079946;C1550512|National origin;Participation Type - origin|origin
Finding|Intellectual Product|History of Present Illness|774,780|false|false|false|C0079946;C1550512|National origin;Participation Type - origin|origin
Drug|Organic Chemical|History of Present Illness|840,845|false|false|false|C0590690|Imdur|Imdur
Drug|Pharmacologic Substance|History of Present Illness|840,845|false|false|false|C0590690|Imdur|Imdur
Finding|Functional Concept|History of Present Illness|850,860|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Finding|Genetic Function|History of Present Illness|850,860|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Finding|Mental Process|History of Present Illness|850,860|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Drug|Organic Chemical|History of Present Illness|864,872|false|false|false|C0126174|losartan|losartan
Drug|Pharmacologic Substance|History of Present Illness|864,872|false|false|false|C0126174|losartan|losartan
Finding|Idea or Concept|History of Present Illness|877,883|false|false|false|C1550462|Observation Interpretation - better|better
Drug|Organic Chemical|History of Present Illness|887,894|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|History of Present Illness|887,894|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|History of Present Illness|887,894|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Finding|Conceptual Entity|History of Present Illness|887,894|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|History of Present Illness|887,894|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|History of Present Illness|887,894|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Intellectual Product|History of Present Illness|901,906|false|false|false|C4050225|Often - answer to question|often
Attribute|Clinical Attribute|History of Present Illness|911,917|false|false|false|C2926611||angina
Finding|Finding|History of Present Illness|911,917|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Finding|Sign or Symptom|History of Present Illness|911,917|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Disorder|Disease or Syndrome|History of Present Illness|911,925|false|false|false|C0002965;C0152172|Angina decubitus;Angina, Unstable|angina at rest
Finding|Functional Concept|History of Present Illness|918,925|false|false|false|C0443144|At rest (qualifier value)|at rest
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|921,925|false|false|false|C1742913|REST protein, human|rest
Drug|Biologically Active Substance|History of Present Illness|921,925|false|false|false|C1742913|REST protein, human|rest
Finding|Daily or Recreational Activity|History of Present Illness|921,925|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Gene or Genome|History of Present Illness|921,925|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Molecular Function|History of Present Illness|921,925|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Drug|Biomedical or Dental Material|History of Present Illness|944,952|false|false|false|C0168634|BaseLine dental cement|baseline
Finding|Idea or Concept|History of Present Illness|944,952|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Drug|Organic Chemical|History of Present Illness|960,973|false|false|false|C0017887|nitroglycerin|nitroglycerin
Drug|Pharmacologic Substance|History of Present Illness|960,973|false|false|false|C0017887|nitroglycerin|nitroglycerin
Anatomy|Body Location or Region|History of Present Illness|1047,1052|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|1047,1052|false|false|false|C0741025|Chest problem|chest
Finding|Sign or Symptom|History of Present Illness|1047,1058|false|false|false|C0008031|Chest Pain|chest pains
Finding|Sign or Symptom|History of Present Illness|1053,1058|false|false|false|C0030193|Pain|pains
Finding|Intellectual Product|History of Present Illness|1089,1096|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|History of Present Illness|1089,1096|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Attribute|Clinical Attribute|History of Present Illness|1097,1103|false|false|false|C2926611||angina
Finding|Finding|History of Present Illness|1097,1103|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Finding|Sign or Symptom|History of Present Illness|1097,1103|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Finding|Finding|History of Present Illness|1111,1118|false|false|false|C3888388|Usually|usually
Anatomy|Body Location or Region|History of Present Illness|1123,1128|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|1123,1128|false|false|false|C0741025|Chest problem|chest
Finding|Intellectual Product|History of Present Illness|1170,1176|false|false|false|C1546717||needle
Disorder|Injury or Poisoning|History of Present Illness|1177,1183|false|false|false|C0033119|Puncture wound|pricks
Finding|Finding|History of Present Illness|1177,1183|false|false|false|C0439821|Pricking sensation quality|pricks
Attribute|Clinical Attribute|History of Present Illness|1186,1190|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|1186,1190|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1186,1190|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Idea or Concept|History of Present Illness|1238,1249|false|true|false|C0750502|Significant|significant
Drug|Organic Chemical|History of Present Illness|1250,1256|true|true|false|C0723011|Relief brand of phenylephrine|relief
Drug|Pharmacologic Substance|History of Present Illness|1250,1256|true|true|false|C0723011|Relief brand of phenylephrine|relief
Finding|Finding|History of Present Illness|1250,1256|true|true|false|C0564405|Feeling relief|relief
Finding|Finding|History of Present Illness|1281,1286|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Idea or Concept|History of Present Illness|1281,1286|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Attribute|Clinical Attribute|History of Present Illness|1292,1296|false|false|false|C4318566|Deep Resection Margin|deep
Finding|Finding|History of Present Illness|1292,1306|false|false|false|C1321587;C1328799|Breathing abnormally deep;Deep breathing|deep breathing
Finding|Sign or Symptom|History of Present Illness|1292,1306|false|false|false|C1321587;C1328799|Breathing abnormally deep;Deep breathing|deep breathing
Attribute|Clinical Attribute|History of Present Illness|1297,1306|false|false|false|C5885990||breathing
Finding|Finding|History of Present Illness|1297,1306|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|History of Present Illness|1297,1306|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|History of Present Illness|1297,1306|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|History of Present Illness|1297,1306|false|false|false|C1160636|respiratory system process|breathing
Finding|Finding|History of Present Illness|1317,1325|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|History of Present Illness|1317,1325|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|History of Present Illness|1317,1325|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|History of Present Illness|1317,1325|false|false|false|C0033095||pressure
Disorder|Disease or Syndrome|History of Present Illness|1329,1337|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Anatomy|Body Location or Region|History of Present Illness|1329,1343|false|false|false|C0230132|Anterior chest wall structure|anterior chest
Anatomy|Body Location or Region|History of Present Illness|1338,1343|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|1338,1343|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|1383,1387|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|1383,1387|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1383,1387|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1407,1411|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Attribute|Clinical Attribute|History of Present Illness|1419,1423|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|1419,1423|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1419,1423|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1484,1487|false|false|false|C0013404|Dyspnea|SOB
Finding|Finding|History of Present Illness|1492,1503|false|true|false|C0700590|Increased sweating|diaphoresis
Attribute|Clinical Attribute|History of Present Illness|1522,1528|false|false|false|C4255480||nausea
Finding|Sign or Symptom|History of Present Illness|1522,1528|false|false|false|C0027497|Nausea|nausea
Finding|Finding|History of Present Illness|1535,1547|false|false|false|C0030252|Palpitations|palpitations
Finding|Finding|History of Present Illness|1582,1589|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|History of Present Illness|1582,1589|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Finding|History of Present Illness|1591,1600|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Finding|Sign or Symptom|History of Present Illness|1591,1600|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Anatomy|Body Location or Region|History of Present Illness|1602,1607|false|false|false|C0003086;C0003087;C4284979|Ankle;Ankle joint structure;Lower extremity>Ankle|ankle
Anatomy|Body Space or Junction|History of Present Illness|1602,1607|false|false|false|C0003086;C0003087;C4284979|Ankle;Ankle joint structure;Lower extremity>Ankle|ankle
Finding|Pathologic Function|History of Present Illness|1602,1613|false|false|false|C0235439|Ankle edema (finding)|ankle edema
Attribute|Clinical Attribute|History of Present Illness|1608,1613|false|false|false|C1717255||edema
Finding|Pathologic Function|History of Present Illness|1608,1613|false|false|false|C0013604|Edema|edema
Finding|Finding|History of Present Illness|1615,1627|false|false|false|C0030252|Palpitations|palpitations
Finding|Sign or Symptom|History of Present Illness|1629,1636|false|false|false|C0039070|Syncope|syncope
Finding|Sign or Symptom|History of Present Illness|1641,1651|false|false|false|C0700200|Presyncope|presyncope
Disorder|Disease or Syndrome|History of Present Illness|1699,1703|false|false|false|C0009443;C0024117|Chronic Obstructive Airway Disease;Common Cold|cold
Drug|Organic Chemical|History of Present Illness|1699,1703|false|false|false|C0719425|Cold brand of chlorpheniramine-phenylpropanolamine|cold
Drug|Pharmacologic Substance|History of Present Illness|1699,1703|false|false|false|C0719425|Cold brand of chlorpheniramine-phenylpropanolamine|cold
Finding|Organism Function|History of Present Illness|1699,1703|false|false|false|C0234192|Cold Sensation|cold
Phenomenon|Natural Phenomenon or Process|History of Present Illness|1699,1703|false|false|false|C0009264|Cold Temperature|cold
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1699,1703|false|false|false|C0010412|Cold Therapy|cold
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1725,1728|false|false|false|C0028723;C2985261|NUT Family Member 1, human;Nuts|nut
Drug|Biologically Active Substance|History of Present Illness|1725,1728|false|false|false|C0028723;C2985261|NUT Family Member 1, human;Nuts|nut
Drug|Food|History of Present Illness|1725,1728|false|false|false|C0028723;C2985261|NUT Family Member 1, human;Nuts|nut
Finding|Gene or Genome|History of Present Illness|1725,1728|false|false|false|C1837033;C2985260|NUTM1 gene;NUTM1 wt Allele|nut
Finding|Sign or Symptom|History of Present Illness|1740,1746|true|false|false|C0015967|Fever|fevers
Finding|Sign or Symptom|History of Present Illness|1750,1756|true|false|false|C0085593|Chills|chills
Finding|Intellectual Product|History of Present Illness|1768,1775|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|History of Present Illness|1768,1775|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Drug|Organic Chemical|History of Present Illness|1788,1793|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|1788,1793|false|false|false|C3815497|Cough (guaifenesin)|cough
Finding|Sign or Symptom|History of Present Illness|1788,1793|false|false|false|C0010200|Coughing|cough
Finding|Finding|History of Present Illness|1817,1827|false|false|false|C5441521|Complaint (finding)|complaints
Finding|Body Substance|History of Present Illness|1843,1850|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1843,1850|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1843,1850|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|History of Present Illness|1887,1891|false|false|false|C5890125|Loss (adaptation)|loss
Finding|Functional Concept|History of Present Illness|1897,1906|false|false|false|C1516691|Cognitive|cognitive
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|1897,1917|false|false|false|C0338656|Impaired cognition|cognitive impairment
Finding|Finding|History of Present Illness|1907,1917|false|false|false|C0221099;C0684336|Impaired;Impaired health|impairment
Finding|Functional Concept|History of Present Illness|1907,1917|false|false|false|C0221099;C0684336|Impaired;Impaired health|impairment
Finding|Intellectual Product|History of Present Illness|1972,1975|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|History of Present Illness|1972,1975|false|false|false|C1623258|Electrocardiography|EKG
Anatomy|Body Space or Junction|History of Present Illness|1977,1982|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|History of Present Illness|1977,1982|false|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|History of Present Illness|1977,1982|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|History of Present Illness|1977,1982|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|1997,2008|false|false|false|C0011570|Mental Depression|depressions
Finding|Finding|History of Present Illness|2030,2033|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|History of Present Illness|2030,2033|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Functional Concept|History of Present Illness|2035,2043|false|false|false|C0475224|Ischemic|ischemic
Lab|Laboratory or Test Result|History of Present Illness|2050,2054|false|false|false|C0587081|Laboratory test finding|Labs
Finding|Finding|History of Present Illness|2074,2077|false|false|false|C5848551|Neg - answer|neg
Procedure|Diagnostic Procedure|History of Present Illness|2082,2085|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Intellectual Product|History of Present Illness|2090,2095|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2126,2133|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|Past Medical History|2126,2133|false|false|false|C1314974|Cardiac attachment|CARDIAC
Finding|Finding|Past Medical History|2126,2138|false|false|false|C3176821|CARD.RISK|CARDIAC RISK
Finding|Finding|Past Medical History|2126,2146|false|false|false|C2024776|cardiac risk factors|CARDIAC RISK FACTORS
Finding|Idea or Concept|Past Medical History|2134,2138|false|false|false|C0035647|Risk|RISK
Attribute|Clinical Attribute|Past Medical History|2134,2146|false|false|false|C1830376||RISK FACTORS
Finding|Finding|Past Medical History|2134,2146|false|false|false|C0035648;C0455624;C1553898|History of - risk factor;risk factors;risk factors - observation list|RISK FACTORS
Finding|Intellectual Product|Past Medical History|2134,2146|false|false|false|C0035648;C0455624;C1553898|History of - risk factor;risk factors;risk factors - observation list|RISK FACTORS
Disorder|Disease or Syndrome|Past Medical History|2151,2159|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|Diabetes
Disorder|Disease or Syndrome|Past Medical History|2164,2176|false|false|false|C0242339|Dyslipidemias|Dyslipidemia
Disorder|Disease or Syndrome|Past Medical History|2181,2184|false|false|false|C0020538|Hypertensive disease|HTN
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2190,2197|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|Past Medical History|2190,2197|false|false|false|C1314974|Cardiac attachment|CARDIAC
Anatomy|Body Part, Organ, or Organ Component|Patient History|2210,2218|false|false|false|C0018787|Heart|Coronary
Anatomy|Body Part, Organ, or Organ Component|Patient History|2210,2225|false|false|false|C0205042|Coronary artery|Coronary artery
Disorder|Disease or Syndrome|Patient History|2210,2233|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|Coronary artery disease
Anatomy|Body Part, Organ, or Organ Component|Patient History|2219,2225|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|Patient History|2219,2225|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Disorder|Disease or Syndrome|Patient History|2219,2233|false|false|false|C0852949|Arteriopathic disease|artery disease
Disorder|Disease or Syndrome|Patient History|2226,2233|false|false|false|C0012634|Disease|disease
Attribute|Clinical Attribute|Patient History|2237,2246|false|false|false|C0012000|Diastole|Diastolic
Disorder|Disease or Syndrome|Patient History|2237,2271|false|false|false|C2183328|diastolic congestive heart failure|Diastolic congestive heart failure
Disorder|Disease or Syndrome|Patient History|2247,2271|false|false|false|C0018802|Congestive heart failure|congestive heart failure
Anatomy|Body Part, Organ, or Organ Component|Patient History|2258,2263|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Patient History|2258,2263|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Patient History|2258,2263|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|Patient History|2258,2271|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Finding|Functional Concept|Patient History|2264,2271|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|Patient History|2264,2271|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|Patient History|2264,2271|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Procedure|Therapeutic or Preventive Procedure|Patient History|2275,2279|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Procedure|Therapeutic or Preventive Procedure|Patient History|2281,2285|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Procedure|Therapeutic or Preventive Procedure|Patient History|2291,2322|false|false|false|C1449706|Coronary Artery Bypass, Off-Pump|Off pump coronary artery bypass
Finding|Molecular Function|Patient History|2295,2299|false|false|false|C1150186|matrix metalloproteinase 7 activity|pump
Anatomy|Body Part, Organ, or Organ Component|Patient History|2300,2308|false|false|false|C0018787|Heart|coronary
Anatomy|Body Part, Organ, or Organ Component|Patient History|2300,2315|false|false|false|C0205042|Coronary artery|coronary artery
Procedure|Therapeutic or Preventive Procedure|Patient History|2300,2322|false|false|false|C0010055|Coronary Artery Bypass Surgery|coronary artery bypass
Procedure|Therapeutic or Preventive Procedure|Patient History|2300,2328|false|false|false|C0010055|Coronary Artery Bypass Surgery|coronary artery bypass graft
Anatomy|Body Part, Organ, or Organ Component|Patient History|2309,2315|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|Patient History|2309,2315|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Procedure|Therapeutic or Preventive Procedure|Patient History|2309,2328|false|false|false|C5886769|Arterial bypass graft|artery bypass graft
Procedure|Therapeutic or Preventive Procedure|Patient History|2316,2322|false|false|false|C0813207|Creation of shunt|bypass
Procedure|Therapeutic or Preventive Procedure|Patient History|2316,2328|false|false|false|C0185098|Bypass graft|bypass graft
Anatomy|Tissue|Patient History|2323,2328|false|false|false|C0332835|Transplanted tissue|graft
Drug|Biomedical or Dental Material|Patient History|2323,2328|false|false|false|C0181074;C1705210|Graft Dosage Form;Graft material|graft
Finding|Intellectual Product|Patient History|2323,2328|false|false|false|C1546653|Graft - Specimen Source Codes|graft
Procedure|Therapeutic or Preventive Procedure|Patient History|2323,2328|false|false|false|C1961139;C3683798|Graft Procedures on the Head;Grafting procedure|graft
Finding|Functional Concept|Patient History|2333,2337|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Patient History|2341,2364|false|false|false|C0226276|Structure of internal thoracic artery|internal mammary artery
Anatomy|Body Part, Organ, or Organ Component|Patient History|2350,2357|false|false|false|C0006141;C0929301|Breast;Mammary gland|mammary
Anatomy|Body Part, Organ, or Organ Component|Patient History|2350,2364|false|false|false|C0024661|Mammary Arteries|mammary artery
Anatomy|Body Part, Organ, or Organ Component|Patient History|2358,2364|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|Patient History|2358,2364|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Finding|Functional Concept|Patient History|2368,2372|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Patient History|2368,2399|false|false|false|C0226032;C1321506|Anterior descending branch of left coronary artery|left anterior descending artery
Disorder|Disease or Syndrome|Patient History|2373,2381|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Finding|Functional Concept|Patient History|2382,2392|false|false|false|C1547177|Sequencing - Descending|descending
Anatomy|Body Part, Organ, or Organ Component|Patient History|2393,2399|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|Patient History|2393,2399|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body Part, Organ, or Organ Component|Patient History|2406,2420|false|false|false|C0036186;C0392907|Great saphenous vein structure;Saphenous Vein|saphenous vein
Anatomy|Body Part, Organ, or Organ Component|Patient History|2416,2420|false|false|false|C0042449|Veins|vein
Anatomy|Tissue|Patient History|2421,2427|false|false|false|C0332835|Transplanted tissue|grafts
Drug|Biomedical or Dental Material|Patient History|2421,2427|false|false|false|C0181074|Graft material|grafts
Finding|Finding|Patient History|2452,2460|false|false|false|C1550517|Target Awareness - marginal|marginal
Anatomy|Body Part, Organ, or Organ Component|Patient History|2461,2469|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Anatomy|Body System|Patient History|2461,2469|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Procedure|Health Care Activity|Patient History|2461,2469|false|false|false|C0397581|Procedure on artery|arteries
Finding|Functional Concept|Patient History|2475,2487|false|false|false|C1522243|Percutaneous Route of Drug Administration|PERCUTANEOUS
Procedure|Therapeutic or Preventive Procedure|Patient History|2475,2510|false|false|false|C1532338|Percutaneous Coronary Intervention|PERCUTANEOUS CORONARY INTERVENTIONS
Anatomy|Body Part, Organ, or Organ Component|Patient History|2488,2496|false|false|false|C0018787|Heart|CORONARY
Attribute|Clinical Attribute|Patient History|2497,2510|false|false|false|C2979881||INTERVENTIONS
Procedure|Health Care Activity|Patient History|2497,2510|false|false|false|C0886296;C1273869|Intervention regimes;Nursing interventions|INTERVENTIONS
Disorder|Disease or Syndrome|Patient History|2512,2515|false|false|false|C0006430|Burning Mouth Syndrome|BMS
Attribute|Clinical Attribute|Patient History|2519,2527|false|false|false|C4489236|Proximal Resection Margin|proximal
Anatomy|Body Part, Organ, or Organ Component|Patient History|2528,2531|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|Patient History|2528,2531|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|Patient History|2528,2531|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Disorder|Disease or Syndrome|Patient History|2539,2542|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|Patient History|2539,2542|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|Patient History|2539,2542|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|Patient History|2539,2542|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|Patient History|2539,2542|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|Patient History|2539,2542|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Finding|Gene or Genome|Patient History|2539,2542|false|false|false|C1413980|DES gene|DES
Anatomy|Body Part, Organ, or Organ Component|Patient History|2550,2553|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|Patient History|2550,2553|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|Patient History|2550,2553|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Disorder|Disease or Syndrome|Patient History|2559,2562|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|Patient History|2559,2562|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|Patient History|2559,2562|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|Patient History|2559,2562|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|Patient History|2559,2562|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|Patient History|2559,2562|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Finding|Gene or Genome|Patient History|2559,2562|false|false|false|C1413980|DES gene|DES
Finding|Conceptual Entity|Patient History|2566,2570|false|false|false|C2697523|Graph Edge|edge
Anatomy|Body Part, Organ, or Organ Component|Patient History|2582,2585|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|Patient History|2582,2585|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|Patient History|2582,2585|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Disorder|Disease or Syndrome|Patient History|2586,2589|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|Patient History|2586,2589|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|Patient History|2586,2589|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|Patient History|2586,2589|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|Patient History|2586,2589|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|Patient History|2586,2589|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Finding|Gene or Genome|Patient History|2586,2589|false|false|false|C1413980|DES gene|DES
Finding|Pathologic Function|Patient History|2596,2604|false|false|false|C1261287|Stenosis|stenosis
Attribute|Clinical Attribute|Patient History|2605,2611|false|false|false|C4522154|Distal Resection Margin|distal
Disorder|Disease or Syndrome|Patient History|2626,2629|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|Patient History|2626,2629|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|Patient History|2626,2629|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|Patient History|2626,2629|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|Patient History|2626,2629|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|Patient History|2626,2629|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Finding|Gene or Genome|Patient History|2626,2629|false|false|false|C1413980|DES gene|DES
Finding|Individual Behavior|Patient History|2645,2651|false|false|false|C0562458|Pacing up and down|PACING
Disorder|Disease or Syndrome|Patient History|2652,2655|false|false|false|C0020725;C0021122|Disruptive, Impulse Control, and Conduct Disorders;Type II Mucolipidosis|ICD
Disorder|Mental or Behavioral Dysfunction|Patient History|2652,2655|false|false|false|C0020725;C0021122|Disruptive, Impulse Control, and Conduct Disorders;Type II Mucolipidosis|ICD
Finding|Gene or Genome|Patient History|2652,2655|false|false|false|C0870733;C5891008|GNPTAB wt Allele;International Classification of Diseases|ICD
Finding|Intellectual Product|Patient History|2652,2655|false|false|false|C0870733;C5891008|GNPTAB wt Allele;International Classification of Diseases|ICD
Procedure|Therapeutic or Preventive Procedure|Patient History|2652,2655|false|false|false|C5575277|Icd Regimen|ICD
Disorder|Disease or Syndrome|Patient History|2663,2677|false|false|false|C0028756|Morbid obesity|Morbid obesity
Disorder|Disease or Syndrome|Patient History|2670,2677|false|false|false|C0028754|Obesity|obesity
Finding|Finding|Patient History|2670,2677|false|false|false|C4759928|BODY MASS INDEX QUANTITATIVE TRAIT LOCUS 20|obesity
Disorder|Disease or Syndrome|Patient History|2681,2685|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Patient History|2681,2685|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|Patient History|2681,2685|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|Patient History|2688,2692|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Finding|Functional Concept|Patient History|2695,2700|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Location or Region|Patient History|2695,2713|false|false|false|C0828608|Right tendinous cuff|Right rotator cuff
Anatomy|Body Part, Organ, or Organ Component|Patient History|2701,2713|false|false|false|C0085515|Rotator Cuff|rotator cuff
Disorder|Injury or Poisoning|Patient History|2701,2720|false|false|false|C0851122|Rotator Cuff Injuries|rotator cuff injury
Anatomy|Body Part, Organ, or Organ Component|Patient History|2709,2713|false|false|false|C1550244|Cuff - body part|cuff
Finding|Pathologic Function|Patient History|2709,2713|false|false|false|C3668885|Cuffing (morphologic abnormality)|cuff
Disorder|Injury or Poisoning|Patient History|2714,2720|false|false|false|C3263722;C3263723|Traumatic AND/OR non-traumatic injury;Traumatic injury|injury
Disorder|Disease or Syndrome|Patient History|2721,2729|false|false|false|C0006444|Bursitis|bursitis
Disorder|Disease or Syndrome|Patient History|2732,2741|false|false|false|C0149931|Migraine Disorders|Migraines
Disorder|Mental or Behavioral Dysfunction|Patient History|2744,2754|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|Depression
Finding|Functional Concept|Patient History|2744,2754|false|false|false|C0460137;C1579931|Depression - motion|Depression
Finding|Sign or Symptom|Patient History|2744,2754|false|false|false|C0460137;C1579931|Depression - motion|Depression
Disorder|Disease or Syndrome|Patient History|2757,2760|false|false|false|C0029408|Degenerative polyarthritis|DJD
Disorder|Disease or Syndrome|Patient History|2763,2774|false|false|false|C0019112|Hemorrhoids|Hemorrhoids
Disorder|Disease or Syndrome|Patient History|2777,2784|false|false|false|C0035854|Rosacea|Rosacea
Drug|Amino Acid, Peptide, or Protein|Family Medical History|2870,2880|false|true|false|C3812393|ErbB Receptors|her family
Drug|Enzyme|Family Medical History|2870,2880|false|true|false|C3812393|ErbB Receptors|her family
Finding|Receptor|Family Medical History|2870,2880|false|true|false|C3812393|ErbB Receptors|her family
Finding|Classification|Family Medical History|2874,2880|true|true|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Family Medical History|2874,2880|true|true|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Family Medical History|2874,2880|true|true|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Family Medical History|2874,2880|true|true|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Procedure|Health Care Activity|General Exam|2902,2911|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Finding|Functional Concept|General Exam|2912,2916|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|2912,2916|false|false|false|C0582103|Medical Examination|EXAM
Finding|Classification|General Exam|2965,2972|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|General Exam|2965,2972|false|false|false|C3812897|General medical service|GENERAL
Finding|Finding|General Exam|2974,2982|false|false|false|C1961028|Oriented to place|Oriented
Attribute|Clinical Attribute|General Exam|2987,2991|false|false|false|C2713234||Mood
Finding|Conceptual Entity|General Exam|2987,2991|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Finding|Finding|General Exam|2987,2991|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Finding|Mental Process|General Exam|2987,2991|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Anatomy|Body Location or Region|General Exam|3015,3020|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|General Exam|3028,3034|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|General Exam|3028,3034|false|false|false|C0036412|Scleral Diseases|Sclera
Procedure|Health Care Activity|General Exam|3028,3034|false|false|false|C2228481|examination of sclera|Sclera
Finding|Finding|General Exam|3035,3044|false|false|false|C0205180|Anicteric|anicteric
Finding|Finding|General Exam|3046,3051|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Anatomy|Body Part, Organ, or Organ Component|General Exam|3059,3070|false|false|false|C0009758;C0229274|Structure of palpebral conjunctiva;conjunctiva|Conjunctiva
Disorder|Disease or Syndrome|General Exam|3059,3070|false|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|Conjunctiva
Disorder|Neoplastic Process|General Exam|3059,3070|false|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|Conjunctiva
Finding|Body Substance|General Exam|3059,3070|false|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|Conjunctiva
Finding|Intellectual Product|General Exam|3059,3070|false|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|Conjunctiva
Procedure|Health Care Activity|General Exam|3059,3070|false|false|false|C0872390;C2228431|Procedure on conjunctiva;examination of conjunctiva|Conjunctiva
Finding|Finding|General Exam|3086,3092|true|false|false|C0241137|Pallor of skin|pallor
Finding|Sign or Symptom|General Exam|3096,3104|true|false|false|C0010520|Cyanosis|cyanosis
Anatomy|Body Space or Junction|General Exam|3112,3116|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|General Exam|3112,3116|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|General Exam|3112,3116|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|General Exam|3112,3116|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Anatomy|Body Part, Organ, or Organ Component|General Exam|3112,3123|false|false|false|C0026639|Oral mucous membrane structure|oral mucosa
Anatomy|Tissue|General Exam|3117,3123|false|false|false|C0026724|Mucous Membrane|mucosa
Finding|Intellectual Product|General Exam|3117,3123|false|false|false|C1561514||mucosa
Disorder|Disease or Syndrome|General Exam|3128,3139|true|false|false|C0155210;C0302314|Eyelid Xanthoma;Xanthoma|xanthelasma
Anatomy|Body Location or Region|General Exam|3144,3148|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|General Exam|3144,3148|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|General Exam|3144,3148|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Finding|Functional Concept|General Exam|3150,3156|false|false|false|C0332254|Supple|Supple
Finding|Finding|General Exam|3162,3165|false|false|false|C0428897|Jugular venous pressure|JVP
Anatomy|Body Location or Region|General Exam|3177,3182|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|General Exam|3177,3182|false|false|false|C0741025|Chest problem|Chest
Finding|Idea or Concept|General Exam|3184,3195|false|false|false|C0750502|Significant|significant
Disorder|Disease or Syndrome|General Exam|3204,3207|false|false|false|C0034155;C1268935|Congenital Thrombotic Thrombocytopenic Purpura;Purpura, Thrombotic Thrombocytopenic|TTP
Drug|Amino Acid, Peptide, or Protein|General Exam|3204,3207|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Drug|Biologically Active Substance|General Exam|3204,3207|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Drug|Organic Chemical|General Exam|3204,3207|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Drug|Vitamin|General Exam|3204,3207|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Finding|Gene or Genome|General Exam|3204,3207|false|false|false|C1413036;C1421571;C3539814|ADAMTS13 gene;ZFP36 gene;ZFP36 wt Allele|TTP
Disorder|Disease or Syndrome|General Exam|3213,3221|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Anatomy|Body Location or Region|General Exam|3213,3227|false|false|false|C0230132|Anterior chest wall structure|anterior chest
Anatomy|Body Location or Region|General Exam|3213,3232|false|false|false|C0230132;C1305714|Anterior chest wall structure|anterior chest wall
Anatomy|Body Part, Organ, or Organ Component|General Exam|3213,3232|false|false|false|C0230132;C1305714|Anterior chest wall structure|anterior chest wall
Anatomy|Body Location or Region|General Exam|3222,3227|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|General Exam|3222,3227|false|false|false|C0741025|Chest problem|chest
Anatomy|Body Location or Region|General Exam|3222,3232|false|false|false|C0205076;C4266615|Chest wall structure;Chest>Chest wall|chest wall
Anatomy|Body Part, Organ, or Organ Component|General Exam|3222,3232|false|false|false|C0205076;C4266615|Chest wall structure;Chest>Chest wall|chest wall
Anatomy|Body Part, Organ, or Organ Component|General Exam|3236,3243|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|General Exam|3236,3243|false|false|false|C1314974|Cardiac attachment|CARDIAC
Procedure|Therapeutic or Preventive Procedure|General Exam|3249,3253|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Finding|Finding|General Exam|3271,3278|true|false|false|C0232269|Cardiac thrill (finding)|thrills
Anatomy|Body Part, Organ, or Organ Component|General Exam|3303,3308|false|false|false|C0024109|Lung|LUNGS
Finding|Functional Concept|General Exam|3317,3321|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Finding|General Exam|3330,3338|false|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Finding|Idea or Concept|General Exam|3352,3362|false|true|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|General Exam|3352,3367|false|true|false|C0332290|Consistent with|consistent with
Anatomy|Tissue|General Exam|3369,3376|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|General Exam|3369,3376|false|false|false|C0032226|Pleural Diseases|pleural
Anatomy|Body Part, Organ, or Organ Component|General Exam|3377,3384|false|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|General Exam|3377,3384|false|false|false|C1951340|Process Pharmacologic Substance|process
Finding|Functional Concept|General Exam|3377,3384|false|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|General Exam|3377,3384|false|false|false|C1522240|Process|process
Procedure|Diagnostic Procedure|General Exam|3393,3396|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Idea or Concept|General Exam|3408,3412|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Drug|Inorganic Chemical|General Exam|3413,3416|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|General Exam|3413,3416|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|General Exam|3413,3416|false|false|false|C0001861;C3536832|Air (substance);air|air
Finding|Finding|General Exam|3413,3416|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|General Exam|3413,3416|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|General Exam|3413,3416|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Phenomenon|Natural Phenomenon or Process|General Exam|3413,3425|false|false|false|C0001868|Air Movements|air movement
Finding|Organism Function|General Exam|3417,3425|false|false|false|C0026649|Movement|movement
Finding|Sign or Symptom|General Exam|3435,3442|false|false|false|C0043144|Wheezing|wheezes
Finding|Finding|General Exam|3446,3453|false|false|false|C0035508|Rhonchi|rhonchi
Anatomy|Body Location or Region|General Exam|3457,3464|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|General Exam|3457,3464|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Finding|Finding|General Exam|3457,3464|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|General Exam|3466,3470|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Finding|Gene or Genome|General Exam|3481,3484|true|false|false|C1537594|LRRC4B gene|HSM
Finding|Mental Process|General Exam|3488,3498|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|General Exam|3488,3498|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Anatomy|Body Location or Region|General Exam|3500,3503|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|Abd
Disorder|Cell or Molecular Dysfunction|General Exam|3500,3503|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|Abd
Anatomy|Body Part, Organ, or Organ Component|General Exam|3504,3509|false|false|false|C0003483;C4037978|Aorta;Chest+Abdomen>Aorta|aorta
Procedure|Health Care Activity|General Exam|3504,3509|false|false|false|C0869784|Procedure on aorta|aorta
Procedure|Diagnostic Procedure|General Exam|3527,3536|false|false|false|C0030247|Palpation|palpation
Anatomy|Body Location or Region|General Exam|3541,3550|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|General Exam|3541,3557|true|false|false|C0221755|Abdominal bruit|abdominal bruits
Finding|Finding|General Exam|3551,3557|true|false|false|C0006318|Bruit|bruits
Anatomy|Body Part, Organ, or Organ Component|General Exam|3561,3572|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Anatomy|Body Part, Organ, or Organ Component|General Exam|3587,3594|false|false|false|C0015811|Femur|femoral
Finding|Finding|General Exam|3595,3601|true|false|false|C0006318|Bruit|bruits
Anatomy|Body System|General Exam|3605,3609|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|General Exam|3605,3609|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|General Exam|3605,3609|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Finding|Body Substance|General Exam|3605,3609|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|General Exam|3605,3609|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Pathologic Function|General Exam|3614,3620|false|false|false|C0333138|Stasis|stasis
Disorder|Disease or Syndrome|General Exam|3614,3631|true|false|false|C0011620|Stasis dermatitis|stasis dermatitis
Disorder|Disease or Syndrome|General Exam|3621,3631|true|false|false|C0011603|Dermatitis|dermatitis
Finding|Pathologic Function|General Exam|3633,3639|true|false|false|C0041582|Ulcer|ulcers
Finding|Finding|General Exam|3641,3646|true|false|false|C0241158;C2004491|Cicatrix;Scar Tissue|scars
Finding|Pathologic Function|General Exam|3641,3646|true|false|false|C0241158;C2004491|Cicatrix;Scar Tissue|scars
Disorder|Disease or Syndrome|General Exam|3651,3660|true|false|false|C0302314|Xanthoma|xanthomas
Drug|Food|General Exam|3664,3670|false|false|false|C5890763||PULSES
Finding|Physiologic Function|General Exam|3664,3670|false|false|false|C0391850|Physiologic pulse|PULSES
Procedure|Health Care Activity|General Exam|3664,3670|false|false|false|C0034107|Pulse taking|PULSES
Finding|Body Substance|General Exam|3722,3731|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|3722,3731|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|3722,3731|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|3722,3731|false|false|false|C0030685|Patient Discharge|DISCHARGE
Finding|Functional Concept|General Exam|3732,3736|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|3732,3736|false|false|false|C0582103|Medical Examination|EXAM
Finding|Classification|General Exam|3790,3797|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|General Exam|3790,3797|false|false|false|C3812897|General medical service|GENERAL
Finding|Finding|General Exam|3799,3807|false|false|false|C1961028|Oriented to place|Oriented
Attribute|Clinical Attribute|General Exam|3812,3816|false|false|false|C2713234||Mood
Finding|Conceptual Entity|General Exam|3812,3816|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Finding|Finding|General Exam|3812,3816|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Finding|Mental Process|General Exam|3812,3816|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Finding|Finding|General Exam|3834,3845|false|false|false|C0233471|Flat affect|flat affect
Finding|Mental Process|General Exam|3839,3845|false|false|false|C0001721|Affect (mental function)|affect
Procedure|Health Care Activity|General Exam|3839,3845|false|false|false|C2237113|assessment of affect|affect
Disorder|Disease or Syndrome|General Exam|3848,3851|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|3848,3851|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|3848,3851|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|3848,3851|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|3848,3851|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Finding|Finding|General Exam|3848,3851|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|General Exam|3854,3859|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|General Exam|3867,3873|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|General Exam|3867,3873|false|false|false|C0036412|Scleral Diseases|Sclera
Procedure|Health Care Activity|General Exam|3867,3873|false|false|false|C2228481|examination of sclera|Sclera
Finding|Finding|General Exam|3874,3883|false|false|false|C0205180|Anicteric|anicteric
Finding|Finding|General Exam|3885,3890|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Anatomy|Body Part, Organ, or Organ Component|General Exam|3898,3909|false|false|false|C0009758;C0229274|Structure of palpebral conjunctiva;conjunctiva|Conjunctiva
Disorder|Disease or Syndrome|General Exam|3898,3909|false|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|Conjunctiva
Disorder|Neoplastic Process|General Exam|3898,3909|false|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|Conjunctiva
Finding|Body Substance|General Exam|3898,3909|false|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|Conjunctiva
Finding|Intellectual Product|General Exam|3898,3909|false|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|Conjunctiva
Procedure|Health Care Activity|General Exam|3898,3909|false|false|false|C0872390;C2228431|Procedure on conjunctiva;examination of conjunctiva|Conjunctiva
Finding|Finding|General Exam|3925,3931|true|false|false|C0241137|Pallor of skin|pallor
Finding|Sign or Symptom|General Exam|3935,3943|true|false|false|C0010520|Cyanosis|cyanosis
Anatomy|Body Space or Junction|General Exam|3951,3955|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|General Exam|3951,3955|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|General Exam|3951,3955|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|General Exam|3951,3955|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Anatomy|Body Part, Organ, or Organ Component|General Exam|3951,3962|false|false|false|C0026639|Oral mucous membrane structure|oral mucosa
Anatomy|Tissue|General Exam|3956,3962|false|false|false|C0026724|Mucous Membrane|mucosa
Finding|Intellectual Product|General Exam|3956,3962|false|false|false|C1561514||mucosa
Disorder|Disease or Syndrome|General Exam|3967,3978|true|false|false|C0155210;C0302314|Eyelid Xanthoma;Xanthoma|xanthelasma
Finding|Functional Concept|General Exam|3982,3986|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|General Exam|3982,3993|false|false|false|C0229124|Structure of cornea of left eye|Left cornea
Anatomy|Body Part, Organ, or Organ Component|General Exam|3987,3993|false|false|false|C0010031|Cornea|cornea
Disorder|Disease or Syndrome|General Exam|3987,3993|false|false|false|C0010034;C0153629;C0154026|Benign neoplasm of cornea;Corneal Diseases;Malignant neoplasm of cornea|cornea
Disorder|Neoplastic Process|General Exam|3987,3993|false|false|false|C0010034;C0153629;C0154026|Benign neoplasm of cornea;Corneal Diseases;Malignant neoplasm of cornea|cornea
Finding|Body Substance|General Exam|3987,3993|false|false|false|C1550625|SpecimenType - Cornea|cornea
Finding|Finding|General Exam|3999,4003|false|false|false|C0241158;C1419736;C2004491|Cicatrix;RPS4X gene;Scar Tissue|scar
Finding|Gene or Genome|General Exam|3999,4003|false|false|false|C0241158;C1419736;C2004491|Cicatrix;RPS4X gene;Scar Tissue|scar
Finding|Pathologic Function|General Exam|3999,4003|false|false|false|C0241158;C1419736;C2004491|Cicatrix;RPS4X gene;Scar Tissue|scar
Finding|Finding|General Exam|3999,4010|false|false|false|C0241158;C2004491|Cicatrix;Scar Tissue|scar tissue
Finding|Pathologic Function|General Exam|3999,4010|false|false|false|C0241158;C2004491|Cicatrix;Scar Tissue|scar tissue
Anatomy|Tissue|General Exam|4004,4010|false|false|false|C0040300|Body tissue|tissue
Finding|Intellectual Product|General Exam|4004,4010|false|false|false|C1547928|Tissue Specimen Code|tissue
Anatomy|Body Location or Region|General Exam|4026,4030|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|General Exam|4026,4030|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|General Exam|4026,4030|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Finding|Functional Concept|General Exam|4032,4038|false|false|false|C0332254|Supple|Supple
Finding|Finding|General Exam|4049,4052|false|false|false|C0428897|Jugular venous pressure|JVP
Disorder|Disease or Syndrome|General Exam|4058,4069|true|false|false|C0018021|Goiter|thyromegaly
Anatomy|Body Location or Region|General Exam|4071,4076|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|CHEST
Finding|Finding|General Exam|4071,4076|false|false|false|C0741025|Chest problem|CHEST
Disorder|Disease or Syndrome|General Exam|4078,4081|false|false|false|C0034155;C1268935|Congenital Thrombotic Thrombocytopenic Purpura;Purpura, Thrombotic Thrombocytopenic|TTP
Drug|Amino Acid, Peptide, or Protein|General Exam|4078,4081|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Drug|Biologically Active Substance|General Exam|4078,4081|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Drug|Organic Chemical|General Exam|4078,4081|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Drug|Vitamin|General Exam|4078,4081|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Finding|Gene or Genome|General Exam|4078,4081|false|false|false|C1413036;C1421571;C3539814|ADAMTS13 gene;ZFP36 gene;ZFP36 wt Allele|TTP
Anatomy|Body Part, Organ, or Organ Component|General Exam|4087,4094|false|false|false|C0038293|Sternum|sternum
Anatomy|Body Part, Organ, or Organ Component|General Exam|4095,4102|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|General Exam|4095,4102|false|false|false|C1314974|Cardiac attachment|CARDIAC
Finding|Pathologic Function|General Exam|4104,4111|false|false|false|C5441917|Distant Metastasis|Distant
Finding|Finding|General Exam|4104,4124|false|false|false|C2198873|distant heart sounds|Distant heart sounds
Anatomy|Body Part, Organ, or Organ Component|General Exam|4112,4117|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|General Exam|4112,4117|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|General Exam|4112,4117|false|false|false|C0795691|HEART PROBLEM|heart
Attribute|Clinical Attribute|General Exam|4112,4124|false|false|false|C4050434||heart sounds
Finding|Organ or Tissue Function|General Exam|4112,4124|false|false|false|C0018820|Heart Sounds|heart sounds
Procedure|Diagnostic Procedure|General Exam|4112,4124|false|false|false|C2230284|auscultation of heart sounds|heart sounds
Phenomenon|Natural Phenomenon or Process|General Exam|4118,4124|false|false|false|C0037709||sounds
Finding|Finding|General Exam|4139,4146|true|false|false|C0232269|Cardiac thrill (finding)|thrills
Anatomy|Body Part, Organ, or Organ Component|General Exam|4171,4176|false|false|false|C0024109|Lung|LUNGS
Drug|Organic Chemical|General Exam|4178,4182|false|false|false|C0951233|cetrimonium bromide|CTAB
Finding|Sign or Symptom|General Exam|4186,4194|true|false|false|C0043144|Wheezing|wheezing
Finding|Finding|General Exam|4196,4201|true|false|false|C0034642;C0240859|Basilar Rales;Rales|rales
Finding|Finding|General Exam|4203,4210|true|false|false|C0035508|Rhonchi|rhonchi
Anatomy|Body Location or Region|General Exam|4213,4220|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|General Exam|4213,4220|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Finding|Finding|General Exam|4213,4220|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|General Exam|4222,4227|false|false|false|C0028754|Obesity|Obese
Disorder|Disease or Syndrome|General Exam|4229,4233|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Finding|Gene or Genome|General Exam|4244,4247|true|false|false|C1537594|LRRC4B gene|HSM
Finding|Mental Process|General Exam|4251,4261|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|General Exam|4251,4261|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Anatomy|Body Location or Region|General Exam|4263,4266|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|Abd
Disorder|Cell or Molecular Dysfunction|General Exam|4263,4266|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|Abd
Anatomy|Body Part, Organ, or Organ Component|General Exam|4267,4272|false|false|false|C0003483;C4037978|Aorta;Chest+Abdomen>Aorta|aorta
Procedure|Health Care Activity|General Exam|4267,4272|false|false|false|C0869784|Procedure on aorta|aorta
Procedure|Diagnostic Procedure|General Exam|4290,4299|false|false|false|C0030247|Palpation|palpation
Anatomy|Body Location or Region|General Exam|4304,4313|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|General Exam|4304,4320|true|false|false|C0221755|Abdominal bruit|abdominal bruits
Finding|Finding|General Exam|4314,4320|true|false|false|C0006318|Bruit|bruits
Anatomy|Body Part, Organ, or Organ Component|General Exam|4324,4335|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Anatomy|Body Part, Organ, or Organ Component|General Exam|4350,4357|false|false|false|C0015811|Femur|femoral
Finding|Finding|General Exam|4358,4364|true|false|false|C0006318|Bruit|bruits
Anatomy|Body System|General Exam|4368,4372|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|General Exam|4368,4372|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|General Exam|4368,4372|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Finding|Body Substance|General Exam|4368,4372|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|General Exam|4368,4372|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Pathologic Function|General Exam|4377,4383|false|false|false|C0333138|Stasis|stasis
Disorder|Disease or Syndrome|General Exam|4377,4394|true|false|false|C0011620|Stasis dermatitis|stasis dermatitis
Disorder|Disease or Syndrome|General Exam|4384,4394|true|false|false|C0011603|Dermatitis|dermatitis
Finding|Pathologic Function|General Exam|4396,4402|true|false|false|C0041582|Ulcer|ulcers
Finding|Finding|General Exam|4404,4409|true|false|false|C0241158;C2004491|Cicatrix;Scar Tissue|scars
Finding|Pathologic Function|General Exam|4404,4409|true|false|false|C0241158;C2004491|Cicatrix;Scar Tissue|scars
Disorder|Disease or Syndrome|General Exam|4414,4423|true|false|false|C0302314|Xanthoma|xanthomas
Drug|Food|General Exam|4427,4433|false|false|false|C5890763||PULSES
Finding|Physiologic Function|General Exam|4427,4433|false|false|false|C0391850|Physiologic pulse|PULSES
Procedure|Health Care Activity|General Exam|4427,4433|false|false|false|C0034107|Pulse taking|PULSES
Finding|Conceptual Entity|General Exam|4438,4444|false|false|false|C0442038;C0920847|Circumpennate;Radial|radial
Finding|Gene or Genome|General Exam|4445,4448|false|false|false|C1414174;C5848994|DSPP gene;DSPP wt Allele|DPP
Finding|Functional Concept|General Exam|4472,4476|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|General Exam|4472,4476|false|false|false|C0582103|Medical Examination|exam
Procedure|Health Care Activity|General Exam|4499,4508|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Lab|Laboratory or Test Result|General Exam|4509,4513|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|General Exam|4528,4533|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4528,4533|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|4534,4537|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|4542,4545|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|4542,4545|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|4542,4545|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|4552,4555|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|4552,4555|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|4552,4555|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|4552,4555|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|4561,4564|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|4561,4564|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|4571,4574|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|General Exam|4571,4574|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|4571,4574|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|4571,4574|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|4578,4581|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|4578,4581|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|General Exam|4578,4581|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|4578,4581|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|4578,4581|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|4588,4592|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|4607,4610|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|4627,4632|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4627,4632|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|4637,4640|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Procedure|Laboratory Procedure|General Exam|4637,4640|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|General Exam|4662,4667|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4662,4667|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|4662,4675|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|4662,4675|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|4662,4675|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|4668,4675|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|4668,4675|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|4668,4675|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|General Exam|4668,4675|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|4668,4675|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|4721,4725|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|4721,4725|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|4721,4725|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|4750,4755|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4750,4755|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|4756,4759|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|4756,4759|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|General Exam|4756,4759|false|false|false|C0001899|Alanine Transaminase|ALT
Finding|Gene or Genome|General Exam|4756,4759|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|General Exam|4756,4759|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|General Exam|4756,4759|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|General Exam|4756,4759|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|General Exam|4763,4766|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|General Exam|4763,4766|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|4763,4766|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|General Exam|4763,4766|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|General Exam|4763,4766|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Finding|Gene or Genome|General Exam|4763,4766|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|4770,4777|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|General Exam|4770,4777|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|General Exam|4805,4810|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4805,4810|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|4811,4817|false|false|false|C0023764|lipase|Lipase
Drug|Enzyme|General Exam|4811,4817|false|false|false|C0023764|lipase|Lipase
Drug|Pharmacologic Substance|General Exam|4811,4817|false|false|false|C0023764|lipase|Lipase
Procedure|Laboratory Procedure|General Exam|4811,4817|false|false|false|C0373670|Lipase measurement|Lipase
Disorder|Disease or Syndrome|General Exam|4834,4839|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4834,4839|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|General Exam|4866,4871|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4866,4871|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|4872,4877|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|General Exam|4872,4877|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|General Exam|4872,4877|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|General Exam|4872,4877|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Finding|Gene or Genome|General Exam|4875,4879|false|false|false|C1413238;C3273407|CD79A gene;CD79A wt Allele|MB-1
Disorder|Disease or Syndrome|General Exam|4906,4911|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4906,4911|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|4906,4919|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|General Exam|4912,4919|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|4912,4919|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|4912,4919|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|4912,4919|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|4912,4919|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Finding|Physiologic Function|General Exam|4912,4919|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|4912,4919|false|false|false|C0201925|Calcium measurement|Calcium
Procedure|Diagnostic Procedure|General Exam|4941,4944|false|false|false|C0039985|Plain chest X-ray|CXR
Anatomy|Body Location or Region|Findings|4995,5000|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Findings|4995,5000|false|false|false|C0741025|Chest problem|chest
Finding|Functional Concept|Findings|5036,5040|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Space or Junction|Findings|5036,5059|false|false|false|C0504100|Left costodiaphragmatic recess|left costophrenic angle
Anatomy|Body Location or Region|Findings|5041,5059|false|false|false|C0230151|Costophrenic angle|costophrenic angle
Finding|Functional Concept|Findings|5070,5080|false|false|false|C0332299|Suggestive of|suggestive
Finding|Functional Concept|Findings|5070,5083|false|false|false|C0332299|Suggestive of|suggestive of
Finding|Pathologic Function|Findings|5096,5104|false|false|false|C0008767;C2004491|Cicatrix;Cicatrization|scarring
Anatomy|Tissue|Findings|5108,5115|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|Findings|5108,5115|false|false|false|C0032226|Pleural Diseases|pleural
Disorder|Disease or Syndrome|Findings|5108,5126|false|false|false|C0264545|Thickening of pleura|pleural thickening
Finding|Finding|Findings|5116,5126|false|false|false|C0205400|Thickened|thickening
Anatomy|Body Part, Organ, or Organ Component|Findings|5133,5138|false|false|false|C0024109|Lung|lungs
Finding|Idea or Concept|Findings|5154,5159|false|false|false|C1550016|Remote control command - Clear|clear
Finding|Functional Concept|Findings|5209,5215|false|false|false|C0439801|Limited (extensiveness)|limits
Procedure|Therapeutic or Preventive Procedure|Findings|5218,5235|false|false|false|C1282959|Median Sternotomy|Median sternotomy
Procedure|Therapeutic or Preventive Procedure|Findings|5225,5235|false|false|false|C0185792|Sternotomy (procedure)|sternotomy
Anatomy|Body Location or Region|Findings|5246,5257|false|false|false|C0025066|Mediastinum|mediastinal
Finding|Intellectual Product|Impression|5297,5302|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Location or Region|Impression|5303,5318|false|false|false|C0553534|Cardiopulmonary|cardiopulmonary
Disorder|Disease or Syndrome|Impression|5303,5318|false|false|false|C4072686|Cardiovascular disease+Pulmonary disease|cardiopulmonary
Anatomy|Body Part, Organ, or Organ Component|Impression|5319,5326|false|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|Impression|5319,5326|true|false|false|C1951340|Process Pharmacologic Substance|process
Finding|Functional Concept|Impression|5319,5326|true|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|Impression|5319,5326|true|false|false|C1522240|Process|process
Finding|Daily or Recreational Activity|Impression|5329,5337|false|false|false|C0015259|Exercise|Exercise
Procedure|Therapeutic or Preventive Procedure|Impression|5329,5337|false|false|false|C1522704|Exercise Pain Management|Exercise
Attribute|Clinical Attribute|Impression|5338,5344|false|false|false|C1718621|W stress|Stress
Drug|Organic Chemical|Impression|5338,5344|false|false|false|C0723460|Stress bismuth subsalicylate|Stress
Drug|Pharmacologic Substance|Impression|5338,5344|false|false|false|C0723460|Stress bismuth subsalicylate|Stress
Finding|Finding|Impression|5338,5344|false|false|false|C0038435|Stress|Stress
Finding|Intellectual Product|Impression|5350,5360|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|Impression|5350,5360|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Finding|Impression|5362,5370|false|false|false|C0741302|atypia morphology|Atypical
Finding|Intellectual Product|Impression|5371,5383|false|false|false|C1272517|Sudden onset (contextual qualifier) (qualifier value)|sudden onset
Finding|Intellectual Product|Impression|5371,5386|false|false|false|C1272517|Sudden onset (contextual qualifier) (qualifier value)|sudden onset of
Anatomy|Body Location or Region|Impression|5387,5392|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Impression|5387,5392|false|false|false|C0741025|Chest problem|chest
Finding|Sign or Symptom|Impression|5387,5402|false|false|false|C0232292|Chest tightness|chest tightness
Finding|Finding|Impression|5422,5432|false|false|false|C0429029|ST segment|ST segment
Finding|Functional Concept|Impression|5433,5440|false|false|false|C0392747|Changing|changes
Finding|Finding|Impression|5453,5456|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Impression|5453,5456|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Daily or Recreational Activity|Impression|5468,5475|false|false|false|C0035253|Rest|Resting
Finding|Intellectual Product|Impression|5476,5480|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Organ or Tissue Function|Impression|5481,5489|false|false|false|C0039155|Systole|systolic
Disorder|Disease or Syndrome|Impression|5481,5502|false|false|false|C0221155|Systolic Hypertension|systolic hypertension
Disorder|Disease or Syndrome|Impression|5490,5502|false|false|false|C0020538|Hypertensive disease|hypertension
Finding|Organ or Tissue Function|Impression|5518,5529|false|false|false|C0019010|Hemodynamics|hemodynamic
Procedure|Laboratory Procedure|Impression|5518,5529|false|false|false|C4281788|hemodynamics (procedure)|hemodynamic
Finding|Finding|Impression|5531,5539|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Intellectual Product|Impression|5531,5539|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Mental Process|Impression|5531,5539|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Organism Function|Impression|5531,5551|false|false|false|C2265833|response to exercise|response to exercise
Finding|Daily or Recreational Activity|Impression|5543,5551|false|false|false|C0015259|Exercise|exercise
Procedure|Therapeutic or Preventive Procedure|Impression|5543,5551|false|false|false|C1522704|Exercise Pain Management|exercise
Procedure|Health Care Activity|Impression|5553,5557|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|Echo
Procedure|Therapeutic or Preventive Procedure|Impression|5553,5557|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|Echo
Attribute|Clinical Attribute|Impression|5558,5564|false|false|false|C4255046||report
Finding|Intellectual Product|Impression|5558,5564|false|false|false|C0684224|Report (document)|report
Procedure|Health Care Activity|Impression|5558,5564|false|false|false|C0700287|Reporting|report
Finding|Daily or Recreational Activity|Impression|5583,5591|false|false|false|C0015259|Exercise|Exercise
Procedure|Therapeutic or Preventive Procedure|Impression|5583,5591|false|false|false|C1522704|Exercise Pain Management|Exercise
Procedure|Health Care Activity|Impression|5592,5596|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|Echo
Procedure|Therapeutic or Preventive Procedure|Impression|5592,5596|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|Echo
Finding|Intellectual Product|Impression|5602,5612|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|Impression|5602,5612|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Intellectual Product|Impression|5614,5618|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|Poor
Finding|Conceptual Entity|Impression|5619,5629|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|functional
Finding|Functional Concept|Impression|5619,5629|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|functional
Finding|Daily or Recreational Activity|Impression|5630,5638|false|false|false|C0015259|Exercise|exercise
Procedure|Therapeutic or Preventive Procedure|Impression|5630,5638|false|false|false|C1522704|Exercise Pain Management|exercise
Drug|Amino Acid, Peptide, or Protein|Impression|5662,5665|false|false|false|C0018064|Equine Gonadotropins|ECG
Drug|Hormone|Impression|5662,5665|false|false|false|C0018064|Equine Gonadotropins|ECG
Drug|Pharmacologic Substance|Impression|5662,5665|false|false|false|C0018064|Equine Gonadotropins|ECG
Finding|Intellectual Product|Impression|5662,5665|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|ECG
Procedure|Diagnostic Procedure|Impression|5662,5665|false|false|false|C1623258|Electrocardiography|ECG
Finding|Functional Concept|Impression|5667,5674|false|false|false|C0392747|Changing|changes
Disorder|Anatomical Abnormality|Impression|5682,5689|false|false|false|C1689985|Absence (morphologic abnormality)|absence
Finding|Functional Concept|Impression|5682,5689|false|false|false|C0332197|Absent|absence
Finding|Functional Concept|Impression|5682,5692|false|false|false|C0332197|Absent|absence of
Finding|Idea or Concept|Impression|5714,5722|false|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Impression|5714,5725|false|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Finding|Functional Concept|Impression|5727,5736|false|false|false|C0205263|Induce (action)|inducible
Finding|Pathologic Function|Impression|5737,5745|false|false|false|C0022116|Ischemia|ischemia
Procedure|Therapeutic or Preventive Procedure|Impression|5737,5745|false|false|false|C4321499|Ischemia Procedure|ischemia
Finding|Finding|Impression|5758,5761|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Impression|5758,5761|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Daily or Recreational Activity|Impression|5772,5779|false|false|false|C0035253|Rest|Resting
Finding|Intellectual Product|Impression|5780,5784|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Organ or Tissue Function|Impression|5786,5794|false|false|false|C0039155|Systole|systolic
Disorder|Disease or Syndrome|Impression|5786,5807|false|false|false|C0221155|Systolic Hypertension|systolic hypertension
Disorder|Disease or Syndrome|Impression|5795,5807|false|false|false|C0020538|Hypertensive disease|hypertension
Finding|Organ or Tissue Function|Impression|5823,5834|false|false|false|C0019010|Hemodynamics|hemodynamic
Procedure|Laboratory Procedure|Impression|5823,5834|false|false|false|C4281788|hemodynamics (procedure)|hemodynamic
Finding|Finding|Impression|5835,5843|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Intellectual Product|Impression|5835,5843|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Mental Process|Impression|5835,5843|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Functional Concept|Impression|5848,5859|false|false|false|C0205463|Physiological|physiologic
Attribute|Clinical Attribute|Impression|5860,5866|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|Impression|5860,5866|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|Impression|5860,5866|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Finding|Finding|Impression|5860,5866|false|false|false|C0038435|Stress|stress
Finding|Body Substance|Impression|5870,5879|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|Impression|5870,5879|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|Impression|5870,5879|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|Impression|5870,5879|false|false|false|C0030685|Patient Discharge|DISCHARGE
Lab|Laboratory or Test Result|Impression|5880,5884|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|Impression|5899,5904|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|Impression|5899,5904|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|Impression|5905,5908|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|Impression|5913,5916|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|Impression|5913,5916|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|Impression|5913,5916|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|Impression|5923,5926|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Impression|5923,5926|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|Impression|5923,5926|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Impression|5923,5926|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|Impression|5932,5935|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|Impression|5932,5935|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|Impression|5943,5946|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|Impression|5943,5946|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|Impression|5943,5946|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|Impression|5943,5946|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|Impression|5950,5953|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|Impression|5950,5953|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|Impression|5950,5953|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|Impression|5950,5953|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|Impression|5950,5953|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|Impression|5960,5964|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|Impression|5979,5982|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|Impression|5999,6004|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|Impression|5999,6004|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Inorganic Chemical|Impression|6034,6038|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|Impression|6034,6038|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|Impression|6034,6038|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|Impression|6064,6069|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|Impression|6064,6069|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|Impression|6101,6105|false|false|false|C0270724|Infantile Neuroaxonal Dystrophy|PLAN
Finding|Functional Concept|Impression|6101,6105|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|PLAN
Finding|Intellectual Product|Impression|6101,6105|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|PLAN
Finding|Mental Process|Impression|6101,6105|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|PLAN
Finding|Finding|Impression|6111,6114|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|pmh
Finding|Finding|Impression|6115,6121|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Impression|6115,6121|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|Impression|6128,6131|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Impression|6128,6131|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Impression|6128,6131|false|false|false|C1504769|DFFB protein, human|CAD
Finding|Gene or Genome|Impression|6128,6131|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Impression|6128,6131|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Impression|6128,6131|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Impression|6128,6131|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Impression|6136,6140|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Finding|Intellectual Product|Impression|6147,6154|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Impression|6147,6154|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Attribute|Clinical Attribute|Impression|6156,6162|false|false|false|C2926611||angina
Finding|Finding|Impression|6156,6162|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Finding|Sign or Symptom|Impression|6156,6162|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Disorder|Disease or Syndrome|Impression|6170,6173|false|false|false|C0020538|Hypertensive disease|HTN
Anatomy|Body Location or Region|Impression|6196,6201|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Impression|6196,6201|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Impression|6196,6206|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Impression|6196,6206|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Impression|6202,6206|false|true|false|C2598155||pain
Finding|Functional Concept|Impression|6202,6206|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Impression|6202,6206|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Hormone|Impression|6223,6232|false|false|false|C3273442|Crescendo|crescendo
Drug|Pharmacologic Substance|Impression|6223,6232|false|false|false|C3273442|Crescendo|crescendo
Disorder|Disease or Syndrome|Impression|6223,6239|false|false|false|C0002965|Angina, Unstable|crescendo angina
Attribute|Clinical Attribute|Impression|6233,6239|false|false|false|C2926611||angina
Finding|Finding|Impression|6233,6239|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Finding|Sign or Symptom|Impression|6233,6239|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Anatomy|Body Location or Region|Impression|6260,6265|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|Impression|6260,6265|false|false|false|C0741025|Chest problem|Chest
Attribute|Clinical Attribute|Impression|6260,6270|false|false|false|C2926613||Chest pain
Finding|Sign or Symptom|Impression|6260,6270|false|false|false|C0008031|Chest Pain|Chest pain
Attribute|Clinical Attribute|Impression|6266,6270|false|false|false|C2598155||pain
Finding|Functional Concept|Impression|6266,6270|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Impression|6266,6270|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Body Substance|Impression|6272,6279|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Impression|6272,6279|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Impression|6272,6279|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|Impression|6285,6289|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|Impression|6285,6289|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|Impression|6285,6289|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Anatomy|Body Part, Organ, or Organ Component|Impression|6290,6298|false|false|false|C0018787|Heart|coronary
Finding|Idea or Concept|Impression|6299,6303|false|false|false|C0035647|Risk|risk
Disorder|Congenital Abnormality|Impression|6320,6323|false|false|false|C0041207|Truncus Arteriosus, Persistent|cat
Drug|Amino Acid, Peptide, or Protein|Impression|6320,6323|false|false|false|C0008169;C1443200;C3530118|CAT protein, human;Cat hair antigen;Chloramphenicol O-Acetyltransferase|cat
Drug|Enzyme|Impression|6320,6323|false|false|false|C0008169;C1443200;C3530118|CAT protein, human;Cat hair antigen;Chloramphenicol O-Acetyltransferase|cat
Drug|Immunologic Factor|Impression|6320,6323|false|false|false|C0008169;C1443200;C3530118|CAT protein, human;Cat hair antigen;Chloramphenicol O-Acetyltransferase|cat
Finding|Gene or Genome|Impression|6320,6323|false|false|false|C1151515;C1366498;C1413138;C4050461;C4758039|CAT gene;Chloramphenicol Acetyl Transferase Gene;Chronic Obstructive Pulmonary Disease Assessment Test scale;Cutaneous Assessment Tool;catalase activity|cat
Finding|Intellectual Product|Impression|6320,6323|false|false|false|C1151515;C1366498;C1413138;C4050461;C4758039|CAT gene;Chloramphenicol Acetyl Transferase Gene;Chronic Obstructive Pulmonary Disease Assessment Test scale;Cutaneous Assessment Tool;catalase activity|cat
Finding|Molecular Function|Impression|6320,6323|false|false|false|C1151515;C1366498;C1413138;C4050461;C4758039|CAT gene;Chloramphenicol Acetyl Transferase Gene;Chronic Obstructive Pulmonary Disease Assessment Test scale;Cutaneous Assessment Tool;catalase activity|cat
Procedure|Diagnostic Procedure|Impression|6320,6323|false|false|false|C0040405;C0280589;C2097305|X-Ray Computed Tomography;allergy testing cat;cytarabine/thioguanine protocol|cat
Procedure|Laboratory Procedure|Impression|6320,6323|false|false|false|C0040405;C0280589;C2097305|X-Ray Computed Tomography;allergy testing cat;cytarabine/thioguanine protocol|cat
Procedure|Therapeutic or Preventive Procedure|Impression|6320,6323|false|false|false|C0040405;C0280589;C2097305|X-Ray Computed Tomography;allergy testing cat;cytarabine/thioguanine protocol|cat
Finding|Gene or Genome|Impression|6334,6337|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Disorder|Disease or Syndrome|Impression|6367,6374|true|false|false|C0012634|Disease|disease
Drug|Amino Acid, Peptide, or Protein|Impression|6377,6381|false|false|false|C5552605|FACT Complex|Fact
Drug|Biologically Active Substance|Impression|6377,6381|false|false|false|C5552605|FACT Complex|Fact
Finding|Gene or Genome|Impression|6377,6381|false|false|false|C1420522;C5551287|SSRP1 wt Allele;SUPT16H gene|Fact
Finding|Finding|Impression|6421,6429|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Finding|Functional Concept|Impression|6421,6429|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Procedure|Health Care Activity|Impression|6421,6429|false|false|false|C0031809|Physical Examination|physical
Finding|Finding|Impression|6421,6434|false|false|false|C1509143|physical examination (physical finding)|physical exam
Procedure|Health Care Activity|Impression|6421,6434|false|false|false|C0031809|Physical Examination|physical exam
Finding|Functional Concept|Impression|6430,6434|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|Impression|6430,6434|false|false|false|C0582103|Medical Examination|exam
Anatomy|Body Part, Organ, or Organ Component|Impression|6449,6456|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|Impression|6449,6456|false|false|false|C1314974|Cardiac attachment|cardiac
Finding|Conceptual Entity|Impression|6457,6462|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Finding|Functional Concept|Impression|6457,6462|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Finding|Functional Concept|Impression|6472,6480|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Impression|6472,6480|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Body Substance|Impression|6500,6507|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Impression|6500,6507|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Impression|6500,6507|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Conceptual Entity|Impression|6511,6518|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Impression|6511,6518|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Impression|6511,6518|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Impression|6511,6521|false|false|false|C0262926|Medical History|history of
Finding|Functional Concept|Impression|6522,6531|false|false|false|C1516691|Cognitive|cognitive
Disorder|Mental or Behavioral Dysfunction|Impression|6522,6542|false|false|false|C0338656|Impaired cognition|cognitive impairment
Finding|Finding|Impression|6532,6542|false|false|false|C0221099;C0684336|Impaired;Impaired health|impairment
Finding|Functional Concept|Impression|6532,6542|false|false|false|C0221099;C0684336|Impaired;Impaired health|impairment
Disorder|Disease or Syndrome|Impression|6557,6560|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Impression|6557,6560|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Impression|6557,6560|false|false|false|C1504769|DFFB protein, human|CAD
Finding|Gene or Genome|Impression|6557,6560|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Impression|6557,6560|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Impression|6557,6560|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Impression|6557,6560|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Finding|Pathologic Function|Impression|6571,6579|false|false|false|C1261287|Stenosis|stenosis
Attribute|Clinical Attribute|Impression|6580,6586|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|Impression|6580,6586|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|Impression|6580,6586|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Finding|Finding|Impression|6580,6586|false|false|false|C0038435|Stress|stress
Procedure|Diagnostic Procedure|Impression|6580,6591|false|false|false|C0920208|Echocardiography, Stress|stress echo
Procedure|Health Care Activity|Impression|6587,6591|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Procedure|Therapeutic or Preventive Procedure|Impression|6587,6591|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Finding|Conceptual Entity|Impression|6620,6630|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|functional
Finding|Functional Concept|Impression|6620,6630|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|functional
Disorder|Congenital Abnormality|Impression|6632,6643|false|false|false|C0000768|Congenital Abnormality|abnormality
Finding|Finding|Impression|6632,6643|false|false|false|C1704258|Abnormality|abnormality
Finding|Organism Function|Impression|6649,6657|false|false|false|C0015264|Exertion|exertion
Procedure|Health Care Activity|Impression|6663,6667|true|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Procedure|Therapeutic or Preventive Procedure|Impression|6663,6667|true|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Disorder|Congenital Abnormality|Impression|6668,6681|true|false|false|C0000768|Congenital Abnormality|abnormalities
Finding|Functional Concept|Impression|6668,6681|true|false|false|C0000769|teratologic|abnormalities
Finding|Finding|Impression|6715,6723|false|false|false|C0741302|atypia morphology|atypical
Finding|Sign or Symptom|Impression|6715,6734|false|true|false|C0262384|Atypical chest pain|atypical chest pain
Anatomy|Body Location or Region|Impression|6724,6729|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Impression|6724,6729|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Impression|6724,6734|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Impression|6724,6734|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Impression|6730,6734|false|true|false|C2598155||pain
Finding|Functional Concept|Impression|6730,6734|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Impression|6730,6734|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|Impression|6740,6746|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|Impression|6740,6746|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|Impression|6740,6746|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Finding|Finding|Impression|6740,6746|false|false|false|C0038435|Stress|stress
Finding|Idea or Concept|Impression|6771,6775|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Impression|6771,6775|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Impression|6771,6775|false|false|false|C1553498|home health encounter|home
Drug|Amino Acid, Peptide, or Protein|Impression|6776,6779|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Enzyme|Impression|6776,6779|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Organic Chemical|Impression|6776,6779|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Pharmacologic Substance|Impression|6776,6779|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Finding|Gene or Genome|Impression|6776,6779|false|false|false|C1412553|ARSA gene|ASA
Drug|Organic Chemical|Impression|6781,6787|false|false|false|C0633084|Plavix|plavix
Drug|Pharmacologic Substance|Impression|6781,6787|false|false|false|C0633084|Plavix|plavix
Drug|Organic Chemical|Impression|6789,6795|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|statin
Drug|Pharmacologic Substance|Impression|6789,6795|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|statin
Finding|Gene or Genome|Impression|6789,6795|false|false|false|C1414273|EEF1A2 gene|statin
Drug|Element, Ion, or Isotope|Impression|6797,6804|false|false|false|C0028125;C0699857;C3848573|Nitrate;Nitrates;nitrate ion|nitrate
Drug|Inorganic Chemical|Impression|6797,6804|false|false|false|C0028125;C0699857;C3848573|Nitrate;Nitrates;nitrate ion|nitrate
Drug|Pharmacologic Substance|Impression|6797,6804|false|false|false|C0028125;C0699857;C3848573|Nitrate;Nitrates;nitrate ion|nitrate
Drug|Organic Chemical|Impression|6809,6819|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|Impression|6809,6819|false|false|false|C0025859|metoprolol|metoprolol
Finding|Idea or Concept|Impression|6827,6835|false|false|false|C4288901|In-House|in-house
Finding|Gene or Genome|Impression|6859,6863|false|false|false|C1420621;C1515258|TCAP gene;Telephone Number|tele
Finding|Intellectual Product|Impression|6859,6863|false|false|false|C1420621;C1515258|TCAP gene;Telephone Number|tele
Finding|Intellectual Product|Impression|6876,6882|true|false|false|C3484361|Alarms (package insert)|alarms
Finding|Idea or Concept|Impression|6905,6909|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Impression|6905,6909|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Impression|6905,6909|false|false|false|C1553498|home health encounter|home
Finding|Classification|Impression|6918,6926|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Impression|6918,6926|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Impression|6918,6926|false|false|false|C5237010|Expression Negative|negative
Attribute|Clinical Attribute|Impression|6927,6933|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|Impression|6927,6933|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|Impression|6927,6933|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Finding|Finding|Impression|6927,6933|false|false|false|C0038435|Stress|stress
Finding|Functional Concept|Impression|6937,6943|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|Impression|6937,6943|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|Impression|6937,6946|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|Impression|6937,6946|false|false|false|C1522577|follow-up|follow-up
Disorder|Disease or Syndrome|Impression|6957,6960|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|Impression|6957,6960|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|Impression|6957,6960|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|Impression|6957,6960|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|Impression|6957,6960|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|Impression|6957,6960|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|Impression|6957,6960|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|Impression|6957,6960|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Finding|Gene or Genome|Impression|6957,6960|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|Impression|6957,6960|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Intellectual Product|Impression|6971,6978|false|false|false|C1547296|Chronic - Admission Level of Care Code|CHRONIC
Procedure|Health Care Activity|Impression|6971,6978|false|false|false|C1555457|Provision of recurring care for chronic illness|CHRONIC
Attribute|Clinical Attribute|Impression|6992,7001|false|false|false|C0012000|Diastole|Diastolic
Disorder|Disease or Syndrome|Impression|6992,7005|false|false|false|C2183328|diastolic congestive heart failure|Diastolic CHF
Anatomy|Body Space or Junction|Impression|7002,7005|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|Impression|7002,7005|false|false|false|C0018802|Congestive heart failure|CHF
Finding|Finding|Impression|7019,7024|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Impression|7019,7024|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Drug|Substance|Impression|7028,7033|true|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Impression|7028,7033|true|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Finding|Impression|7028,7042|true|false|false|C0546817;C5848920|Fluid Overload;Hypervolemia (finding)|fluid overload
Finding|Pathologic Function|Impression|7028,7042|true|false|false|C0546817;C5848920|Fluid Overload;Hypervolemia (finding)|fluid overload
Drug|Biomedical or Dental Material|Impression|7063,7071|false|false|false|C0168634|BaseLine dental cement|baseline
Finding|Idea or Concept|Impression|7063,7071|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Organ or Tissue Function|Impression|7072,7080|false|false|false|C0012797|Diuresis|diuresis
Finding|Idea or Concept|Impression|7104,7108|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Impression|7104,7108|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Impression|7104,7108|false|false|false|C1553498|home health encounter|home
Finding|Finding|Impression|7145,7150|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Impression|7145,7150|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Finding|Impression|7154,7168|false|false|false|C0231187|Decompensation|decompensation
Finding|Organ or Tissue Function|Impression|7186,7194|false|false|false|C0012797|Diuresis|diuresis
Disorder|Disease or Syndrome|Impression|7200,7208|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|Diabetes
Finding|Intellectual Product|Impression|7211,7215|false|false|false|C0019972|Hospital Information Systems|HISS
Finding|Idea or Concept|Impression|7216,7224|false|false|false|C4288901|In-House|in-house
Finding|Idea or Concept|Impression|7252,7256|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Impression|7252,7256|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Impression|7252,7256|false|false|false|C1553498|home health encounter|home
Drug|Amino Acid, Peptide, or Protein|Impression|7258,7265|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|Impression|7258,7265|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|Impression|7258,7265|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Finding|Gene or Genome|Impression|7258,7265|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|Impression|7258,7265|false|false|false|C0202098|Insulin measurement|insulin
Finding|Intellectual Product|Impression|7266,7273|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|Impression|7266,7273|false|false|false|C0040808|Treatment Protocols|regimen
Drug|Amino Acid, Peptide, or Protein|Impression|7282,7288|false|false|false|C0876064|Lantus|lantus
Drug|Pharmacologic Substance|Impression|7282,7288|false|false|false|C0876064|Lantus|lantus
Attribute|Clinical Attribute|Impression|7297,7308|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Impression|7297,7308|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Impression|7297,7308|false|false|false|C4284232|Medications|Medications
Finding|Finding|Impression|7297,7321|false|false|false|C1627937|Medications on admission|Medications on Admission
Procedure|Health Care Activity|Impression|7312,7321|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|Impression|7340,7350|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Impression|7340,7350|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|Impression|7340,7355|false|false|false|C0746470|MEDICATION LIST|Medication list
Finding|Intellectual Product|Impression|7351,7355|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Drug|Organic Chemical|Impression|7372,7380|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Impression|7372,7380|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Impression|7372,7380|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Finding|Functional Concept|Impression|7372,7380|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Impression|7372,7380|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|Impression|7385,7393|false|false|false|C0126174|losartan|Losartan
Drug|Pharmacologic Substance|Impression|7385,7393|false|false|false|C0126174|losartan|Losartan
Drug|Organic Chemical|Impression|7385,7403|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Pharmacologic Substance|Impression|7385,7403|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Biologically Active Substance|Impression|7394,7403|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|Impression|7394,7403|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|Impression|7394,7403|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|Impression|7394,7403|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|Impression|7394,7403|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Finding|Physiologic Function|Impression|7394,7403|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|Impression|7394,7403|false|false|false|C0202194|Potassium measurement|Potassium
Drug|Organic Chemical|Impression|7423,7430|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Impression|7423,7430|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|Impression|7450,7462|false|false|false|C0007248|carisoprodol|carisoprodol
Drug|Pharmacologic Substance|Impression|7450,7462|false|false|false|C0007248|carisoprodol|carisoprodol
Anatomy|Body Space or Junction|Impression|7475,7479|false|false|false|C0226896|Oral cavity|Oral
Drug|Biomedical or Dental Material|Impression|7475,7479|false|false|false|C1272919|Oral Dosage Form|Oral
Finding|Finding|Impression|7475,7479|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Finding|Functional Concept|Impression|7475,7479|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Finding|Gene or Genome|Impression|7484,7489|false|false|false|C0037763;C3812627|KANTR gene;Spasm|spasm
Finding|Sign or Symptom|Impression|7484,7489|false|false|false|C0037763;C3812627|KANTR gene;Spasm|spasm
Drug|Biomedical or Dental Material|Impression|7498,7504|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Gene or Genome|Impression|7519,7522|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Part, Organ, or Organ Component|Impression|7523,7529|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|Impression|7523,7529|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Finding|Sign or Symptom|Impression|7523,7535|false|false|false|C0037763|Spasm|muscle spasm
Finding|Gene or Genome|Impression|7530,7535|false|false|false|C0037763;C3812627|KANTR gene;Spasm|spasm
Finding|Sign or Symptom|Impression|7530,7535|false|false|false|C0037763;C3812627|KANTR gene;Spasm|spasm
Drug|Organic Chemical|Impression|7540,7552|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Pharmacologic Substance|Impression|7540,7552|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Organic Chemical|Impression|7571,7580|false|false|false|C0040805|trazodone|traZODONE
Drug|Pharmacologic Substance|Impression|7571,7580|false|false|false|C0040805|trazodone|traZODONE
Drug|Organic Chemical|Impression|7597,7606|false|false|false|C0030049|oxycodone|Oxycodone
Drug|Pharmacologic Substance|Impression|7597,7606|false|false|false|C0030049|oxycodone|Oxycodone
Procedure|Laboratory Procedure|Impression|7597,7606|false|false|false|C0524222|Oxycodone measurement|Oxycodone
Drug|Pharmacologic Substance|Impression|7597,7620|false|false|false|C0717368|acetaminophen / oxycodone|Oxycodone-Acetaminophen
Drug|Organic Chemical|Impression|7607,7620|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Impression|7607,7620|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Procedure|Laboratory Procedure|Impression|7607,7620|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Biomedical or Dental Material|Impression|7635,7638|false|false|false|C0039225|Tablet Dosage Form|TAB
Finding|Gene or Genome|Impression|7646,7649|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Impression|7650,7654|false|false|false|C2598155||pain
Finding|Functional Concept|Impression|7650,7654|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Impression|7650,7654|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Impression|7659,7671|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Impression|7659,7671|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|Impression|7691,7704|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Pharmacologic Substance|Impression|7691,7704|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Finding|Gene or Genome|Impression|7718,7721|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Location or Region|Impression|7722,7727|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Impression|7722,7727|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Impression|7722,7732|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Impression|7722,7732|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Impression|7728,7732|false|true|false|C2598155||pain
Finding|Functional Concept|Impression|7728,7732|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Impression|7728,7732|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Impression|7737,7747|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|Impression|7737,7747|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|Impression|7737,7757|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Pharmacologic Substance|Impression|7737,7757|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Organic Chemical|Impression|7748,7757|false|false|false|C0038617;C0220918|Succinates;succinate|Succinate
Drug|Organic Chemical|Impression|7782,7792|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|Impression|7782,7792|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|Impression|7782,7804|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|Impression|7782,7804|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Finding|Finding|Impression|7806,7814|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Impression|7806,7814|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Impression|7815,7822|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Impression|7815,7822|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Impression|7815,7822|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Impression|7845,7856|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Pharmacologic Substance|Impression|7845,7856|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Organic Chemical|Impression|7877,7888|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Impression|7877,7888|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Organic Chemical|Impression|7877,7899|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|Impression|7877,7899|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|Impression|7889,7899|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Disorder|Mental or Behavioral Dysfunction|Impression|7917,7920|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Impression|7917,7920|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Impression|7917,7920|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Impression|7917,7920|false|false|false|C1332410|BID gene|BID
Drug|Amino Acid, Peptide, or Protein|Impression|7949,7956|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Hormone|Impression|7949,7956|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Pharmacologic Substance|Impression|7949,7956|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Finding|Gene or Genome|Impression|7949,7956|false|false|false|C1337112|INS gene|Insulin
Procedure|Laboratory Procedure|Impression|7949,7956|false|false|false|C0202098|Insulin measurement|Insulin
Finding|Functional Concept|Impression|7960,7967|false|false|false|C0332246|Sliding|Sliding
Procedure|Therapeutic or Preventive Procedure|Impression|7960,7973|false|false|false|C2937251|sliding scale|Sliding Scale
Anatomy|Body Part, Organ, or Organ Component|Impression|7968,7973|false|false|false|C0222045|Integumentary scale|Scale
Event|Activity|Impression|7968,7973|false|false|false|C1947916|Scaling|Scale
Finding|Conceptual Entity|Impression|7968,7973|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|Scale
Finding|Intellectual Product|Impression|7968,7973|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|Scale
Finding|Functional Concept|Impression|8000,8008|false|false|false|C1547671|Override|Override
Finding|Idea or Concept|Impression|8010,8016|false|false|false|C0392360|Indication of (contextual qualifier)|Reason
Drug|Amino Acid, Peptide, or Protein|Impression|8018,8025|false|false|false|C1314782|Levemir|Levemir
Drug|Hormone|Impression|8018,8025|false|false|false|C1314782|Levemir|Levemir
Drug|Pharmacologic Substance|Impression|8018,8025|false|false|false|C1314782|Levemir|Levemir
Finding|Intellectual Product|Impression|8040,8048|false|false|false|C1547997;C3244303|Diagnostic Service Section ID - Pharmacy;Pharmacy domain|pharmacy
Procedure|Health Care Activity|Impression|8040,8048|false|false|false|C0031321|Pharmaceutical Services|pharmacy
Finding|Intellectual Product|Impression|8049,8053|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Finding|Body Substance|Impression|8057,8066|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Impression|8057,8066|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Impression|8057,8066|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Impression|8057,8066|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Impression|8057,8078|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Impression|8067,8078|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Impression|8067,8078|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Impression|8067,8078|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Impression|8083,8090|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Impression|8083,8090|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|Impression|8110,8122|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Impression|8110,8122|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|Impression|8142,8153|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Pharmacologic Substance|Impression|8142,8153|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Organic Chemical|Impression|8173,8184|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Impression|8173,8184|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Organic Chemical|Impression|8173,8195|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|Impression|8173,8195|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|Impression|8185,8195|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Disorder|Mental or Behavioral Dysfunction|Impression|8213,8216|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Impression|8213,8216|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Impression|8213,8216|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Impression|8213,8216|false|false|false|C1332410|BID gene|BID
Drug|Amino Acid, Peptide, or Protein|Impression|8244,8251|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Hormone|Impression|8244,8251|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Pharmacologic Substance|Impression|8244,8251|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Finding|Gene or Genome|Impression|8244,8251|false|false|false|C1337112|INS gene|Insulin
Procedure|Laboratory Procedure|Impression|8244,8251|false|false|false|C0202098|Insulin measurement|Insulin
Finding|Functional Concept|Impression|8255,8262|false|false|false|C0332246|Sliding|Sliding
Procedure|Therapeutic or Preventive Procedure|Impression|8255,8268|false|false|false|C2937251|sliding scale|Sliding Scale
Anatomy|Body Part, Organ, or Organ Component|Impression|8263,8268|false|false|false|C0222045|Integumentary scale|Scale
Event|Activity|Impression|8263,8268|false|false|false|C1947916|Scaling|Scale
Finding|Conceptual Entity|Impression|8263,8268|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|Scale
Finding|Intellectual Product|Impression|8263,8268|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|Scale
Finding|Functional Concept|Impression|8295,8303|false|false|false|C1547671|Override|Override
Finding|Idea or Concept|Impression|8305,8311|false|false|false|C0392360|Indication of (contextual qualifier)|Reason
Drug|Amino Acid, Peptide, or Protein|Impression|8313,8320|false|false|false|C1314782|Levemir|Levemir
Drug|Hormone|Impression|8313,8320|false|false|false|C1314782|Levemir|Levemir
Drug|Pharmacologic Substance|Impression|8313,8320|false|false|false|C1314782|Levemir|Levemir
Finding|Intellectual Product|Impression|8335,8343|false|false|false|C1547997;C3244303|Diagnostic Service Section ID - Pharmacy;Pharmacy domain|pharmacy
Procedure|Health Care Activity|Impression|8335,8343|false|false|false|C0031321|Pharmaceutical Services|pharmacy
Finding|Intellectual Product|Impression|8344,8348|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Drug|Organic Chemical|Impression|8353,8361|false|false|false|C0126174|losartan|Losartan
Drug|Pharmacologic Substance|Impression|8353,8361|false|false|false|C0126174|losartan|Losartan
Drug|Organic Chemical|Impression|8353,8371|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Pharmacologic Substance|Impression|8353,8371|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Biologically Active Substance|Impression|8362,8371|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|Impression|8362,8371|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|Impression|8362,8371|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|Impression|8362,8371|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|Impression|8362,8371|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Finding|Physiologic Function|Impression|8362,8371|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|Impression|8362,8371|false|false|false|C0202194|Potassium measurement|Potassium
Drug|Organic Chemical|Impression|8391,8404|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Pharmacologic Substance|Impression|8391,8404|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Finding|Gene or Genome|Impression|8418,8421|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Location or Region|Impression|8422,8427|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Impression|8422,8427|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Impression|8422,8432|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Impression|8422,8432|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Impression|8428,8432|false|true|false|C2598155||pain
Finding|Functional Concept|Impression|8428,8432|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Impression|8428,8432|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Impression|8437,8449|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Pharmacologic Substance|Impression|8437,8449|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Organic Chemical|Impression|8468,8477|false|false|false|C0040805|trazodone|traZODONE
Drug|Pharmacologic Substance|Impression|8468,8477|false|false|false|C0040805|trazodone|traZODONE
Drug|Organic Chemical|Impression|8495,8507|false|false|false|C0007248|carisoprodol|carisoprodol
Drug|Pharmacologic Substance|Impression|8495,8507|false|false|false|C0007248|carisoprodol|carisoprodol
Anatomy|Body Space or Junction|Impression|8520,8524|false|false|false|C0226896|Oral cavity|Oral
Drug|Biomedical or Dental Material|Impression|8520,8524|false|false|false|C1272919|Oral Dosage Form|Oral
Finding|Finding|Impression|8520,8524|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Finding|Functional Concept|Impression|8520,8524|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Finding|Gene or Genome|Impression|8529,8534|false|false|false|C0037763;C3812627|KANTR gene;Spasm|spasm
Finding|Sign or Symptom|Impression|8529,8534|false|false|false|C0037763;C3812627|KANTR gene;Spasm|spasm
Drug|Organic Chemical|Impression|8540,8550|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|Impression|8540,8550|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|Impression|8540,8560|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Pharmacologic Substance|Impression|8540,8560|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Organic Chemical|Impression|8551,8560|false|false|false|C0038617;C0220918|Succinates;succinate|Succinate
Drug|Organic Chemical|Impression|8585,8594|false|false|false|C0030049|oxycodone|Oxycodone
Drug|Pharmacologic Substance|Impression|8585,8594|false|false|false|C0030049|oxycodone|Oxycodone
Procedure|Laboratory Procedure|Impression|8585,8594|false|false|false|C0524222|Oxycodone measurement|Oxycodone
Drug|Pharmacologic Substance|Impression|8585,8608|false|false|false|C0717368|acetaminophen / oxycodone|Oxycodone-Acetaminophen
Drug|Organic Chemical|Impression|8595,8608|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Impression|8595,8608|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Procedure|Laboratory Procedure|Impression|8595,8608|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Biomedical or Dental Material|Impression|8623,8626|false|false|false|C0039225|Tablet Dosage Form|TAB
Finding|Gene or Genome|Impression|8634,8637|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Impression|8638,8642|false|false|false|C2598155||pain
Finding|Functional Concept|Impression|8638,8642|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Impression|8638,8642|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Impression|8648,8658|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|Impression|8648,8658|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|Impression|8648,8670|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|Impression|8648,8670|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Finding|Finding|Impression|8672,8680|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Impression|8672,8680|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Impression|8681,8688|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Impression|8681,8688|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Impression|8681,8688|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Finding|Body Substance|Impression|8709,8718|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Impression|8709,8718|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Impression|8709,8718|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Impression|8709,8718|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Impression|8709,8730|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Impression|8709,8730|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Impression|8719,8730|false|false|false|C2926604||Disposition
Procedure|Health Care Activity|Impression|8719,8730|false|false|false|C0184758|Patient disposition|Disposition
Finding|Idea or Concept|Impression|8732,8736|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Impression|8732,8736|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Impression|8732,8736|false|false|false|C1553498|home health encounter|Home
Finding|Body Substance|Impression|8739,8748|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Impression|8739,8748|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Impression|8739,8748|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Impression|8739,8748|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Impression|8739,8758|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Impression|8749,8758|false|false|false|C0945731||Diagnosis
Finding|Classification|Impression|8749,8758|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Impression|8749,8758|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Impression|8749,8758|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Finding|Impression|8760,8768|false|false|false|C0741302|atypia morphology|Atypical
Finding|Sign or Symptom|Impression|8760,8779|false|false|false|C0262384|Atypical chest pain|Atypical Chest Pain
Anatomy|Body Location or Region|Impression|8769,8774|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|Impression|8769,8774|false|false|false|C0741025|Chest problem|Chest
Attribute|Clinical Attribute|Impression|8769,8779|false|false|false|C2926613||Chest Pain
Finding|Sign or Symptom|Impression|8769,8779|false|false|false|C0008031|Chest Pain|Chest Pain
Attribute|Clinical Attribute|Impression|8775,8779|false|true|false|C2598155||Pain
Finding|Functional Concept|Impression|8775,8779|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Impression|8775,8779|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Attribute|Clinical Attribute|Discharge Condition|8804,8826|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|8804,8826|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Finding|Finding|Discharge Condition|8813,8826|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|8813,8826|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|8828,8833|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|8828,8833|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|8828,8833|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|Discharge Condition|8828,8833|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|8828,8833|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|8828,8833|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|8838,8849|false|false|false|C1704675|Interaction|interactive
Finding|Mental Process|Discharge Condition|8851,8857|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|8851,8864|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|8851,8864|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|8858,8864|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|8858,8864|false|false|false|C1546481|What subject filter - Status|Status
Disorder|Mental or Behavioral Dysfunction|Discharge Condition|8866,8874|false|false|false|C0009676|Confusion|Confused
Finding|Finding|Discharge Condition|8866,8874|false|false|false|C0683369;C1547301|Clouded consciousness;Precaution Code - Confused|Confused
Finding|Intellectual Product|Discharge Condition|8866,8874|false|false|false|C0683369;C1547301|Clouded consciousness;Precaution Code - Confused|Confused
Event|Activity|Discharge Condition|8888,8896|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|8888,8896|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|8888,8896|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|8897,8903|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|8897,8903|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|Discharge Condition|8905,8915|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|8905,8915|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|8905,8915|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|8905,8915|false|false|false|C1561560|ambulatory encounter|Ambulatory
Finding|Finding|Discharge Condition|8918,8929|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Condition|8918,8929|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Instructions|8984,8992|false|false|false|C1547192|Organization unit type - Hospital|hospital
Anatomy|Body Location or Region|Discharge Instructions|8998,9003|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Discharge Instructions|8998,9003|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Discharge Instructions|8998,9008|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Discharge Instructions|8998,9008|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Discharge Instructions|9004,9008|false|false|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|9004,9008|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|9004,9008|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Gene or Genome|Discharge Instructions|9019,9022|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|lab
Finding|Intellectual Product|Discharge Instructions|9019,9022|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|lab
Anatomy|Body Location or Region|Discharge Instructions|9023,9029|false|false|false|C0817096|Chest|chests
Finding|Intellectual Product|Discharge Instructions|9035,9038|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|Discharge Instructions|9035,9038|false|false|false|C1623258|Electrocardiography|EKG
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|9089,9094|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|9089,9094|false|true|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Discharge Instructions|9089,9094|false|true|false|C0795691|HEART PROBLEM|heart
Finding|Finding|Discharge Instructions|9096,9102|false|false|false|C1261512;C1304680|Attack (finding);Attack behavior|attack
Finding|Social Behavior|Discharge Instructions|9096,9102|false|false|false|C1261512;C1304680|Attack (finding);Attack behavior|attack
Attribute|Clinical Attribute|Discharge Instructions|9136,9142|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|Discharge Instructions|9136,9142|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|Discharge Instructions|9136,9142|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Finding|Finding|Discharge Instructions|9136,9142|false|false|false|C0038435|Stress|stress
Procedure|Diagnostic Procedure|Discharge Instructions|9136,9147|false|false|false|C0015260;C3494508|Exercise stress test;Stress Test|stress test
Anatomy|Body Location or Region|Discharge Instructions|9143,9147|false|false|false|C4318744|Test - temporal region|test
Finding|Functional Concept|Discharge Instructions|9143,9147|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|Discharge Instructions|9143,9147|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|Discharge Instructions|9143,9147|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|Discharge Instructions|9143,9147|false|false|false|C0022885|Laboratory Procedures|test
Finding|Idea or Concept|Discharge Instructions|9175,9183|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Discharge Instructions|9175,9186|true|true|false|C0332120|Evidence of (contextual qualifier)|evidence of
Finding|Idea or Concept|Discharge Instructions|9187,9196|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|9197,9205|false|false|false|C0018787|Heart|coronary
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|9197,9212|false|false|false|C0205042|Coronary artery|coronary artery
Disorder|Disease or Syndrome|Discharge Instructions|9197,9220|true|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|coronary artery disease
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|9206,9212|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|Discharge Instructions|9206,9212|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Disorder|Disease or Syndrome|Discharge Instructions|9206,9220|false|false|false|C0852949|Arteriopathic disease|artery disease
Disorder|Disease or Syndrome|Discharge Instructions|9213,9220|false|false|false|C0012634|Disease|disease
Anatomy|Body Location or Region|Discharge Instructions|9229,9234|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Discharge Instructions|9229,9234|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Discharge Instructions|9229,9239|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Discharge Instructions|9229,9239|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Discharge Instructions|9235,9239|false|false|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|9235,9239|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|9235,9239|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Functional Concept|Discharge Instructions|9262,9270|false|false|false|C2584295|Touching|touching
Anatomy|Body Location or Region|Discharge Instructions|9276,9281|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Discharge Instructions|9276,9281|false|false|false|C0741025|Chest problem|chest
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|9308,9316|false|false|false|C0018787|Heart|coronary
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|9308,9323|false|false|false|C0205042|Coronary artery|coronary artery
Disorder|Disease or Syndrome|Discharge Instructions|9308,9331|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|coronary artery disease
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|9317,9323|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|Discharge Instructions|9317,9323|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Disorder|Disease or Syndrome|Discharge Instructions|9317,9331|false|false|false|C0852949|Arteriopathic disease|artery disease
Disorder|Disease or Syndrome|Discharge Instructions|9324,9331|false|false|false|C0012634|Disease|disease
Attribute|Clinical Attribute|Discharge Instructions|9332,9336|false|false|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|9332,9336|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|9332,9336|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Discharge Instructions|9344,9350|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Discharge Instructions|9344,9350|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Drug|Organic Chemical|Discharge Instructions|9355,9362|false|false|false|C0163712|Relate - vinyl resin|related
Finding|Finding|Discharge Instructions|9355,9362|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|Discharge Instructions|9355,9362|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Attribute|Clinical Attribute|Discharge Instructions|9366,9381|false|false|false|C2707260||musculoskeletal
Finding|Functional Concept|Discharge Instructions|9366,9381|false|false|false|C0497254|Musculoskeletal|musculoskeletal
Finding|Finding|Discharge Instructions|9366,9386|false|false|false|C0026858|Musculoskeletal Pain|musculoskeletal pain
Attribute|Clinical Attribute|Discharge Instructions|9382,9386|false|false|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|9382,9386|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|9382,9386|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Functional Concept|Discharge Instructions|9395,9402|false|false|false|C0392747|Changing|changes
Drug|Pharmacologic Substance|Discharge Instructions|9426,9436|false|false|false|C0013227|Pharmaceutical Preparations|medication
Finding|Intellectual Product|Discharge Instructions|9426,9436|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Finding|Intellectual Product|Discharge Instructions|9426,9441|false|false|false|C0746470|MEDICATION LIST|medication list
Finding|Intellectual Product|Discharge Instructions|9437,9441|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Procedure|Health Care Activity|Discharge Instructions|9452,9460|false|false|false|C1522577|follow-up|followup
Drug|Pharmacologic Substance|Discharge Instructions|9496,9506|false|false|false|C0013227|Pharmaceutical Preparations|medication
Finding|Intellectual Product|Discharge Instructions|9496,9506|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Finding|Functional Concept|Discharge Instructions|9507,9514|false|false|false|C0392747|Changing|changes
Procedure|Health Care Activity|Discharge Instructions|9518,9526|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|9527,9539|false|false|false|C3263700||Instructions
Finding|Intellectual Product|Discharge Instructions|9527,9539|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

