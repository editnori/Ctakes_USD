 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|29,33
No|34,36
:|36,37
_|40,41
_|41,42
_|42,43
<EOL>|43,44
<EOL>|45,46
Admission|46,55
Date|56,60
:|60,61
_|63,64
_|64,65
_|65,66
Discharge|80,89
Date|90,94
:|94,95
_|98,99
_|99,100
_|100,101
<EOL>|101,102
<EOL>|103,104
Date|104,108
of|109,111
Birth|112,117
:|117,118
_|120,121
_|121,122
_|122,123
Sex|136,139
:|139,140
F|143,144
<EOL>|144,145
<EOL>|146,147
Service|147,154
:|154,155
MEDICINE|156,164
<EOL>|164,165
<EOL>|166,167
Allergies|167,176
:|176,177
<EOL>|178,179
Codeine|179,186
<EOL>|186,187
<EOL>|188,189
Attending|189,198
:|198,199
_|200,201
_|201,202
_|202,203
<EOL>|203,204
<EOL>|205,206
Chief|206,211
Complaint|212,221
:|221,222
<EOL>|222,223
Difficulty|223,233
in|234,236
breathing|237,246
<EOL>|246,247
<EOL>|248,249
Major|249,254
Surgical|255,263
or|264,266
Invasive|267,275
Procedure|276,285
:|285,286
<EOL>|286,287
none|287,291
<EOL>|291,292
<EOL>|292,293
<EOL>|294,295
History|295,302
of|303,305
Present|306,313
Illness|314,321
:|321,322
<EOL>|322,323
The|323,326
patient|327,334
is|335,337
a|338,339
_|340,341
_|341,342
_|342,343
year|344,348
-|348,349
old|349,352
female|353,359
with|360,364
a|365,366
history|367,374
of|375,377
NSCLC|378,383
<EOL>|384,385
(|385,386
stage|386,391
IV|392,394
)|394,395
who|396,399
presents|400,408
with|409,413
shortness|414,423
of|424,426
breath|427,433
.|433,434
<EOL>|434,435
.|435,436
<EOL>|436,437
The|437,440
patient|441,448
was|449,452
in|453,455
her|456,459
usual|460,465
state|466,471
of|472,474
health|475,481
until|482,487
the|488,491
evening|492,499
<EOL>|500,501
before|501,507
admission|508,517
when|518,522
she|523,526
began|527,532
to|533,535
feel|536,540
somewhat|541,549
short|550,555
of|556,558
<EOL>|559,560
breath|560,566
.|566,567
The|569,572
next|573,577
morning|578,585
,|585,586
this|587,591
sensation|592,601
persisted|602,611
,|611,612
so|613,615
she|616,619
<EOL>|620,621
became|621,627
concerned|628,637
.|637,638
She|640,643
also|644,648
reports|649,656
a|657,658
few|659,662
day|663,666
history|667,674
of|675,677
a|678,679
<EOL>|680,681
non-productive|681,695
cough|696,701
.|701,702
Denies|704,710
sick|711,715
contacts|716,724
,|724,725
recent|726,732
travel|733,739
or|740,742
<EOL>|743,744
sedentary|744,753
lifestyle|754,763
.|763,764
She|766,769
denied|770,776
chest|777,782
pain|783,787
,|787,788
fever|789,794
,|794,795
chills|796,802
,|802,803
<EOL>|804,805
dizziness|805,814
,|814,815
lightheadedness|816,831
or|832,834
syncope|835,842
.|842,843
She|845,848
presented|849,858
to|859,861
the|862,865
ED|866,868
<EOL>|869,870
where|870,875
she|876,879
was|880,883
found|884,889
to|890,892
be|893,895
hypoxic|896,903
to|904,906
the|907,910
_|911,912
_|912,913
_|913,914
on|915,917
room|918,922
air|923,926
.|926,927
<EOL>|927,928
.|928,929
<EOL>|931,932
In|932,934
the|935,938
ED|939,941
,|941,942
she|943,946
was|947,950
placed|951,957
on|958,960
a|961,962
non-rebreather|963,977
with|978,982
sats|983,987
up|988,990
to|991,993
<EOL>|994,995
the|995,998
high|999,1003
90's|1004,1008
.|1008,1009
Attempts|1011,1019
were|1020,1024
made|1025,1029
to|1030,1032
wean|1033,1037
her|1038,1041
to|1042,1044
NC|1045,1047
but|1048,1051
they|1052,1056
<EOL>|1057,1058
were|1058,1062
unsuccessful|1063,1075
,|1075,1076
as|1077,1079
she|1080,1083
was|1084,1087
satting|1088,1095
88|1096,1098
%|1098,1099
on|1100,1102
4L|1103,1105
NC|1106,1108
.|1108,1109
She|1111,1114
<EOL>|1115,1116
remained|1116,1124
afebrile|1125,1133
in|1134,1136
the|1137,1140
ED|1141,1143
but|1144,1147
was|1148,1151
found|1152,1157
to|1158,1160
have|1161,1165
WBC|1166,1169
of|1170,1172
17|1173,1175
.|1175,1176
<EOL>|1178,1179
Given|1179,1184
that|1185,1189
,|1189,1190
she|1191,1194
received|1195,1203
levofloxacin|1204,1216
and|1217,1220
vancomycin|1221,1231
.|1231,1232
Blood|1234,1239
<EOL>|1240,1241
cultures|1241,1249
were|1250,1254
drawn|1255,1260
prior|1261,1266
to|1267,1269
antibiotic|1270,1280
administration|1281,1295
.|1295,1296
CXR|1298,1301
did|1302,1305
<EOL>|1306,1307
not|1307,1310
show|1311,1315
PNA|1316,1319
,|1319,1320
but|1321,1324
demonstrated|1325,1337
progression|1338,1349
of|1350,1352
known|1353,1358
lung|1359,1363
cancer|1364,1370
.|1370,1371
<EOL>|1372,1373
She|1374,1377
underwent|1378,1387
a|1388,1389
CT|1390,1392
head|1393,1397
to|1398,1400
rule|1401,1405
out|1406,1409
metastases|1410,1420
,|1420,1421
which|1422,1427
was|1428,1431
<EOL>|1432,1433
negative|1433,1441
.|1441,1442
On|1444,1446
transfer|1447,1455
,|1455,1456
patient|1457,1464
was|1465,1468
afebrile|1469,1477
with|1478,1482
HR|1483,1485
-|1485,1486
77|1487,1489
,|1489,1490
BP|1491,1493
-|1493,1494
<EOL>|1495,1496
112|1496,1499
/|1499,1500
49|1500,1502
,|1502,1503
RR|1504,1506
-|1506,1507
16|1508,1510
,|1510,1511
SaO2|1512,1516
-|1516,1517
98|1518,1520
%|1520,1521
on|1522,1524
15L|1525,1528
NRB|1529,1532
<EOL>|1534,1535
.|1535,1536
<EOL>|1536,1537
On|1537,1539
transfer|1540,1548
to|1549,1551
the|1552,1555
ICU|1556,1559
,|1559,1560
the|1561,1564
patient|1565,1572
was|1573,1576
stable|1577,1583
and|1584,1587
comfortable|1588,1599
.|1599,1600
<EOL>|1602,1603
Sats|1603,1607
were|1608,1612
97|1613,1615
%|1615,1616
on|1617,1619
5L|1620,1622
NC|1623,1625
and|1626,1629
95|1630,1632
%|1632,1633
high|1634,1638
-|1638,1639
flow|1639,1643
with|1644,1648
a|1649,1650
face|1651,1655
-|1655,1656
tent|1656,1660
.|1660,1661
<EOL>|1663,1664
.|1664,1665
<EOL>|1667,1668
ROS|1668,1671
:|1671,1672
The|1673,1676
patient|1677,1684
denies|1685,1691
any|1692,1695
fevers|1696,1702
,|1702,1703
chills|1704,1710
,|1710,1711
weight|1712,1718
change|1719,1725
,|1725,1726
<EOL>|1727,1728
nausea|1728,1734
,|1734,1735
vomiting|1736,1744
,|1744,1745
abdominal|1746,1755
pain|1756,1760
,|1760,1761
diarrhea|1762,1770
,|1770,1771
constipation|1772,1784
,|1784,1785
<EOL>|1786,1787
melena|1787,1793
,|1793,1794
hematochezia|1795,1807
,|1807,1808
chest|1809,1814
pain|1815,1819
,|1819,1820
orthopnea|1821,1830
,|1830,1831
PND|1832,1835
,|1835,1836
lower|1837,1842
<EOL>|1843,1844
extremity|1844,1853
edema|1854,1859
,|1859,1860
cough|1861,1866
,|1866,1867
urinary|1868,1875
frequency|1876,1885
,|1885,1886
urgency|1887,1894
,|1894,1895
dysuria|1896,1903
,|1903,1904
<EOL>|1905,1906
lightheadedness|1906,1921
,|1921,1922
gait|1923,1927
unsteadiness|1928,1940
,|1940,1941
focal|1942,1947
weakness|1948,1956
,|1956,1957
vision|1958,1964
<EOL>|1965,1966
changes|1966,1973
,|1973,1974
headache|1975,1983
,|1983,1984
rash|1985,1989
or|1990,1992
skin|1993,1997
changes|1998,2005
.|2005,2006
<EOL>|2008,2009
.|2009,2010
<EOL>|2012,2013
<EOL>|2013,2014
<EOL>|2015,2016
Past|2016,2020
Medical|2021,2028
History|2029,2036
:|2036,2037
<EOL>|2037,2038
CAD|2038,2041
s|2042,2043
/|2043,2044
p|2044,2045
MI|2046,2048
_|2049,2050
_|2050,2051
_|2051,2052
s|2053,2054
/|2054,2055
p|2055,2056
CABG|2057,2061
_|2062,2063
_|2063,2064
_|2064,2065
<EOL>|2065,2066
Hypertension|2066,2078
<EOL>|2078,2079
Dyslipidemia|2079,2091
<EOL>|2091,2092
CVA|2092,2095
:|2095,2096
small|2097,2102
left|2103,2107
posterior|2108,2117
frontal|2118,2125
infarct|2126,2133
in|2134,2136
_|2137,2138
_|2138,2139
_|2139,2140
<EOL>|2140,2141
Macular|2141,2148
Degeneration|2149,2161
<EOL>|2161,2162
NSCLC|2162,2167
-|2167,2168
stage|2169,2174
IV|2175,2177
(|2178,2179
oncology|2179,2187
history|2188,2195
below|2196,2201
)|2201,2202
<EOL>|2202,2203
.|2203,2204
<EOL>|2204,2205
-|2205,2206
-|2206,2207
_|2208,2209
_|2209,2210
_|2210,2211
presented|2212,2221
in|2222,2224
with|2225,2229
unresolving|2230,2241
right|2242,2247
-|2247,2248
sided|2248,2253
pulmonary|2254,2263
<EOL>|2264,2265
infiltrate|2265,2275
and|2276,2279
an|2280,2282
unrelated|2283,2292
myocardial|2293,2303
infarction|2304,2314
.|2314,2315
<EOL>|2315,2316
-|2316,2317
-|2317,2318
_|2319,2320
_|2320,2321
_|2321,2322
Sputumcytology|2323,2337
confirmed|2338,2347
adenocarcinoma|2348,2362
with|2363,2367
a|2368,2369
<EOL>|2370,2371
pattern|2371,2378
of|2379,2381
stainpositivity|2382,2397
consistent|2398,2408
with|2409,2413
lung|2414,2418
origin|2419,2425
(|2426,2427
CK7|2427,2430
and|2431,2434
<EOL>|2435,2436
TTF|2436,2439
-|2439,2440
1|2440,2441
positive|2442,2450
)|2450,2451
.|2451,2452
She|2453,2456
had|2457,2460
stage|2461,2466
IV|2467,2469
nonsmall|2470,2478
cell|2479,2483
lung|2484,2488
cancer|2489,2495
,|2495,2496
<EOL>|2497,2498
based|2498,2503
on|2504,2506
the|2507,2510
multiple|2511,2519
intrapulmonary|2520,2534
lesions|2535,2542
.|2542,2543
She|2544,2547
has|2548,2551
no|2552,2554
<EOL>|2555,2556
evidence|2556,2564
of|2565,2567
extrathoracic|2568,2581
or|2582,2584
central|2585,2592
nervous|2593,2600
system|2601,2607
involvement|2608,2619
<EOL>|2620,2621
with|2621,2625
metastasis|2626,2636
.|2636,2637
<EOL>|2637,2638
-|2638,2639
-|2639,2640
_|2641,2642
_|2642,2643
_|2643,2644
:|2644,2645
Status|2646,2652
post|2653,2657
6|2658,2659
cycles|2660,2666
of|2667,2669
pemetrexed|2670,2680
<EOL>|2681,2682
500|2682,2685
-|2685,2686
>|2686,2687
400|2687,2690
>|2690,2691
200|2691,2694
mg|2695,2697
/|2697,2698
m2|2698,2700
on|2701,2703
_|2704,2705
_|2705,2706
_|2706,2707
,|2707,2708
<EOL>|2709,2710
_|2710,2711
_|2711,2712
_|2712,2713
,|2713,2714
and|2715,2718
_|2719,2720
_|2720,2721
_|2721,2722
.|2722,2723
Her|2725,2728
course|2729,2735
was|2736,2739
complicated|2740,2751
by|2752,2754
<EOL>|2755,2756
cytopenias|2756,2766
and|2767,2770
development|2771,2782
of|2783,2785
increased|2786,2795
creatinine|2796,2806
levels|2807,2813
.|2813,2814
<EOL>|2815,2816
-|2816,2817
-|2817,2818
_|2819,2820
_|2820,2821
_|2821,2822
Chest|2823,2828
CT|2829,2831
showed|2832,2838
partial|2839,2846
response|2847,2855
with|2856,2860
interval|2861,2869
<EOL>|2870,2871
improvement|2871,2882
in|2883,2885
the|2886,2889
consolidation|2890,2903
of|2904,2906
the|2907,2910
superior|2911,2919
segment|2920,2927
of|2928,2930
the|2931,2934
<EOL>|2935,2936
right|2936,2941
lower|2942,2947
lobe|2948,2952
and|2953,2956
nodular|2957,2964
densities|2965,2974
of|2975,2977
the|2978,2981
left|2982,2986
lower|2987,2992
lobe|2993,2997
.|2997,2998
<EOL>|3000,3001
Still|3001,3006
widely|3007,3013
disseminated|3014,3026
BAC|3027,3030
.|3030,3031
<EOL>|3032,3033
-|3033,3034
-|3034,3035
_|3036,3037
_|3037,3038
_|3038,3039
CT|3040,3042
Chest|3043,3048
shows|3049,3054
increased|3055,3064
density|3065,3072
of|3073,3075
right|3076,3081
lower|3082,3087
lobe|3088,3092
<EOL>|3092,3093
consolidation|3093,3106
and|3107,3110
worsened|3111,3119
peribronchiolar|3120,3135
ground|3136,3142
-|3142,3143
glass|3143,3148
<EOL>|3149,3150
opacities|3150,3159
<EOL>|3159,3160
in|3160,3162
the|3163,3166
lingula|3167,3174
are|3175,3178
most|3179,3183
consistent|3184,3194
with|3195,3199
worsening|3200,3209
of|3210,3212
widely|3213,3219
<EOL>|3219,3220
disseminated|3220,3232
non-small|3233,3242
cell|3243,3247
lung|3248,3252
cancer|3253,3259
,|3259,3260
much|3261,3265
less|3266,3270
likely|3271,3277
due|3278,3281
to|3282,3284
<EOL>|3284,3285
infection|3285,3294
.|3294,3295
<EOL>|3296,3297
-|3297,3298
-|3298,3299
_|3300,3301
_|3301,3302
_|3302,3303
Chest|3304,3309
CT|3310,3312
:|3312,3313
slight|3314,3320
interval|3321,3329
progression|3330,3341
of|3342,3344
known|3345,3350
<EOL>|3351,3352
disease|3352,3359
,|3359,3360
no|3361,3363
new|3364,3367
sites|3368,3373
.|3373,3374
<EOL>|3374,3375
<EOL>|3375,3376
<EOL>|3377,3378
Social|3378,3384
History|3385,3392
:|3392,3393
<EOL>|3393,3394
_|3394,3395
_|3395,3396
_|3396,3397
<EOL>|3397,3398
Family|3398,3404
History|3405,3412
:|3412,3413
<EOL>|3413,3414
Her|3414,3417
father|3418,3424
died|3425,3429
due|3430,3433
to|3434,3436
CAD|3437,3440
at|3441,3443
age|3444,3447
_|3448,3449
_|3449,3450
_|3450,3451
.|3451,3452
Her|3453,3456
mother|3457,3463
had|3464,3467
stomach|3468,3475
<EOL>|3476,3477
cancer|3477,3483
and|3484,3487
osteosarcoma|3488,3500
.|3500,3501
No|3502,3504
history|3505,3512
of|3513,3515
lung|3516,3520
cancer|3521,3527
,|3527,3528
colon|3529,3534
cancer|3535,3541
<EOL>|3542,3543
or|3543,3545
breast|3546,3552
cancer|3553,3559
.|3559,3560
<EOL>|3560,3561
<EOL>|3562,3563
Physical|3563,3571
Exam|3572,3576
:|3576,3577
<EOL>|3577,3578
On|3578,3580
Admission|3581,3590
:|3590,3591
<EOL>|3591,3592
Vitals|3592,3598
:|3598,3599
T|3600,3601
:|3601,3602
96.9|3603,3607
BP|3608,3610
:|3610,3611
118|3612,3615
/|3615,3616
51|3616,3618
HR|3619,3621
:|3621,3622
94|3623,3625
RR|3626,3628
:|3628,3629
18|3630,3632
O2Sat|3633,3638
:|3638,3639
94|3640,3642
%|3642,3643
on|3644,3646
5L|3647,3649
with|3650,3654
<EOL>|3655,3656
face|3656,3660
tent|3661,3665
<EOL>|3667,3668
GEN|3668,3671
:|3671,3672
Well|3673,3677
-|3677,3678
appearing|3678,3687
female|3688,3694
in|3695,3697
no|3698,3700
acute|3701,3706
distress|3707,3715
<EOL>|3717,3718
HEENT|3718,3723
:|3723,3724
EOMI|3725,3729
,|3729,3730
PERRL|3731,3736
,|3736,3737
sclera|3738,3744
anicteric|3745,3754
,|3754,3755
MMM|3756,3759
,|3759,3760
OP|3761,3763
Clear|3764,3769
<EOL>|3771,3772
NECK|3772,3776
:|3776,3777
No|3778,3780
JVD|3781,3784
,|3784,3785
no|3786,3788
cervical|3789,3797
lymphadenopathy|3798,3813
,|3813,3814
trachea|3815,3822
midline|3823,3830
<EOL>|3832,3833
COR|3833,3836
:|3836,3837
Regular|3838,3845
rate|3846,3850
and|3851,3854
rhythm|3855,3861
,|3861,3862
no|3863,3865
M|3866,3867
/|3867,3868
G|3868,3869
/|3869,3870
R|3870,3871
,|3871,3872
normal|3873,3879
S1|3880,3882
S2|3883,3885
<EOL>|3885,3886
PULM|3886,3890
:|3890,3891
Decreased|3892,3901
breath|3902,3908
sounds|3909,3915
throughout|3916,3926
.|3926,3927
minimally|3929,3938
faint|3939,3944
<EOL>|3945,3946
bibasilar|3946,3955
crackles|3956,3964
.|3964,3965
Good|3967,3971
effort|3972,3978
.|3978,3979
<EOL>|3983,3984
ABD|3984,3987
:|3987,3988
Soft|3989,3993
,|3993,3994
NT|3995,3997
,|3997,3998
ND|3999,4001
,|4001,4002
+|4003,4004
BS|4004,4006
,|4006,4007
no|4008,4010
HSM|4011,4014
,|4014,4015
<EOL>|4015,4016
EXT|4016,4019
:|4019,4020
No|4021,4023
C|4024,4025
/|4025,4026
C|4026,4027
/|4027,4028
E|4028,4029
<EOL>|4031,4032
NEURO|4032,4037
:|4037,4038
alert|4039,4044
,|4044,4045
oriented|4046,4054
to|4055,4057
person|4058,4064
,|4064,4065
place|4066,4071
,|4071,4072
and|4073,4076
time|4077,4081
.|4081,4082
CN|4083,4085
II|4086,4088
|4089,4090
XII|4091,4094
<EOL>|4095,4096
grossly|4096,4103
intact|4104,4110
.|4110,4111
Moves|4112,4117
all|4118,4121
4|4122,4123
extremities|4124,4135
.|4135,4136
<EOL>|4138,4139
SKIN|4139,4143
:|4143,4144
No|4145,4147
jaundice|4148,4156
,|4156,4157
cyanosis|4158,4166
,|4166,4167
or|4168,4170
gross|4171,4176
dermatitis|4177,4187
.|4187,4188
No|4189,4191
ecchymoses|4192,4202
.|4202,4203
<EOL>|4204,4205
<EOL>|4206,4207
.|4207,4208
<EOL>|4210,4211
<EOL>|4211,4212
<EOL>|4213,4214
Pertinent|4214,4223
Results|4224,4231
:|4231,4232
<EOL>|4232,4233
_|4233,4234
_|4234,4235
_|4235,4236
08|4237,4239
:|4239,4240
30PM|4240,4244
WBC|4247,4250
-|4250,4251
17|4251,4253
.|4253,4254
9|4254,4255
*|4255,4256
#|4256,4257
RBC|4258,4261
-|4261,4262
3|4262,4263
.|4263,4264
36|4264,4266
*|4266,4267
#|4267,4268
HGB|4269,4272
-|4272,4273
8|4273,4274
.|4274,4275
1|4275,4276
*|4276,4277
HCT|4278,4281
-|4281,4282
25|4282,4284
.|4284,4285
5|4285,4286
*|4286,4287
<EOL>|4288,4289
MCV|4289,4292
-|4292,4293
76|4293,4295
*|4295,4296
MCH|4297,4300
-|4300,4301
24|4301,4303
.|4303,4304
2|4304,4305
*|4305,4306
MCHC|4307,4311
-|4311,4312
31.8|4312,4316
RDW|4317,4320
-|4320,4321
15|4321,4323
.|4323,4324
8|4324,4325
*|4325,4326
<EOL>|4326,4327
_|4327,4328
_|4328,4329
_|4329,4330
08|4331,4333
:|4333,4334
30PM|4334,4338
PLT|4341,4344
COUNT|4345,4350
-|4350,4351
341|4351,4354
<EOL>|4354,4355
_|4355,4356
_|4356,4357
_|4357,4358
08|4359,4361
:|4361,4362
30PM|4362,4366
NEUTS|4369,4374
-|4374,4375
84|4375,4377
*|4377,4378
BANDS|4379,4384
-|4384,4385
7|4385,4386
*|4386,4387
LYMPHS|4388,4394
-|4394,4395
2|4395,4396
*|4396,4397
MONOS|4398,4403
-|4403,4404
7|4404,4405
EOS|4406,4409
-|4409,4410
0|4410,4411
<EOL>|4412,4413
BASOS|4413,4418
-|4418,4419
0|4419,4420
_|4421,4422
_|4422,4423
_|4423,4424
MYELOS|4425,4431
-|4431,4432
0|4432,4433
<EOL>|4433,4434
_|4434,4435
_|4435,4436
_|4436,4437
08|4438,4440
:|4440,4441
30PM|4441,4445
HYPOCHROM|4448,4457
-|4457,4458
3|4458,4459
+|4459,4460
ANISOCYT|4461,4469
-|4469,4470
1|4470,4471
+|4471,4472
POIKILOCY|4473,4482
-|4482,4483
NORMAL|4483,4489
<EOL>|4490,4491
MACROCYT|4491,4499
-|4499,4500
1|4500,4501
+|4501,4502
MICROCYT|4503,4511
-|4511,4512
2|4512,4513
+|4513,4514
POLYCHROM|4515,4524
-|4524,4525
1|4525,4526
+|4526,4527
OVALOCYT|4528,4536
-|4536,4537
1|4537,4538
+|4538,4539
TEARDROP|4540,4548
-|4548,4549
1|4549,4550
+|4550,4551
<EOL>|4552,4553
ENVELOP|4553,4560
-|4560,4561
1|4561,4562
+|4562,4563
<EOL>|4563,4564
_|4564,4565
_|4565,4566
_|4566,4567
08|4568,4570
:|4570,4571
30PM|4571,4575
_|4578,4579
_|4579,4580
_|4580,4581
PTT|4582,4585
-|4585,4586
26.5|4586,4590
_|4591,4592
_|4592,4593
_|4593,4594
<EOL>|4594,4595
_|4595,4596
_|4596,4597
_|4597,4598
08|4599,4601
:|4601,4602
30PM|4602,4606
GLUCOSE|4609,4616
-|4616,4617
117|4617,4620
*|4620,4621
UREA|4622,4626
N|4627,4628
-|4628,4629
71|4629,4631
*|4631,4632
CREAT|4633,4638
-|4638,4639
2|4639,4640
.|4640,4641
8|4641,4642
*|4642,4643
SODIUM|4644,4650
-|4650,4651
135|4651,4654
<EOL>|4655,4656
POTASSIUM|4656,4665
-|4665,4666
4.9|4666,4669
CHLORIDE|4670,4678
-|4678,4679
98|4679,4681
TOTAL|4682,4687
CO2|4688,4691
-|4691,4692
23|4692,4694
ANION|4695,4700
GAP|4701,4704
-|4704,4705
19|4705,4707
<EOL>|4707,4708
_|4708,4709
_|4709,4710
_|4710,4711
08|4712,4714
:|4714,4715
43PM|4715,4719
LACTATE|4722,4729
-|4729,4730
2|4730,4731
.|4731,4732
6|4732,4733
*|4733,4734
<EOL>|4734,4735
_|4735,4736
_|4736,4737
_|4737,4738
08|4739,4741
:|4741,4742
30PM|4742,4746
cTropnT|4749,4756
-|4756,4757
<|4757,4758
0|4758,4759
.|4759,4760
01|4760,4762
<EOL>|4762,4763
_|4763,4764
_|4764,4765
_|4765,4766
10|4767,4769
:|4769,4770
46PM|4770,4774
URINE|4775,4780
COLOR|4782,4787
-|4787,4788
Straw|4788,4793
APPEAR|4794,4800
-|4800,4801
Clear|4801,4806
SP|4807,4809
_|4810,4811
_|4811,4812
_|4812,4813
<EOL>|4813,4814
_|4814,4815
_|4815,4816
_|4816,4817
10|4818,4820
:|4820,4821
46PM|4821,4825
URINE|4826,4831
BLOOD|4833,4838
-|4838,4839
NEG|4839,4842
NITRITE|4843,4850
-|4850,4851
NEG|4851,4854
PROTEIN|4855,4862
-|4862,4863
NEG|4863,4866
<EOL>|4867,4868
GLUCOSE|4868,4875
-|4875,4876
NEG|4876,4879
KETONE|4880,4886
-|4886,4887
NEG|4887,4890
BILIRUBIN|4891,4900
-|4900,4901
NEG|4901,4904
UROBILNGN|4905,4914
-|4914,4915
NEG|4915,4918
PH|4919,4921
-|4921,4922
5.0|4922,4925
<EOL>|4926,4927
LEUK|4927,4931
-|4931,4932
NEG|4932,4935
<EOL>|4935,4936
.|4936,4937
<EOL>|4937,4938
Micro|4938,4943
:|4943,4944
<EOL>|4944,4945
Legionella|4945,4955
Urinary|4956,4963
Antigen|4964,4971
(|4973,4974
Final|4974,4979
_|4980,4981
_|4981,4982
_|4982,4983
:|4983,4984
<EOL>|4985,4986
NEGATIVE|4992,5000
FOR|5001,5004
LEGIONELLA|5005,5015
SEROGROUP|5016,5025
1|5026,5027
ANTIGEN|5028,5035
<EOL>|5035,5036
.|5036,5037
<EOL>|5037,5038
Urine|5038,5043
cx|5044,5046
:|5046,5047
URINE|5050,5055
CULTURE|5056,5063
(|5064,5065
Final|5065,5070
_|5071,5072
_|5072,5073
_|5073,5074
:|5074,5075
NO|5079,5081
GROWTH|5082,5088
.|5088,5089
<EOL>|5089,5090
<EOL>|5090,5091
Blood|5091,5096
cx|5097,5099
:|5099,5100
NGTD|5101,5105
<EOL>|5105,5106
.|5106,5107
<EOL>|5107,5108
Studies|5108,5115
/|5115,5116
Imaging|5116,5123
:|5123,5124
<EOL>|5124,5125
.|5125,5126
<EOL>|5126,5127
EKG|5127,5130
:|5130,5131
_|5132,5133
_|5133,5134
_|5134,5135
<EOL>|5135,5136
Sinus|5136,5141
rhythm|5142,5148
at|5149,5151
68|5152,5154
bpm|5155,5158
,|5158,5159
normal|5160,5166
axis|5167,5171
,|5171,5172
normal|5173,5179
intervals|5180,5189
,|5189,5190
poor|5191,5195
<EOL>|5196,5197
R|5197,5198
-|5198,5199
wave|5199,5203
progresion|5204,5214
,|5214,5215
ST|5216,5218
-|5218,5219
depressions|5219,5230
in|5231,5233
V4|5234,5236
-|5236,5237
V6|5237,5239
.|5239,5240
<EOL>|5240,5241
.|5241,5242
<EOL>|5242,5243
CXR|5243,5246
:|5246,5247
_|5248,5249
_|5249,5250
_|5250,5251
<EOL>|5251,5252
SINGLE|5252,5258
AP|5259,5261
VIEW|5262,5266
OF|5267,5269
THE|5270,5273
CHEST|5274,5279
:|5279,5280
Patient|5281,5288
is|5289,5291
status|5292,5298
post|5299,5303
median|5304,5310
<EOL>|5311,5312
sternotomy|5312,5322
.|5322,5323
The|5324,5327
<EOL>|5328,5329
cardiac|5329,5336
,|5336,5337
mediastinal|5338,5349
and|5350,5353
hilar|5354,5359
contours|5360,5368
are|5369,5372
unchanged|5373,5382
.|5382,5383
There|5384,5389
<EOL>|5390,5391
continues|5391,5400
to|5401,5403
be|5404,5406
progression|5407,5418
of|5419,5421
disease|5422,5429
with|5430,5434
increased|5435,5444
extent|5445,5451
of|5452,5454
<EOL>|5455,5456
consolidative|5456,5469
opacity|5470,5477
within|5478,5484
the|5485,5488
right|5489,5494
lung|5495,5499
base|5500,5504
.|5504,5505
Ill|5506,5509
-|5509,5510
defined|5510,5517
<EOL>|5518,5519
opacities|5519,5528
within|5529,5535
the|5536,5539
lingula|5540,5547
and|5548,5551
left|5552,5556
lower|5557,5562
lobe|5563,5567
are|5568,5571
similar|5572,5579
to|5580,5582
<EOL>|5583,5584
prior|5584,5589
.|5589,5590
Small|5591,5596
right|5597,5602
pleural|5603,5610
effusion|5611,5619
is|5620,5622
present|5623,5630
.|5630,5631
There|5632,5637
is|5638,5640
no|5641,5643
<EOL>|5644,5645
pneumothorax|5645,5657
.|5657,5658
There|5659,5664
is|5665,5667
hyperinflation|5668,5682
of|5683,5685
the|5686,5689
lungs|5690,5695
.|5695,5696
<EOL>|5697,5698
IMPRESSION|5698,5708
:|5708,5709
Evidence|5710,5718
of|5719,5721
disease|5722,5729
progression|5730,5741
.|5741,5742
<EOL>|5743,5744
.|5744,5745
<EOL>|5745,5746
CT|5746,5748
Head|5749,5753
:|5753,5754
_|5755,5756
_|5756,5757
_|5757,5758
<EOL>|5758,5759
FINDINGS|5759,5767
:|5767,5768
There|5769,5774
is|5775,5777
no|5778,5780
evidence|5781,5789
of|5790,5792
acute|5793,5798
hemorrhage|5799,5809
,|5809,5810
edema|5811,5816
,|5816,5817
mass|5818,5822
<EOL>|5823,5824
effect|5824,5830
or|5831,5833
<EOL>|5834,5835
recent|5835,5841
infarction|5842,5852
.|5852,5853
An|5854,5856
area|5857,5861
of|5862,5864
encephalomalacia|5865,5881
in|5882,5884
the|5885,5888
left|5889,5893
<EOL>|5894,5895
frontal|5895,5902
lobe|5903,5907
,|5907,5908
<EOL>|5909,5910
compatible|5910,5920
with|5921,5925
chronic|5926,5933
infarct|5934,5941
is|5942,5944
unchanged|5945,5954
.|5954,5955
Prominence|5956,5966
of|5967,5969
the|5970,5973
<EOL>|5974,5975
ventricles|5975,5985
<EOL>|5986,5987
and|5987,5990
sulci|5991,5996
reflects|5997,6005
generalized|6006,6017
atrophy|6018,6025
,|6025,6026
notably|6027,6034
in|6035,6037
the|6038,6041
bifrontal|6042,6051
<EOL>|6052,6053
extraaxial|6053,6063
spaces|6064,6070
.|6070,6071
Areas|6072,6077
of|6078,6080
periventricular|6081,6096
and|6097,6100
subcortical|6101,6112
<EOL>|6113,6114
white|6114,6119
matter|6120,6126
hypodensity|6127,6138
likely|6139,6145
reflect|6146,6153
sequela|6154,6161
of|6162,6164
chronic|6165,6172
small|6173,6178
<EOL>|6179,6180
vessel|6180,6186
ischemic|6187,6195
disease|6196,6203
.|6203,6204
No|6205,6207
concerning|6208,6218
osseous|6219,6226
lesion|6227,6233
is|6234,6236
seen|6237,6241
.|6241,6242
<EOL>|6243,6244
There|6244,6249
are|6250,6253
calcifications|6254,6268
of|6269,6271
the|6272,6275
bilateral|6276,6285
carotid|6286,6293
siphons|6294,6301
.|6301,6302
The|6303,6306
<EOL>|6307,6308
visualized|6308,6318
paranasal|6319,6328
sinuses|6329,6336
are|6337,6340
grossly|6341,6348
unremarkable|6349,6361
.|6361,6362
<EOL>|6363,6364
IMPRESSION|6364,6374
:|6374,6375
No|6376,6378
evidence|6379,6387
of|6388,6390
acute|6391,6396
intracranial|6397,6409
process|6410,6417
or|6418,6420
mass|6421,6425
<EOL>|6426,6427
effect|6427,6433
<EOL>|6434,6435
.|6435,6436
<EOL>|6436,6437
LENIs|6437,6442
:|6442,6443
_|6444,6445
_|6445,6446
_|6446,6447
<EOL>|6447,6448
IMPRESSION|6448,6458
:|6458,6459
No|6460,6462
evidence|6463,6471
of|6472,6474
DVT|6475,6478
.|6478,6479
<EOL>|6480,6481
.|6481,6482
<EOL>|6482,6483
CT|6483,6485
chest|6486,6491
_|6492,6493
_|6493,6494
_|6494,6495
<EOL>|6495,6496
IMPRESSION|6496,6506
:|6506,6507
<EOL>|6509,6510
1.|6510,6512
Interval|6513,6521
worsening|6522,6531
of|6532,6534
diffuse|6535,6542
bilateral|6543,6552
ground|6553,6559
-|6559,6560
glass|6560,6565
<EOL>|6566,6567
opacities|6567,6576
,|6576,6577
<EOL>|6578,6579
bronchiolar|6579,6590
nodules|6591,6598
and|6599,6602
dense|6603,6608
consolidation|6609,6622
within|6623,6629
the|6630,6633
lingula|6634,6641
<EOL>|6642,6643
and|6643,6646
right|6647,6652
<EOL>|6653,6654
middle|6654,6660
lobe|6661,6665
.|6665,6666
After|6667,6672
review|6673,6679
of|6680,6682
multiple|6683,6691
recent|6692,6698
prior|6699,6704
chest|6705,6710
x-rays|6711,6717
<EOL>|6718,6719
and|6719,6722
CTs|6723,6726
,|6726,6727
these|6728,6733
findings|6734,6742
can|6743,6746
all|6747,6750
be|6751,6753
explained|6754,6763
by|6764,6766
worsening|6767,6776
<EOL>|6777,6778
bronchioalveolar|6778,6794
carcinoma|6795,6804
,|6804,6805
given|6806,6811
the|6812,6815
absence|6816,6823
of|6824,6826
any|6827,6830
change|6831,6837
<EOL>|6838,6839
rapid|6839,6844
enough|6845,6851
to|6852,6854
suggest|6855,6862
pneumonia|6863,6872
.|6872,6873
Of|6874,6876
course|6877,6883
pneumonia|6884,6893
might|6894,6899
be|6900,6902
<EOL>|6903,6904
present|6904,6911
and|6912,6915
unrecognized|6916,6928
,|6928,6929
and|6930,6933
treatment|6934,6943
should|6944,6950
be|6951,6953
made|6954,6958
on|6959,6961
the|6962,6965
<EOL>|6966,6967
basis|6967,6972
of|6973,6975
clinical|6976,6984
findings|6985,6993
.|6993,6994
<EOL>|6995,6996
2.|6996,6998
Stable|6999,7005
mild|7006,7010
cardiomegaly|7011,7023
.|7023,7024
<EOL>|7025,7026
3.|7026,7028
Moderate|7029,7037
emphysema|7038,7047
.|7047,7048
<EOL>|7049,7050
4.|7050,7052
Cholelithiasis|7053,7067
without|7068,7075
evidence|7076,7084
of|7085,7087
cholecystitis|7088,7101
.|7101,7102
<EOL>|7103,7104
<EOL>|7104,7105
<EOL>|7106,7107
Brief|7107,7112
Hospital|7113,7121
Course|7122,7128
:|7128,7129
<EOL>|7129,7130
_|7130,7131
_|7131,7132
_|7132,7133
female|7134,7140
with|7141,7145
NSCLC|7146,7151
stage|7152,7157
IV|7158,7160
presents|7161,7169
with|7170,7174
hypoxia|7175,7182
.|7182,7183
<EOL>|7183,7184
.|7184,7185
<EOL>|7185,7186
#|7186,7187
.|7187,7188
Hypoxia|7189,7196
.|7196,7197
On|7198,7200
admission|7201,7210
patient|7211,7218
with|7219,7223
chief|7224,7229
complaints|7230,7240
of|7241,7243
<EOL>|7244,7245
progressive|7245,7256
shortness|7257,7266
of|7267,7269
breath|7270,7276
and|7277,7280
non-productive|7281,7295
cough|7296,7301
.|7301,7302
No|7303,7305
<EOL>|7306,7307
home|7307,7311
oxygen|7312,7318
requirement|7319,7330
at|7331,7333
baseline|7334,7342
.|7342,7343
On|7344,7346
admission|7347,7356
she|7357,7360
was|7361,7364
placed|7365,7371
<EOL>|7372,7373
on|7373,7375
NRB|7376,7379
for|7380,7383
treatment|7384,7393
of|7394,7396
O2|7397,7399
saturations|7400,7411
in|7412,7414
_|7415,7416
_|7416,7417
_|7417,7418
saturations|7419,7430
in|7431,7433
the|7434,7437
<EOL>|7438,7439
_|7439,7440
_|7440,7441
_|7441,7442
.|7442,7443
Admission|7445,7454
CXR|7455,7458
with|7459,7463
no|7464,7466
definite|7467,7475
infiltrate|7476,7486
,|7486,7487
though|7488,7494
concern|7495,7502
<EOL>|7503,7504
for|7504,7507
progression|7508,7519
of|7520,7522
her|7523,7526
known|7527,7532
lung|7533,7537
disease|7538,7545
.|7545,7546
In|7547,7549
setting|7550,7557
of|7558,7560
<EOL>|7561,7562
elevated|7562,7570
WBC|7571,7574
.|7574,7575
concern|7576,7583
for|7584,7587
infectious|7588,7598
process|7599,7606
and|7607,7610
empirically|7611,7622
<EOL>|7623,7624
treated|7624,7631
with|7632,7636
levofloxacin|7637,7649
and|7650,7653
vancomycin|7654,7664
in|7665,7667
the|7668,7671
ED|7672,7674
.|7674,7675
Transitioned|7676,7688
<EOL>|7689,7690
to|7690,7692
monotherapy|7693,7704
with|7705,7709
levofloxacin|7710,7722
on|7723,7725
_|7726,7727
_|7727,7728
_|7728,7729
and|7730,7733
ceftriaxone|7734,7745
was|7746,7749
<EOL>|7750,7751
later|7751,7756
added|7757,7762
on|7763,7765
_|7766,7767
_|7767,7768
_|7768,7769
.|7769,7770
CXR|7771,7774
on|7775,7777
_|7778,7779
_|7779,7780
_|7780,7781
demonstrates|7782,7794
new|7795,7798
left|7799,7803
lower|7804,7809
<EOL>|7810,7811
lobe|7811,7815
consolidation|7816,7829
.|7829,7830
Additional|7831,7841
hypoxia|7842,7849
work|7850,7854
-|7854,7855
up|7855,7857
notable|7858,7865
for|7866,7869
<EOL>|7870,7871
negative|7871,7879
biomarkers|7880,7890
,|7890,7891
negative|7892,7900
LENIs|7901,7906
;|7906,7907
unable|7908,7914
to|7915,7917
perform|7918,7925
CTA|7926,7929
due|7930,7933
<EOL>|7934,7935
to|7935,7937
chronic|7938,7945
kidney|7946,7952
disease|7953,7960
and|7961,7964
creatinine|7965,7975
2.8|7976,7979
.|7979,7980
Patient|7981,7988
was|7989,7992
able|7993,7997
<EOL>|7998,7999
to|7999,8001
be|8002,8004
weaned|8005,8011
back|8012,8016
to|8017,8019
room|8020,8024
air|8025,8028
by|8029,8031
the|8032,8035
end|8036,8039
of|8040,8042
her|8043,8046
FICU|8047,8051
stay|8052,8056
.|8056,8057
She|8058,8061
<EOL>|8062,8063
was|8063,8066
transferred|8067,8078
to|8079,8081
the|8082,8085
medical|8086,8093
floor|8094,8099
on|8100,8102
_|8103,8104
_|8104,8105
_|8105,8106
,|8106,8107
where|8108,8113
she|8114,8117
<EOL>|8118,8119
demonstrated|8119,8131
exertional|8132,8142
hypoxia|8143,8150
,|8150,8151
usually|8152,8159
asymptomatic|8160,8172
.|8172,8173
Home|8174,8178
O2|8179,8181
<EOL>|8182,8183
was|8183,8186
arranged|8187,8195
.|8195,8196
<EOL>|8196,8197
.|8197,8198
<EOL>|8198,8199
#|8199,8200
Post-obstructive|8201,8217
pneumonia|8218,8227
.|8227,8228
Consolidation|8229,8242
of|8243,8245
left|8246,8250
lower|8251,8256
lobe|8257,8261
<EOL>|8262,8263
evident|8263,8270
on|8271,8273
_|8274,8275
_|8275,8276
_|8276,8277
likely|8278,8284
secondary|8285,8294
to|8295,8297
infection|8298,8307
rather|8308,8314
than|8315,8319
<EOL>|8320,8321
progression|8321,8332
of|8333,8335
disease|8336,8343
due|8344,8347
to|8348,8350
short|8351,8356
time|8357,8361
course|8362,8368
of|8369,8371
infiltrate|8372,8382
<EOL>|8383,8384
development|8384,8395
(|8396,8397
although|8397,8405
on|8406,8408
CT|8409,8411
scan|8412,8416
of|8417,8419
_|8420,8421
_|8421,8422
_|8422,8423
,|8423,8424
the|8425,8428
radiologist|8429,8440
<EOL>|8441,8442
concluded|8442,8451
the|8452,8455
opposite|8456,8464
:|8464,8465
that|8466,8470
changes|8471,8478
seen|8479,8483
were|8484,8488
likely|8489,8495
caused|8496,8502
by|8503,8505
<EOL>|8506,8507
her|8507,8510
NSCLC|8511,8516
,|8516,8517
though|8518,8524
pneumonia|8525,8534
could|8535,8540
not|8541,8544
be|8545,8547
absolutely|8548,8558
ruled|8559,8564
out|8565,8568
)|8568,8569
.|8569,8570
<EOL>|8571,8572
Continued|8572,8581
course|8582,8588
of|8589,8591
ceftriaxone|8592,8603
,|8603,8604
levofloxacin|8605,8617
,|8617,8618
which|8619,8624
was|8625,8628
<EOL>|8629,8630
eventually|8630,8640
narrowed|8641,8649
to|8650,8652
levofloxacin|8653,8665
alone|8666,8671
.|8671,8672
Blood|8673,8678
cultures|8679,8687
no|8688,8690
<EOL>|8691,8692
growth|8692,8698
to|8699,8701
date|8702,8706
.|8706,8707
Multiple|8708,8716
sputum|8717,8723
cultures|8724,8732
obtained|8733,8741
;|8741,8742
however|8743,8750
,|8750,8751
all|8752,8755
<EOL>|8756,8757
contaminated|8757,8769
with|8770,8774
oral|8775,8779
flora|8780,8785
.|8785,8786
Urine|8787,8792
legionella|8793,8803
negative|8804,8812
.|8812,8813
Patient|8814,8821
<EOL>|8822,8823
did|8823,8826
improve|8827,8834
clinically|8835,8845
with|8846,8850
antibiotics|8851,8862
,|8862,8863
so|8864,8866
she|8867,8870
should|8871,8877
complete|8878,8886
<EOL>|8887,8888
a|8888,8889
_|8890,8891
_|8891,8892
_|8892,8893
day|8894,8897
course|8898,8904
of|8905,8907
levofloxacin|8908,8920
.|8920,8921
<EOL>|8921,8922
.|8922,8923
<EOL>|8923,8924
#|8924,8925
NSCLC|8927,8932
-|8932,8933
stage|8934,8939
IV|8940,8942
.|8942,8943
Not|8944,8947
currently|8948,8957
receiving|8958,8967
chemotherapy|8968,8980
.|8980,8981
<EOL>|8983,8984
Outpatient|8984,8994
oncologist|8995,9005
Dr.|9006,9009
_|9010,9011
_|9011,9012
_|9012,9013
is|9014,9016
planning|9017,9025
on|9026,9028
continued|9029,9038
<EOL>|9039,9040
surveillance|9040,9052
with|9053,9057
plan|9058,9062
for|9063,9066
possible|9067,9075
further|9076,9083
palliative|9084,9094
systemic|9095,9103
<EOL>|9104,9105
chemotherapy|9105,9117
if|9118,9120
symptomatic|9121,9132
progression|9133,9144
of|9145,9147
her|9148,9151
disease|9152,9159
is|9160,9162
noted|9163,9168
.|9168,9169
<EOL>|9170,9171
CT|9171,9173
scan|9174,9178
for|9179,9182
evaluation|9183,9193
of|9194,9196
disease|9197,9204
progression|9205,9216
was|9217,9220
obtained|9221,9229
and|9230,9233
<EOL>|9234,9235
did|9235,9238
show|9239,9243
further|9244,9251
progression|9252,9263
.|9263,9264
Dr.|9265,9268
_|9269,9270
_|9270,9271
_|9271,9272
plans|9273,9278
to|9279,9281
weigh|9282,9287
the|9288,9291
risks|9292,9297
<EOL>|9298,9299
and|9299,9302
benefits|9303,9311
of|9312,9314
additional|9315,9325
chemotherapy|9326,9338
,|9338,9339
as|9340,9342
it|9343,9345
will|9346,9350
be|9351,9353
<EOL>|9354,9355
complicated|9355,9366
by|9367,9369
her|9370,9373
kidney|9374,9380
dysfunction|9381,9392
and|9393,9396
other|9397,9402
comorbidities|9403,9416
.|9416,9417
<EOL>|9418,9419
He|9419,9421
plans|9422,9427
to|9428,9430
repeat|9431,9437
her|9438,9441
CT|9442,9444
scan|9445,9449
once|9450,9454
she|9455,9458
completes|9459,9468
her|9469,9472
<EOL>|9473,9474
antibiotics|9474,9485
to|9486,9488
further|9489,9496
evaluate|9497,9505
the|9506,9509
rate|9510,9514
of|9515,9517
disease|9518,9525
progression|9526,9537
.|9537,9538
<EOL>|9538,9539
.|9539,9540
<EOL>|9544,9545
#|9545,9546
CAD|9548,9551
s|9552,9553
/|9553,9554
p|9554,9555
MI|9556,9558
.|9558,9559
Patient|9560,9567
without|9568,9575
chest|9576,9581
pain|9582,9586
;|9586,9587
however|9588,9595
,|9595,9596
EKG|9597,9600
with|9601,9605
new|9606,9609
<EOL>|9610,9611
ST|9611,9613
-|9613,9614
depressions|9614,9625
.|9625,9626
Biomarkers|9627,9637
cycled|9638,9644
and|9645,9648
negative|9649,9657
x2|9658,9660
.|9660,9661
Patient|9662,9669
<EOL>|9670,9671
continued|9671,9680
on|9681,9683
home|9684,9688
beta|9689,9693
-|9693,9694
blocker|9694,9701
at|9702,9704
a|9705,9706
decreased|9707,9716
dose|9717,9721
due|9722,9725
to|9726,9728
<EOL>|9729,9730
relative|9730,9738
hypotension|9739,9750
.|9750,9751
She|9752,9755
was|9756,9759
maintained|9760,9770
on|9771,9773
aspirin|9774,9781
,|9781,9782
plavix|9783,9789
,|9789,9790
and|9791,9794
<EOL>|9795,9796
statin|9796,9802
.|9802,9803
<EOL>|9803,9804
.|9804,9805
<EOL>|9805,9806
#|9806,9807
chronic|9808,9815
systolic|9816,9824
CHF|9825,9828
(|9829,9830
LVEF|9830,9834
_|9835,9836
_|9836,9837
_|9837,9838
by|9839,9841
TTE|9842,9845
_|9846,9847
_|9847,9848
_|9848,9849
:|9849,9850
<EOL>|9851,9852
Well|9852,9856
-|9856,9857
compensated|9857,9868
.|9868,9869
As|9870,9872
described|9873,9882
below|9883,9888
,|9888,9889
lasix|9890,9895
was|9896,9899
held|9900,9904
but|9905,9908
<EOL>|9909,9910
B|9910,9911
-|9911,9912
blocker|9912,9919
was|9920,9923
given|9924,9929
at|9930,9932
a|9933,9934
lower|9935,9940
dose|9941,9945
given|9946,9951
relative|9952,9960
hypotension|9961,9972
<EOL>|9973,9974
and|9974,9977
exertional|9978,9988
tachycardia|9989,10000
.|10000,10001
<EOL>|10001,10002
.|10002,10003
<EOL>|10003,10004
#|10004,10005
CKD|10007,10010
stage|10011,10016
III|10017,10020
:|10020,10021
Creatinine|10022,10032
on|10033,10035
admission|10036,10045
2.8|10046,10049
,|10049,10050
down|10051,10055
to|10056,10058
2.4|10059,10062
by|10063,10065
<EOL>|10066,10067
the|10067,10070
time|10071,10075
of|10076,10078
discharge|10079,10088
.|10088,10089
She|10090,10093
was|10094,10097
given|10098,10103
minimal|10104,10111
IV|10112,10114
fluids|10115,10121
in|10122,10124
the|10125,10128
<EOL>|10129,10130
ICU|10130,10133
and|10134,10137
her|10138,10141
lasix|10142,10147
was|10148,10151
held|10152,10156
.|10156,10157
Throughout|10158,10168
stay|10169,10173
,|10173,10174
patient|10175,10182
had|10183,10186
<EOL>|10187,10188
adequate|10188,10196
urine|10197,10202
output|10203,10209
.|10209,10210
<EOL>|10211,10212
.|10212,10213
<EOL>|10213,10214
#|10214,10215
Microcytic|10217,10227
anemia|10228,10234
.|10234,10235
On|10236,10238
presentation|10239,10251
,|10251,10252
patient|10253,10260
's|10260,10262
Hct|10263,10266
likely|10267,10273
<EOL>|10274,10275
hemoconcentrated|10275,10291
.|10291,10292
Follow|10293,10299
-|10299,10300
up|10300,10302
Hct|10303,10306
found|10307,10312
to|10313,10315
be|10316,10318
20|10319,10321
.|10321,10322
No|10323,10325
signs|10326,10331
of|10332,10334
<EOL>|10335,10336
bleeding|10336,10344
on|10345,10347
exam|10348,10352
.|10352,10353
Patient|10354,10361
transfused|10362,10372
2units|10373,10379
of|10380,10382
pRBC|10383,10387
due|10388,10391
to|10392,10394
<EOL>|10395,10396
history|10396,10403
of|10404,10406
CAD|10407,10410
with|10411,10415
appropriate|10416,10427
elevation|10428,10437
in|10438,10440
hematocrit|10441,10451
.|10451,10452
The|10453,10456
<EOL>|10457,10458
hematocrit|10458,10468
did|10469,10472
remain|10473,10479
steady|10480,10486
during|10487,10493
FICU|10494,10498
course|10499,10505
following|10506,10515
<EOL>|10516,10517
tranfusion|10517,10527
.|10527,10528
Just|10529,10533
before|10534,10540
transfer|10541,10549
from|10550,10554
_|10555,10556
_|10556,10557
_|10557,10558
,|10558,10559
the|10560,10563
patient|10564,10571
's|10571,10573
stool|10574,10579
<EOL>|10580,10581
guaiac|10581,10587
was|10588,10591
positive|10592,10600
,|10600,10601
which|10602,10607
may|10608,10611
call|10612,10616
for|10617,10620
further|10621,10628
work|10629,10633
-|10633,10634
up|10634,10636
.|10636,10637
The|10638,10641
<EOL>|10642,10643
patient|10643,10650
's|10650,10652
anemia|10653,10659
is|10660,10662
most|10663,10667
likely|10668,10674
secondary|10675,10684
to|10685,10687
acute|10688,10693
inflammation|10694,10706
<EOL>|10707,10708
in|10708,10710
the|10711,10714
setting|10715,10722
of|10723,10725
underlying|10726,10736
chronic|10737,10744
disease|10745,10752
.|10752,10753
<EOL>|10754,10755
.|10755,10756
<EOL>|10756,10757
<EOL>|10758,10759
Medications|10759,10770
on|10771,10773
Admission|10774,10783
:|10783,10784
<EOL>|10784,10785
amlodipine|10785,10795
5|10796,10797
mg|10798,10800
Tablet|10801,10807
-|10807,10808
one|10809,10812
Tablet|10813,10819
(|10819,10820
s|10820,10821
)|10821,10822
by|10823,10825
mouth|10826,10831
one|10832,10835
daily|10836,10841
<EOL>|10843,10844
atorvastatin|10844,10856
[|10857,10858
Lipitor|10858,10865
]|10865,10866
80|10867,10869
mg|10870,10872
Tablet|10873,10879
-|10879,10880
one|10881,10884
Tablet|10885,10891
(|10891,10892
s|10892,10893
)|10893,10894
by|10895,10897
mouth|10898,10903
one|10904,10907
<EOL>|10908,10909
daily|10909,10914
<EOL>|10915,10916
calcitriol|10916,10926
0.25|10927,10931
mcg|10932,10935
Capsule|10936,10943
-|10943,10944
1|10945,10946
Capsule|10947,10954
(|10954,10955
s|10955,10956
)|10956,10957
by|10958,10960
mouth|10961,10966
once|10967,10971
a|10972,10973
day|10974,10977
<EOL>|10977,10978
clopidogrel|10978,10989
[|10990,10991
Plavix|10991,10997
]|10997,10998
75|10999,11001
mg|11002,11004
Tablet|11005,11011
1|11012,11013
Tablet|11014,11020
(|11020,11021
s|11021,11022
)|11022,11023
by|11024,11026
mouth|11027,11032
once|11033,11037
a|11038,11039
<EOL>|11040,11041
day|11041,11044
<EOL>|11045,11046
folic|11046,11051
acid|11052,11056
-|11056,11057
1|11058,11059
mg|11060,11062
Tablet|11063,11069
one|11070,11073
Tablet|11074,11080
(|11080,11081
s|11081,11082
)|11082,11083
by|11084,11086
mouth|11087,11092
one|11093,11096
daily|11097,11102
<EOL>|11103,11104
furosemide|11104,11114
40|11115,11117
mg|11118,11120
Tablet|11121,11127
-|11127,11128
1|11129,11130
Tablet|11131,11137
(|11137,11138
s|11138,11139
)|11139,11140
by|11141,11143
mouth|11144,11149
daily|11150,11155
<EOL>|11155,11156
loperamide|11156,11166
2|11167,11168
mg|11169,11171
Capsule|11172,11179
-|11179,11180
one|11181,11184
Capsule|11185,11192
(|11192,11193
s|11193,11194
)|11194,11195
by|11196,11198
mouth|11199,11204
one|11205,11208
twice|11209,11214
daily|11215,11220
<EOL>|11221,11222
as|11222,11224
needed|11225,11231
<EOL>|11232,11233
lorazepam|11233,11242
0.5|11243,11246
mg|11247,11249
Tablet|11250,11256
_|11257,11258
_|11258,11259
_|11259,11260
Tablet|11261,11267
(|11267,11268
s|11268,11269
)|11269,11270
by|11271,11273
mouth|11274,11279
q6|11280,11282
hours|11283,11288
as|11289,11291
<EOL>|11292,11293
needed|11293,11299
for|11300,11303
Nausea|11304,11310
<EOL>|11311,11312
metoprolol|11312,11322
tartrate|11323,11331
[|11332,11333
Lopressor|11333,11342
]|11342,11343
50|11344,11346
mg|11347,11349
Tablet|11350,11356
-|11356,11357
one|11358,11361
Tablet|11362,11368
(|11368,11369
s|11369,11370
)|11370,11371
by|11372,11374
<EOL>|11375,11376
mouth|11376,11381
_|11382,11383
_|11383,11384
_|11384,11385
AM|11386,11388
and|11389,11392
one|11393,11396
in|11397,11399
_|11400,11401
_|11401,11402
_|11402,11403
<EOL>|11404,11405
tramadol|11405,11413
50|11414,11416
mg|11417,11419
Tablet|11420,11426
-|11426,11427
0.5|11428,11431
(|11432,11433
One|11433,11436
half|11437,11441
)|11441,11442
Tablet|11443,11449
(|11449,11450
s|11450,11451
)|11451,11452
by|11453,11455
mouth|11456,11461
three|11462,11467
<EOL>|11468,11469
times|11469,11474
a|11475,11476
day|11477,11480
as|11481,11483
needed|11484,11490
for|11491,11494
Pain|11495,11499
<EOL>|11501,11502
trazodone|11502,11511
50|11512,11514
mg|11515,11517
Tablet|11518,11524
-|11524,11525
one|11526,11529
Tablet|11530,11536
(|11536,11537
s|11537,11538
)|11538,11539
by|11540,11542
mouth|11543,11548
one|11549,11552
daily|11553,11558
as|11559,11561
<EOL>|11562,11563
needed|11563,11569
<EOL>|11570,11571
aspirin|11571,11578
81|11579,11581
mg|11582,11584
Tablet|11585,11591
,|11591,11592
Chewable|11593,11601
-|11601,11602
2|11603,11604
Tablet|11605,11611
(|11611,11612
s|11612,11613
)|11613,11614
by|11615,11617
mouth|11618,11623
one|11624,11627
daily|11628,11633
<EOL>|11634,11635
ranitidine|11635,11645
HCl|11646,11649
[|11650,11651
Acid|11651,11655
Control|11656,11663
]|11663,11664
150|11665,11668
mg|11669,11671
Tablet|11672,11678
-|11678,11679
one|11680,11683
Tablet|11684,11690
(|11690,11691
s|11691,11692
)|11692,11693
by|11694,11696
<EOL>|11697,11698
mouth|11698,11703
one|11704,11707
daily|11708,11713
<EOL>|11714,11715
<EOL>|11716,11717
Discharge|11717,11726
Medications|11727,11738
:|11738,11739
<EOL>|11739,11740
1.|11740,11742
oxygen|11743,11749
<EOL>|11749,11750
_|11750,11751
_|11751,11752
_|11752,11753
continuous|11754,11764
,|11764,11765
pulse|11766,11771
dose|11772,11776
for|11777,11780
portability|11781,11792
<EOL>|11792,11793
Dx|11793,11795
:|11795,11796
lung|11797,11801
cancer|11802,11808
<EOL>|11808,11809
2.|11809,11811
levofloxacin|11812,11824
500|11825,11828
mg|11829,11831
Tablet|11832,11838
Sig|11839,11842
:|11842,11843
One|11844,11847
(|11848,11849
1|11849,11850
)|11850,11851
Tablet|11852,11858
PO|11859,11861
Q48H|11862,11866
(|11867,11868
every|11868,11873
<EOL>|11874,11875
48|11875,11877
hours|11878,11883
)|11883,11884
for|11885,11888
2|11889,11890
weeks|11891,11896
:|11896,11897
last|11898,11902
day|11903,11906
_|11907,11908
_|11908,11909
_|11909,11910
.|11910,11911
<EOL>|11911,11912
Disp|11912,11916
:|11916,11917
*|11917,11918
4|11918,11919
Tablet|11920,11926
(|11926,11927
s|11927,11928
)|11928,11929
*|11929,11930
Refills|11931,11938
:|11938,11939
*|11939,11940
0|11940,11941
*|11941,11942
<EOL>|11942,11943
3.|11943,11945
atorvastatin|11946,11958
40|11959,11961
mg|11962,11964
Tablet|11965,11971
Sig|11972,11975
:|11975,11976
Two|11977,11980
(|11981,11982
2|11982,11983
)|11983,11984
Tablet|11985,11991
PO|11992,11994
DAILY|11995,12000
<EOL>|12001,12002
(|12002,12003
Daily|12003,12008
)|12008,12009
.|12009,12010
<EOL>|12012,12013
4.|12013,12015
metoprolol|12016,12026
tartrate|12027,12035
25|12036,12038
mg|12039,12041
Tablet|12042,12048
Sig|12049,12052
:|12052,12053
One|12054,12057
(|12058,12059
1|12059,12060
)|12060,12061
Tablet|12062,12068
PO|12069,12071
twice|12072,12077
<EOL>|12078,12079
a|12079,12080
day|12081,12084
:|12084,12085
PLEASE|12086,12092
NOTE|12093,12097
THIS|12098,12102
IS|12103,12105
A|12106,12107
CHANGE|12108,12114
FROM|12115,12119
YOUR|12120,12124
PREVIOUS|12125,12133
EVENING|12134,12141
<EOL>|12142,12143
DOSING|12143,12149
.|12149,12150
<EOL>|12152,12153
5.|12153,12155
docusate|12156,12164
sodium|12165,12171
100|12172,12175
mg|12176,12178
Capsule|12179,12186
Sig|12187,12190
:|12190,12191
One|12192,12195
(|12196,12197
1|12197,12198
)|12198,12199
Capsule|12200,12207
PO|12208,12210
BID|12211,12214
(|12215,12216
2|12216,12217
<EOL>|12218,12219
times|12219,12224
a|12225,12226
day|12227,12230
)|12230,12231
:|12231,12232
hold|12233,12237
if|12238,12240
loose|12241,12246
stools|12247,12253
.|12253,12254
<EOL>|12256,12257
6.|12257,12259
trazodone|12260,12269
50|12270,12272
mg|12273,12275
Tablet|12276,12282
Sig|12283,12286
:|12286,12287
One|12288,12291
(|12292,12293
1|12293,12294
)|12294,12295
Tablet|12296,12302
PO|12303,12305
HS|12306,12308
(|12309,12310
at|12310,12312
bedtime|12313,12320
)|12320,12321
<EOL>|12322,12323
as|12323,12325
needed|12326,12332
for|12333,12336
insomnia|12337,12345
.|12345,12346
<EOL>|12348,12349
7.|12349,12351
clopidogrel|12352,12363
75|12364,12366
mg|12367,12369
Tablet|12370,12376
Sig|12377,12380
:|12380,12381
One|12382,12385
(|12386,12387
1|12387,12388
)|12388,12389
Tablet|12390,12396
PO|12397,12399
DAILY|12400,12405
<EOL>|12406,12407
(|12407,12408
Daily|12408,12413
)|12413,12414
.|12414,12415
<EOL>|12417,12418
8.|12418,12420
ranitidine|12421,12431
HCl|12432,12435
150|12436,12439
mg|12440,12442
Tablet|12443,12449
Sig|12450,12453
:|12453,12454
One|12455,12458
(|12459,12460
1|12460,12461
)|12461,12462
Tablet|12463,12469
PO|12470,12472
DAILY|12473,12478
<EOL>|12479,12480
(|12480,12481
Daily|12481,12486
)|12486,12487
.|12487,12488
<EOL>|12490,12491
9.|12491,12493
calcitriol|12494,12504
0.25|12505,12509
mcg|12510,12513
Capsule|12514,12521
Sig|12522,12525
:|12525,12526
One|12527,12530
(|12531,12532
1|12532,12533
)|12533,12534
Capsule|12535,12542
PO|12543,12545
DAILY|12546,12551
<EOL>|12552,12553
(|12553,12554
Daily|12554,12559
)|12559,12560
.|12560,12561
<EOL>|12563,12564
10.|12564,12567
folic|12568,12573
acid|12574,12578
1|12579,12580
mg|12581,12583
Tablet|12584,12590
Sig|12591,12594
:|12594,12595
One|12596,12599
(|12600,12601
1|12601,12602
)|12602,12603
Tablet|12604,12610
PO|12611,12613
DAILY|12614,12619
(|12620,12621
Daily|12621,12626
)|12626,12627
.|12627,12628
<EOL>|12629,12630
<EOL>|12631,12632
11.|12632,12635
aspirin|12636,12643
81|12644,12646
mg|12647,12649
Tablet|12650,12656
,|12656,12657
Chewable|12658,12666
Sig|12667,12670
:|12670,12671
One|12672,12675
(|12676,12677
1|12677,12678
)|12678,12679
Tablet|12680,12686
,|12686,12687
Chewable|12688,12696
<EOL>|12697,12698
PO|12698,12700
DAILY|12701,12706
(|12707,12708
Daily|12708,12713
)|12713,12714
.|12714,12715
<EOL>|12717,12718
<EOL>|12718,12719
<EOL>|12720,12721
Discharge|12721,12730
Disposition|12731,12742
:|12742,12743
<EOL>|12743,12744
Home|12744,12748
With|12749,12753
Service|12754,12761
<EOL>|12761,12762
<EOL>|12763,12764
Facility|12764,12772
:|12772,12773
<EOL>|12773,12774
_|12774,12775
_|12775,12776
_|12776,12777
<EOL>|12777,12778
<EOL>|12779,12780
Discharge|12780,12789
Diagnosis|12790,12799
:|12799,12800
<EOL>|12800,12801
#|12801,12802
post-obstructive|12803,12819
pneumonia|12820,12829
<EOL>|12829,12830
#|12830,12831
non|12832,12835
small|12836,12841
cell|12842,12846
lung|12847,12851
cancer|12852,12858
stage|12859,12864
IV|12865,12867
,|12867,12868
progressing|12869,12880
<EOL>|12880,12881
.|12881,12882
<EOL>|12882,12883
SECONDARY|12883,12892
DIAGNOSES|12893,12902
:|12902,12903
<EOL>|12903,12904
#|12904,12905
anemia|12906,12912
of|12913,12915
acute|12916,12921
inflammation|12922,12934
<EOL>|12934,12935
#|12935,12936
CAD|12937,12940
s|12941,12942
/|12942,12943
p|12943,12944
MI|12945,12947
<EOL>|12947,12948
#|12948,12949
chronic|12950,12957
systolic|12958,12966
CHF|12967,12970
<EOL>|12970,12971
#|12971,12972
HTN|12973,12976
<EOL>|12976,12977
#|12977,12978
CKD|12979,12982
stage|12983,12988
III|12989,12992
<EOL>|12992,12993
<EOL>|12993,12994
<EOL>|12995,12996
Discharge|12996,13005
Condition|13006,13015
:|13015,13016
<EOL>|13016,13017
Mental|13017,13023
Status|13024,13030
:|13030,13031
Clear|13032,13037
and|13038,13041
coherent|13042,13050
.|13050,13051
<EOL>|13051,13052
Level|13052,13057
of|13058,13060
Consciousness|13061,13074
:|13074,13075
Alert|13076,13081
and|13082,13085
interactive|13086,13097
.|13097,13098
<EOL>|13098,13099
Activity|13099,13107
Status|13108,13114
:|13114,13115
Ambulatory|13116,13126
-|13127,13128
requires|13129,13137
assistance|13138,13148
or|13149,13151
aid|13152,13155
(|13156,13157
walker|13157,13163
<EOL>|13164,13165
or|13165,13167
cane|13168,13172
)|13172,13173
.|13173,13174
<EOL>|13174,13175
<EOL>|13175,13176
<EOL>|13177,13178
Discharge|13178,13187
Instructions|13188,13200
:|13200,13201
<EOL>|13201,13202
You|13202,13205
were|13206,13210
admitted|13211,13219
with|13220,13224
cough|13225,13230
and|13231,13234
found|13235,13240
to|13241,13243
have|13244,13248
low|13249,13252
oxygen|13253,13259
levels|13260,13266
<EOL>|13267,13268
which|13268,13273
required|13274,13282
the|13283,13286
Intensive|13287,13296
Care|13297,13301
Unit|13302,13306
.|13306,13307
Your|13308,13312
CT|13313,13315
shows|13316,13321
<EOL>|13322,13323
progression|13323,13334
of|13335,13337
your|13338,13342
lung|13343,13347
cancer|13348,13354
with|13355,13359
a|13360,13361
probable|13362,13370
superimposed|13371,13383
<EOL>|13384,13385
pneumonia|13385,13394
.|13394,13395
You|13396,13399
were|13400,13404
treated|13405,13412
with|13413,13417
antibiotics|13418,13429
and|13430,13433
oxygen|13434,13440
and|13441,13444
<EOL>|13445,13446
improved|13446,13454
,|13454,13455
and|13456,13459
you|13460,13463
were|13464,13468
tranferred|13469,13479
to|13480,13482
the|13483,13486
medical|13487,13494
floor|13495,13500
.|13500,13501
You|13502,13505
were|13506,13510
<EOL>|13511,13512
continued|13512,13521
on|13522,13524
antibiotics|13525,13536
,|13536,13537
and|13538,13541
your|13542,13546
oxygen|13547,13553
levels|13554,13560
were|13561,13565
monitored|13566,13575
<EOL>|13576,13577
closely|13577,13584
.|13584,13585
We|13586,13588
communicated|13589,13601
with|13602,13606
your|13607,13611
primary|13612,13619
oncologist|13620,13630
,|13630,13631
Dr|13632,13634
.|13634,13635
<EOL>|13636,13637
_|13637,13638
_|13638,13639
_|13639,13640
,|13640,13641
who|13642,13645
will|13646,13650
weigh|13651,13656
the|13657,13660
risks|13661,13666
and|13667,13670
benefits|13671,13679
of|13680,13682
<EOL>|13683,13684
additional|13684,13694
chemotherapy|13695,13707
,|13707,13708
as|13709,13711
it|13712,13714
will|13715,13719
be|13720,13722
complicated|13723,13734
by|13735,13737
your|13738,13742
<EOL>|13743,13744
kidney|13744,13750
dysfunction|13751,13762
and|13763,13766
other|13767,13772
medical|13773,13780
problems|13781,13789
.|13789,13790
He|13791,13793
plans|13794,13799
to|13800,13802
<EOL>|13803,13804
repeat|13804,13810
your|13811,13815
CT|13816,13818
scan|13819,13823
once|13824,13828
you|13829,13832
finish|13833,13839
your|13840,13844
antibiotics|13845,13856
to|13857,13859
further|13860,13867
<EOL>|13868,13869
evaluate|13869,13877
the|13878,13881
rate|13882,13886
of|13887,13889
your|13890,13894
disease|13895,13902
progression|13903,13914
.|13914,13915
<EOL>|13915,13916
<EOL>|13916,13917
Your|13917,13921
congestive|13922,13932
heart|13933,13938
failure|13939,13946
has|13947,13950
been|13951,13955
stable|13956,13962
.|13962,13963
Please|13964,13970
note|13971,13975
we|13976,13978
<EOL>|13979,13980
stopped|13980,13987
your|13988,13992
lasix|13993,13998
and|13999,14002
amlodipine|14003,14013
for|14014,14017
now|14018,14021
,|14021,14022
and|14023,14026
you|14027,14030
will|14031,14035
need|14036,14040
to|14041,14043
<EOL>|14044,14045
be|14045,14047
re-evaluated|14048,14060
by|14061,14063
your|14064,14068
PCP|14069,14072
to|14073,14075
see|14076,14079
when|14080,14084
you|14085,14088
should|14089,14095
restart|14096,14103
them|14104,14108
.|14108,14109
<EOL>|14110,14111
We|14111,14113
also|14114,14118
decreased|14119,14128
your|14129,14133
evening|14134,14141
dose|14142,14146
of|14147,14149
metoprolol|14150,14160
.|14160,14161
As|14162,14164
usual|14165,14170
,|14170,14171
<EOL>|14172,14173
please|14173,14179
weigh|14180,14185
yourself|14186,14194
every|14195,14200
morning|14201,14208
,|14208,14209
and|14210,14213
call|14214,14218
MD|14219,14221
if|14222,14224
weight|14225,14231
goes|14232,14236
<EOL>|14237,14238
up|14238,14240
more|14241,14245
than|14246,14250
3|14251,14252
lbs|14253,14256
.|14256,14257
<EOL>|14257,14258
<EOL>|14259,14260
Followup|14260,14268
Instructions|14269,14281
:|14281,14282
<EOL>|14282,14283
_|14283,14284
_|14284,14285
_|14285,14286
<EOL>|14286,14287

