 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|43,52|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|43,52|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|43,57|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|77,86|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|77,86|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|77,91|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|133,136|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|144,151|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|144,151|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|153,161|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Drug|Organic Chemical|Allergies|176,183|false|false|false|C0591292|Corgard|Corgard
Drug|Pharmacologic Substance|Allergies|176,183|false|false|false|C0591292|Corgard|Corgard
Drug|Amino Acid, Peptide, or Protein|Allergies|186,193|false|false|false|C0728763|Vasotec|Vasotec
Drug|Pharmacologic Substance|Allergies|186,193|false|false|false|C0728763|Vasotec|Vasotec
Event|Event|Allergies|196,205|false|false|false|||Attending
Finding|Functional Concept|Allergies|196,205|false|false|false|C1999232|Attending (action)|Attending
Event|Event|Chief Complaint|231,238|false|false|false|||Dyspnea
Finding|Finding|Chief Complaint|231,238|false|false|false|C0013404;C2024878|Dyspnea|Dyspnea
Finding|Sign or Symptom|Chief Complaint|231,238|false|false|false|C0013404;C2024878|Dyspnea|Dyspnea
Finding|Sign or Symptom|Chief Complaint|231,250|false|false|false|C0231807|Dyspnea on exertion|Dyspnea on Exertion
Event|Event|Chief Complaint|242,250|false|false|false|||Exertion
Finding|Organism Function|Chief Complaint|242,250|false|false|false|C0015264|Exertion|Exertion
Finding|Classification|Chief Complaint|253,258|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|259,267|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|259,267|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|271,289|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|280,289|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|280,289|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|280,289|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|280,289|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|280,289|false|false|false|C0184661|Interventional procedure|Procedure
Finding|Functional Concept|History of Present Illness|391,398|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|FAILURE
Finding|Idea or Concept|History of Present Illness|391,398|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|FAILURE
Finding|Individual Behavior|History of Present Illness|391,398|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|FAILURE
Procedure|Health Care Activity|History of Present Illness|399,408|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|History of Present Illness|409,413|false|false|false|||NOTE
Event|Event|History of Present Illness|475,485|false|false|false|||OUTPATIENT
Finding|Classification|History of Present Illness|475,485|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|OUTPATIENT
Finding|Idea or Concept|History of Present Illness|475,485|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|OUTPATIENT
Anatomy|Body System|History of Present Illness|514,524|false|false|false|C0007226|Cardiovascular system|cardiology
Anatomy|Body Space or Junction|History of Present Illness|541,544|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|History of Present Illness|541,544|false|false|false|C0018802|Congestive heart failure|CHF
Disorder|Disease or Syndrome|History of Present Illness|546,549|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|546,549|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|History of Present Illness|546,549|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|546,549|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|History of Present Illness|546,549|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|History of Present Illness|546,549|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|History of Present Illness|546,549|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|History of Present Illness|546,549|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|History of Present Illness|546,549|false|false|false|||PCP
Finding|Gene or Genome|History of Present Illness|546,549|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|History of Present Illness|546,549|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Finding|History of Present Illness|562,577|false|false|false|C0277786|Chief complaint (finding)|CHIEF COMPLAINT
Attribute|Clinical Attribute|History of Present Illness|568,577|false|false|false|C3864418||COMPLAINT
Finding|Finding|History of Present Illness|568,577|false|false|false|C5441521|Complaint (finding)|COMPLAINT
Event|Event|History of Present Illness|580,587|false|false|false|||Dyspnea
Finding|Finding|History of Present Illness|580,587|false|false|false|C0013404;C2024878|Dyspnea|Dyspnea
Finding|Sign or Symptom|History of Present Illness|580,587|false|false|false|C0013404;C2024878|Dyspnea|Dyspnea
Finding|Sign or Symptom|History of Present Illness|580,599|false|false|false|C0231807|Dyspnea on exertion|Dyspnea on Exertion
Event|Event|History of Present Illness|591,599|false|false|false|||Exertion
Finding|Organism Function|History of Present Illness|591,599|false|false|false|C0015264|Exertion|Exertion
Event|Event|History of Present Illness|600,607|false|false|false|||HISTORY
Finding|Conceptual Entity|History of Present Illness|600,607|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|HISTORY
Finding|Finding|History of Present Illness|600,607|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|HISTORY
Finding|Functional Concept|History of Present Illness|600,607|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|HISTORY
Finding|Finding|History of Present Illness|600,610|false|false|false|C0262926|Medical History|HISTORY OF
Finding|Idea or Concept|History of Present Illness|611,621|true|false|false|C0449450|Presentation|PRESENTING
Event|Event|History of Present Illness|622,629|false|false|false|||ILLNESS
Finding|Sign or Symptom|History of Present Illness|622,629|false|false|false|C0221423|Illness (finding)|ILLNESS
Event|Event|History of Present Illness|672,679|false|false|false|||medical
Finding|Functional Concept|History of Present Illness|672,679|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|History of Present Illness|672,679|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|History of Present Illness|672,679|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|History of Present Illness|672,679|false|false|false|C0199168|Medical service|medical
Event|Event|History of Present Illness|680,687|false|false|false|||history
Finding|Conceptual Entity|History of Present Illness|680,687|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|680,687|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|680,687|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Event|Event|History of Present Illness|688,697|false|false|false|||pertinent
Event|Event|History of Present Illness|702,707|false|false|false|||HFrEF
Disorder|Disease or Syndrome|History of Present Illness|717,720|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|717,720|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|History of Present Illness|717,720|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|History of Present Illness|717,720|false|false|false|||CAD
Finding|Gene or Genome|History of Present Illness|717,720|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|History of Present Illness|717,720|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|History of Present Illness|717,720|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|717,720|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|725,729|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|745,748|false|false|false|C2713669|SERPINA5 protein, human|PCI
Drug|Biologically Active Substance|History of Present Illness|745,748|false|false|false|C2713669|SERPINA5 protein, human|PCI
Event|Event|History of Present Illness|745,748|false|false|false|||PCI
Finding|Gene or Genome|History of Present Illness|745,748|false|false|false|C1418370;C1705930;C4049621|Peritoneal Cancer Index;SERPINA5 gene;SERPINA5 wt Allele|PCI
Finding|Intellectual Product|History of Present Illness|745,748|false|false|false|C1418370;C1705930;C4049621|Peritoneal Cancer Index;SERPINA5 gene;SERPINA5 wt Allele|PCI
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|745,748|false|false|false|C1514496;C1532338;C4724254|Percutaneous Coronary Intervention;Prophylactic Cranial Irradiation;photochemical internalization|PCI
Finding|Finding|History of Present Illness|750,758|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|History of Present Illness|750,758|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Finding|History of Present Illness|750,782|false|false|false|C3276922|Tricuspid regurgitation, moderate|moderate tricuspid regurgitation
Disorder|Disease or Syndrome|History of Present Illness|759,782|false|false|false|C0040961|Tricuspid Valve Insufficiency|tricuspid regurgitation
Event|Event|History of Present Illness|769,782|false|false|false|||regurgitation
Finding|Finding|History of Present Illness|769,782|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|History of Present Illness|769,782|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|History of Present Illness|769,782|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Event|Event|History of Present Illness|784,789|false|false|false|||right
Finding|Functional Concept|History of Present Illness|784,789|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|790,801|false|false|false|C0018827|Heart Ventricle|ventricular
Finding|Pathologic Function|History of Present Illness|790,813|false|false|false|C0242973|Ventricular Dysfunction|ventricular dysfunction
Disorder|Disease or Syndrome|History of Present Illness|802,813|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Event|Event|History of Present Illness|802,813|false|false|false|||dysfunction
Finding|Conceptual Entity|History of Present Illness|802,813|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|History of Present Illness|802,813|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|History of Present Illness|802,813|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Finding|History of Present Illness|815,823|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|History of Present Illness|815,823|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Pathologic Function|History of Present Illness|815,846|false|false|false|C5395246|Moderate pulmonary hypertension|moderate pulmonary hypertension
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|824,833|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|History of Present Illness|824,833|false|false|false|C2707265||pulmonary
Finding|Finding|History of Present Illness|824,833|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|History of Present Illness|824,846|false|false|false|C0020542|Pulmonary Hypertension|pulmonary hypertension
Disorder|Disease or Syndrome|History of Present Illness|834,846|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|History of Present Illness|834,846|false|false|false|||hypertension
Disorder|Disease or Syndrome|History of Present Illness|852,882|false|false|false|C0235480|Paroxysmal atrial fibrillation|paroxysmal atrial fibrillation
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|863,869|false|false|false|C0018792|Heart Atrium|atrial
Attribute|Clinical Attribute|History of Present Illness|863,882|false|false|false|C2926591||atrial fibrillation
Disorder|Disease or Syndrome|History of Present Illness|863,882|false|false|false|C0004238|Atrial Fibrillation|atrial fibrillation
Lab|Laboratory or Test Result|History of Present Illness|863,882|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|atrial fibrillation
Disorder|Disease or Syndrome|History of Present Illness|870,882|false|false|false|C0232197|Fibrillation|fibrillation
Event|Event|History of Present Illness|870,882|false|false|false|||fibrillation
Drug|Organic Chemical|History of Present Illness|886,894|false|false|false|C1831808|apixaban|apixaban
Drug|Pharmacologic Substance|History of Present Illness|886,894|false|false|false|C1831808|apixaban|apixaban
Event|Event|History of Present Illness|886,894|false|false|false|||apixaban
Attribute|Clinical Attribute|History of Present Illness|896,901|false|false|false|C1300072|Tumor stage|stage
Event|Event|History of Present Illness|906,913|false|false|false|||chronic
Finding|Intellectual Product|History of Present Illness|906,913|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|History of Present Illness|906,913|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|914,920|false|false|false|C0022646;C0227665|Both kidneys;Kidney|kidney
Disorder|Neoplastic Process|History of Present Illness|914,920|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|kidney
Finding|Sign or Symptom|History of Present Illness|914,920|false|false|false|C0812426|Kidney problem|kidney
Procedure|Diagnostic Procedure|History of Present Illness|914,920|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|914,920|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Disorder|Disease or Syndrome|History of Present Illness|914,928|false|false|false|C0022658|Kidney Diseases|kidney disease
Disorder|Disease or Syndrome|History of Present Illness|921,928|false|false|false|C0012634|Disease|disease
Event|Event|History of Present Illness|921,928|false|false|false|||disease
Drug|Biomedical or Dental Material|History of Present Illness|930,938|false|false|false|C0168634|BaseLine dental cement|Baseline
Finding|Idea or Concept|History of Present Illness|930,938|false|false|false|C1552824|baseline - TableCellVerticalAlign|Baseline
Disorder|Disease or Syndrome|History of Present Illness|952,975|false|false|false|C0007820|Cerebrovascular Disorders|cerebrovascular disease
Disorder|Disease or Syndrome|History of Present Illness|968,975|false|false|false|C0012634|Disease|disease
Event|Event|History of Present Illness|968,975|false|false|false|||disease
Finding|Functional Concept|History of Present Illness|981,991|false|false|false|C0036525;C1522484|Metastatic to;metastatic qualifier|metastatic
Disorder|Neoplastic Process|History of Present Illness|981,1000|false|false|false|C0278883|Metastatic melanoma|metastatic melanoma
Disorder|Neoplastic Process|History of Present Illness|992,1000|false|false|false|C0025202|melanoma|melanoma
Drug|Immunologic Factor|History of Present Illness|992,1000|false|false|false|C0796561|Melanoma vaccine|melanoma
Drug|Pharmacologic Substance|History of Present Illness|992,1000|false|false|false|C0796561|Melanoma vaccine|melanoma
Event|Event|History of Present Illness|992,1000|false|false|false|||melanoma
Disorder|Neoplastic Process|History of Present Illness|992,1019|false|false|false|C4745280|Melanoma of Unknown Primary|melanoma of unknown primary
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1004,1011|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Immunologic Factor|History of Present Illness|1004,1011|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Pharmacologic Substance|History of Present Illness|1004,1011|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Event|Event|History of Present Illness|1004,1011|false|false|false|||unknown
Finding|Finding|History of Present Illness|1004,1011|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Functional Concept|History of Present Illness|1004,1011|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Idea or Concept|History of Present Illness|1004,1011|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Intellectual Product|History of Present Illness|1004,1011|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Event|Event|History of Present Illness|1023,1033|false|false|false|||checkpoint
Finding|Cell Function|History of Present Illness|1023,1033|false|false|false|C1155874|Cell Cycle Checkpoints|checkpoint
Drug|Biologically Active Substance|History of Present Illness|1034,1043|false|false|false|C1999216|Inhibitor|inhibitor
Event|Event|History of Present Illness|1034,1043|false|false|false|||inhibitor
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1044,1057|false|false|false|C3658706|pembrolizumab|pembrolizumab
Drug|Immunologic Factor|History of Present Illness|1044,1057|false|false|false|C3658706|pembrolizumab|pembrolizumab
Drug|Pharmacologic Substance|History of Present Illness|1044,1057|false|false|false|C3658706|pembrolizumab|pembrolizumab
Event|Event|History of Present Illness|1044,1057|false|false|false|||pembrolizumab
Event|Event|History of Present Illness|1066,1071|false|false|false|||found
Finding|Intellectual Product|History of Present Illness|1072,1078|false|false|false|C1705102|Volume (publication)|volume
Event|Event|History of Present Illness|1105,1108|false|false|false|||DOE
Finding|Sign or Symptom|History of Present Illness|1105,1108|false|false|false|C0231807|Dyspnea on exertion|DOE
Event|Event|History of Present Illness|1110,1118|false|false|false|||admitted
Event|Event|History of Present Illness|1133,1141|false|false|false|||diuresis
Finding|Organ or Tissue Function|History of Present Illness|1133,1141|false|false|false|C0012797|Diuresis|diuresis
Finding|Idea or Concept|History of Present Illness|1149,1171|false|false|false|C1546461|Most recent outpatient|most recent outpatient
Finding|Classification|History of Present Illness|1161,1171|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|History of Present Illness|1161,1171|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Anatomy|Body Space or Junction|History of Present Illness|1172,1175|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|History of Present Illness|1172,1175|false|false|false|C0018802|Congestive heart failure|CHF
Event|Event|History of Present Illness|1176,1181|false|false|false|||notes
Event|Event|History of Present Illness|1191,1195|false|false|false|||seen
Anatomy|Cell Component|History of Present Illness|1211,1214|false|false|false|C1166663|actomyosin contractile ring|car
Disorder|Disease or Syndrome|History of Present Illness|1211,1214|false|false|false|C0406810|Carney Complex|car
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1211,1214|false|false|false|C3539542;C4039583;C5890846|Chimeric antigen receptor;Coxsackievirus and Adenovirus Receptor, human;Extracellular Calcium-Sensing Receptor, Human|car
Drug|Biologically Active Substance|History of Present Illness|1211,1214|false|false|false|C3539542;C4039583;C5890846|Chimeric antigen receptor;Coxsackievirus and Adenovirus Receptor, human;Extracellular Calcium-Sensing Receptor, Human|car
Drug|Immunologic Factor|History of Present Illness|1211,1214|false|false|false|C3539542;C4039583;C5890846|Chimeric antigen receptor;Coxsackievirus and Adenovirus Receptor, human;Extracellular Calcium-Sensing Receptor, Human|car
Finding|Gene or Genome|History of Present Illness|1211,1214|false|false|false|C1413828;C1417827;C1420354;C1547285;C1706434;C1858724;C2239319;C3273602;C3540475;C3811749;C4039583;C5890846;C5890847;C5960871|CASR wt Allele;CXADR gene;CXADR wt Allele;CXADRP1 gene;Car - Mode of Arrival Code;Caronte Gene;Chimeric antigen receptor;Extracellular Calcium-Sensing Receptor, Human;NR1I3 gene;NR1I3 wt Allele;PRKAR1A wt Allele;SPG7 gene;SPG7 wt Allele;TRIM13 wt Allele|car
Finding|Intellectual Product|History of Present Illness|1211,1214|false|false|false|C1413828;C1417827;C1420354;C1547285;C1706434;C1858724;C2239319;C3273602;C3540475;C3811749;C4039583;C5890846;C5890847;C5960871|CASR wt Allele;CXADR gene;CXADR wt Allele;CXADRP1 gene;Car - Mode of Arrival Code;Caronte Gene;Chimeric antigen receptor;Extracellular Calcium-Sensing Receptor, Human;NR1I3 gene;NR1I3 wt Allele;PRKAR1A wt Allele;SPG7 gene;SPG7 wt Allele;TRIM13 wt Allele|car
Finding|Receptor|History of Present Illness|1211,1214|false|false|false|C1413828;C1417827;C1420354;C1547285;C1706434;C1858724;C2239319;C3273602;C3540475;C3811749;C4039583;C5890846;C5890847;C5960871|CASR wt Allele;CXADR gene;CXADR wt Allele;CXADRP1 gene;Car - Mode of Arrival Code;Caronte Gene;Chimeric antigen receptor;Extracellular Calcium-Sensing Receptor, Human;NR1I3 gene;NR1I3 wt Allele;PRKAR1A wt Allele;SPG7 gene;SPG7 wt Allele;TRIM13 wt Allele|car
Event|Event|History of Present Illness|1223,1235|false|false|false|||Cardiologist
Finding|Finding|History of Present Illness|1245,1262|false|false|false|C2673338|Increased fatigue|increased fatigue
Event|Event|History of Present Illness|1255,1262|false|false|false|||fatigue
Finding|Sign or Symptom|History of Present Illness|1255,1262|false|false|false|C0015672|Fatigue|fatigue
Finding|Sign or Symptom|History of Present Illness|1267,1277|false|false|false|C0239313|exercise induced|exertional
Finding|Sign or Symptom|History of Present Illness|1267,1285|false|false|false|C0231807|Dyspnea on exertion|exertional dyspnea
Event|Event|History of Present Illness|1278,1285|false|false|false|||dyspnea
Finding|Finding|History of Present Illness|1278,1285|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|History of Present Illness|1278,1285|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Event|Event|History of Present Illness|1306,1310|false|false|false|||felt
Attribute|Clinical Attribute|History of Present Illness|1315,1319|false|false|false|C0428772|Left ventricular ejection fraction|LVEF
Event|Event|History of Present Illness|1315,1319|false|false|false|||LVEF
Procedure|Diagnostic Procedure|History of Present Illness|1315,1319|false|false|false|C3837267|LVEF (procedure)|LVEF
Event|Event|History of Present Illness|1333,1340|false|false|false|||reduced
Event|Event|History of Present Illness|1360,1367|false|false|false|||started
Finding|Finding|History of Present Illness|1371,1374|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|History of Present Illness|1371,1374|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Procedure|Research Activity|History of Present Illness|1371,1379|false|false|false|C1708745|Low-Dose Treatment|low-dose
Drug|Organic Chemical|History of Present Illness|1380,1388|false|false|false|C4033616|Entresto|Entresto
Drug|Pharmacologic Substance|History of Present Illness|1380,1388|false|false|false|C4033616|Entresto|Entresto
Event|Event|History of Present Illness|1380,1388|false|false|false|||Entresto
Event|Event|History of Present Illness|1403,1411|true|false|false|||tolerate
Event|Event|History of Present Illness|1425,1436|true|false|false|||prospective
Drug|Organic Chemical|History of Present Illness|1459,1467|false|false|false|C0126174|losartan|losartan
Drug|Pharmacologic Substance|History of Present Illness|1459,1467|false|false|false|C0126174|losartan|losartan
Event|Event|History of Present Illness|1459,1467|false|false|false|||losartan
Event|Event|History of Present Illness|1478,1485|false|false|false|||stopped
Event|Event|History of Present Illness|1498,1513|false|false|false|||lightheadedness
Finding|Sign or Symptom|History of Present Illness|1498,1513|false|false|false|C0220870|Lightheadedness|lightheadedness
Event|Event|History of Present Illness|1515,1524|false|false|false|||dizziness
Finding|Sign or Symptom|History of Present Illness|1515,1524|false|false|false|C0012833;C0042571|Dizziness;Vertigo|dizziness
Event|Event|History of Present Illness|1529,1538|false|false|false|||worsening
Finding|Idea or Concept|History of Present Illness|1529,1538|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1539,1544|false|false|false|C0022646|Kidney|renal
Disorder|Disease or Syndrome|History of Present Illness|1539,1544|false|false|false|C0042075|Urologic Diseases|renal
Event|Event|History of Present Illness|1545,1553|false|false|false|||function
Finding|Finding|History of Present Illness|1545,1553|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|History of Present Illness|1545,1553|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|History of Present Illness|1545,1553|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|History of Present Illness|1545,1553|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Event|Event|History of Present Illness|1563,1570|false|false|false|||concern
Finding|Idea or Concept|History of Present Illness|1563,1570|false|false|false|C2699424|Concern|concern
Disorder|Disease or Syndrome|History of Present Illness|1596,1607|false|false|false|C0027059|Myocarditis|myocarditis
Event|Event|History of Present Illness|1596,1607|false|false|false|||myocarditis
Disorder|Neoplastic Process|History of Present Illness|1608,1617|false|false|false|C0027627|Neoplasm Metastasis|secondary
Event|Event|History of Present Illness|1608,1617|false|false|false|||secondary
Finding|Functional Concept|History of Present Illness|1608,1617|false|false|false|C1522484|metastatic qualifier|secondary
Finding|Cell Function|History of Present Illness|1625,1635|false|false|false|C1155874|Cell Cycle Checkpoints|checkpoint
Drug|Biologically Active Substance|History of Present Illness|1636,1645|false|false|false|C1999216|Inhibitor|inhibitor
Event|Event|History of Present Illness|1636,1645|false|false|false|||inhibitor
Disorder|Neoplastic Process|History of Present Illness|1676,1684|false|false|false|C0027651|Neoplasms|Oncology
Procedure|Health Care Activity|History of Present Illness|1676,1684|false|false|false|C1555459|oncology services|Oncology
Event|Event|History of Present Illness|1702,1710|false|false|false|||symptoms
Finding|Functional Concept|History of Present Illness|1702,1710|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|History of Present Illness|1702,1710|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Finding|History of Present Illness|1716,1724|false|false|false|C2984079|Somewhat|somewhat
Event|Event|History of Present Illness|1725,1733|false|false|false|||improved
Finding|Finding|History of Present Illness|1725,1733|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Finding|Intellectual Product|History of Present Illness|1725,1733|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1735,1742|false|false|false|C0018787|Heart|Cardiac
Finding|Intellectual Product|History of Present Illness|1735,1742|false|false|false|C1314974|Cardiac attachment|Cardiac
Attribute|Clinical Attribute|History of Present Illness|1735,1753|false|false|false|C2735101;C2735102|Cardiac biomarkers|Cardiac biomarkers
Attribute|Clinical Attribute|History of Present Illness|1743,1753|false|false|false|C0005516|Biological Markers|biomarkers
Event|Event|History of Present Illness|1743,1753|false|false|false|||biomarkers
Event|Event|History of Present Illness|1759,1766|false|false|false|||notable
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1780,1788|false|false|false|C0669479|pro-brain natriuretic peptide (1-76)|NTproBNP
Drug|Biologically Active Substance|History of Present Illness|1780,1788|false|false|false|C0669479|pro-brain natriuretic peptide (1-76)|NTproBNP
Event|Event|History of Present Illness|1780,1788|false|false|false|||NTproBNP
Event|Event|History of Present Illness|1793,1796|false|false|false|||10K
Event|Event|History of Present Illness|1801,1807|false|false|false|||normal
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1808,1813|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|History of Present Illness|1808,1813|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|History of Present Illness|1808,1813|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|History of Present Illness|1808,1813|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Event|Event|History of Present Illness|1828,1836|false|false|false|||elevated
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1838,1846|false|false|false|C0041199|Troponin|troponin
Drug|Biologically Active Substance|History of Present Illness|1838,1846|false|false|false|C0041199|Troponin|troponin
Event|Event|History of Present Illness|1838,1846|false|false|false|||troponin
Procedure|Laboratory Procedure|History of Present Illness|1838,1846|false|false|false|C0523952|Troponin measurement|troponin
Event|Event|History of Present Illness|1871,1881|true|false|false|||unexpected
Finding|Intellectual Product|History of Present Illness|1871,1881|true|true|false|C4055646|Unexpected|unexpected
Finding|Mental Process|History of Present Illness|1889,1896|true|false|false|C0542559|contextual factors|setting
Event|Event|History of Present Illness|1918,1925|false|false|false|||failure
Finding|Functional Concept|History of Present Illness|1918,1925|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|History of Present Illness|1918,1925|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|History of Present Illness|1918,1925|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|History of Present Illness|1930,1937|false|false|false|||chronic
Finding|Intellectual Product|History of Present Illness|1930,1937|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|History of Present Illness|1930,1937|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|History of Present Illness|1930,1952|false|false|false|C1561643|Chronic Kidney Diseases|chronic kidney disease
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1938,1944|false|false|false|C0022646;C0227665|Both kidneys;Kidney|kidney
Disorder|Neoplastic Process|History of Present Illness|1938,1944|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|kidney
Finding|Sign or Symptom|History of Present Illness|1938,1944|false|false|false|C0812426|Kidney problem|kidney
Procedure|Diagnostic Procedure|History of Present Illness|1938,1944|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1938,1944|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Disorder|Disease or Syndrome|History of Present Illness|1938,1952|false|false|false|C0022658|Kidney Diseases|kidney disease
Disorder|Disease or Syndrome|History of Present Illness|1945,1952|false|false|false|C0012634|Disease|disease
Event|Event|History of Present Illness|1945,1952|false|false|false|||disease
Event|Event|History of Present Illness|1962,1969|false|false|false|||planned
Drug|Pharmacologic Substance|History of Present Illness|1981,1994|false|false|false|C5848866|Immunotherapy [APC]|immunotherapy
Event|Event|History of Present Illness|1981,1994|false|false|false|||immunotherapy
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1981,1994|false|false|false|C0021083|Immunotherapy|immunotherapy
Event|Event|History of Present Illness|2007,2016|false|false|false|||treatment
Finding|Conceptual Entity|History of Present Illness|2007,2016|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|History of Present Illness|2007,2016|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|History of Present Illness|2007,2016|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|2007,2016|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Event|Event|History of Present Illness|2021,2025|false|false|false|||held
Event|Event|History of Present Illness|2042,2044|false|false|false|||Cr
Event|Event|History of Present Illness|2046,2053|false|false|false|||Recheck
Event|Event|History of Present Illness|2054,2060|false|false|false|||showed
Event|Event|History of Present Illness|2061,2072|false|false|false|||improvement
Finding|Conceptual Entity|History of Present Illness|2061,2072|false|false|false|C2986411|Improvement|improvement
Finding|Body Substance|History of Present Illness|2078,2085|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|2078,2085|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|2078,2085|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|2086,2095|false|false|false|||restarted
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|2096,2109|false|false|false|C3658706|pembrolizumab|pembrolizumab
Drug|Immunologic Factor|History of Present Illness|2096,2109|false|false|false|C3658706|pembrolizumab|pembrolizumab
Drug|Pharmacologic Substance|History of Present Illness|2096,2109|false|false|false|C3658706|pembrolizumab|pembrolizumab
Event|Event|History of Present Illness|2096,2109|false|false|false|||pembrolizumab
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|2118,2131|false|false|false|C3658706|pembrolizumab|Pembrolizumab
Drug|Immunologic Factor|History of Present Illness|2118,2131|false|false|false|C3658706|pembrolizumab|Pembrolizumab
Drug|Pharmacologic Substance|History of Present Illness|2118,2131|false|false|false|C3658706|pembrolizumab|Pembrolizumab
Event|Event|History of Present Illness|2118,2131|false|false|false|||Pembrolizumab
Event|Event|History of Present Illness|2143,2147|false|false|false|||held
Event|Event|History of Present Illness|2159,2167|false|false|false|||diarrhea
Finding|Finding|History of Present Illness|2159,2167|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|History of Present Illness|2159,2167|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Event|Event|History of Present Illness|2181,2185|false|false|false|||LFTs
Finding|Functional Concept|History of Present Illness|2191,2199|false|false|false|C0332287;C1883712|Add - instruction imperative;In addition to|addition
Event|Event|History of Present Illness|2209,2217|false|false|false|||received
Finding|Functional Concept|History of Present Illness|2218,2229|false|false|false|C1522726|Intravenous Route of Administration|intravenous
Event|Event|History of Present Illness|2230,2239|false|false|false|||hydration
Finding|Finding|History of Present Illness|2230,2239|false|false|false|C1321013;C4520800|Hydration;Hydration status|hydration
Finding|Physiologic Function|History of Present Illness|2230,2239|false|false|false|C1321013;C4520800|Hydration;Hydration status|hydration
Event|Event|History of Present Illness|2262,2267|false|false|false|||noted
Event|Event|History of Present Illness|2279,2285|false|false|false|||volume
Finding|Intellectual Product|History of Present Illness|2279,2285|false|false|false|C1705102|Volume (publication)|volume
Finding|Finding|History of Present Illness|2308,2312|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|History of Present Illness|2308,2312|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|History of Present Illness|2308,2312|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Drug|Organic Chemical|History of Present Illness|2313,2322|false|false|false|C0076840|torsemide|Torsemide
Drug|Pharmacologic Substance|History of Present Illness|2313,2322|false|false|false|C0076840|torsemide|Torsemide
Event|Event|History of Present Illness|2313,2322|false|false|false|||Torsemide
Finding|Intellectual Product|History of Present Illness|2355,2359|false|false|false|C1720594|Then - dosing instruction fragment|then
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|2373,2381|false|false|false|C0041199|Troponin|Troponin
Drug|Biologically Active Substance|History of Present Illness|2373,2381|false|false|false|C0041199|Troponin|Troponin
Procedure|Laboratory Procedure|History of Present Illness|2373,2381|false|false|false|C0523952|Troponin measurement|Troponin
Event|Event|History of Present Illness|2382,2389|false|false|false|||testing
Finding|Functional Concept|History of Present Illness|2382,2389|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|testing
Finding|Intellectual Product|History of Present Illness|2382,2389|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|testing
Event|Event|History of Present Illness|2390,2396|false|false|false|||showed
Event|Event|History of Present Illness|2413,2423|false|false|false|||attributed
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2427,2432|false|false|false|C0022646|Kidney|renal
Disorder|Disease or Syndrome|History of Present Illness|2427,2432|false|false|false|C0042075|Urologic Diseases|renal
Event|Event|History of Present Illness|2433,2446|false|false|false|||insufficiency
Finding|Functional Concept|History of Present Illness|2433,2446|false|false|false|C0231179|Insufficiency|insufficiency
Finding|Body Substance|History of Present Illness|2452,2459|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|2452,2459|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|2452,2459|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|2469,2474|false|false|false|||noted
Event|Event|History of Present Illness|2483,2487|false|false|false|||mild
Finding|Intellectual Product|History of Present Illness|2483,2487|false|false|false|C1547225|Mild Severity of Illness Code|mild
Event|Event|History of Present Illness|2488,2500|false|false|false|||hyperkalemia
Finding|Finding|History of Present Illness|2488,2500|false|false|false|C0020461;C5700154|Hyperkalemia;Serum potassium level above reference range|hyperkalemia
Drug|Biologically Active Substance|History of Present Illness|2519,2528|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Element, Ion, or Isotope|History of Present Illness|2519,2528|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Food|History of Present Illness|2519,2528|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Inorganic Chemical|History of Present Illness|2519,2528|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Pharmacologic Substance|History of Present Illness|2519,2528|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Event|Event|History of Present Illness|2519,2528|false|false|false|||potassium
Finding|Physiologic Function|History of Present Illness|2519,2528|false|false|false|C4553027|Potassium metabolic function|potassium
Procedure|Laboratory Procedure|History of Present Illness|2519,2528|false|false|false|C0202194|Potassium measurement|potassium
Drug|Pharmacologic Substance|History of Present Illness|2519,2544|false|false|false|C0561938|Potassium supplementation (product)|potassium supplementation
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|2519,2544|false|false|false|C3541460|Potassium supplement therapy|potassium supplementation
Event|Event|History of Present Illness|2529,2544|false|false|false|||supplementation
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|2529,2544|false|false|false|C0242297|Dietary Supplementation|supplementation
Event|Event|History of Present Illness|2549,2556|false|false|false|||stopped
Drug|Organic Chemical|History of Present Illness|2561,2570|false|false|false|C0076840|torsemide|torsemide
Drug|Pharmacologic Substance|History of Present Illness|2561,2570|false|false|false|C0076840|torsemide|torsemide
Event|Event|History of Present Illness|2571,2575|false|false|false|||dose
Event|Event|History of Present Illness|2576,2585|false|false|false|||increased
Event|Event|History of Present Illness|2599,2603|false|false|false|||seen
Event|Event|History of Present Illness|2611,2620|false|false|false|||Emergency
Finding|Finding|History of Present Illness|2611,2620|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Idea or Concept|History of Present Illness|2611,2620|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Intellectual Product|History of Present Illness|2611,2620|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Pathologic Function|History of Present Illness|2611,2620|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Phenomenon|Phenomenon or Process|History of Present Illness|2611,2620|false|false|false|C0013956|Emergency Situation|Emergency
Procedure|Health Care Activity|History of Present Illness|2611,2620|false|false|false|C1553500|emergency encounter|Emergency
Finding|Idea or Concept|History of Present Illness|2611,2625|false|false|false|C1546435|Encounter Referral Source - emergency room|Emergency room
Event|Event|History of Present Illness|2650,2654|false|false|false|||fall
Finding|Finding|History of Present Illness|2650,2654|false|false|false|C0085639|Falls|fall
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2670,2675|false|false|false|C0036270|Scalp structure|scalp
Disorder|Injury or Poisoning|History of Present Illness|2670,2686|false|false|false|C0240937|Scalp laceration|scalp laceration
Disorder|Injury or Poisoning|History of Present Illness|2676,2686|false|false|false|C0043246|Laceration|laceration
Event|Event|History of Present Illness|2676,2686|false|false|false|||laceration
Attribute|Clinical Attribute|History of Present Illness|2688,2695|false|false|false|C0881943||CT head
Procedure|Diagnostic Procedure|History of Present Illness|2688,2695|false|false|false|C0202691|CAT scan of head|CT head
Anatomy|Body Location or Region|History of Present Illness|2691,2695|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2691,2695|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|History of Present Illness|2691,2695|false|false|false|C0362076|Problems with head|head
Event|Event|History of Present Illness|2691,2695|false|false|false|||head
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|2691,2695|false|false|false|C0876917|Procedure on head|head
Anatomy|Body Location or Region|History of Present Illness|2691,2704|false|false|false|C0460004|Head and neck structure|head and neck
Anatomy|Body Location or Region|History of Present Illness|2700,2704|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|History of Present Illness|2700,2704|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|History of Present Illness|2700,2704|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Event|Event|History of Present Illness|2709,2721|false|false|false|||unremarkable
Event|Event|History of Present Illness|2728,2737|false|false|false|||presented
Event|Event|History of Present Illness|2773,2778|false|false|false|||visit
Finding|Social Behavior|History of Present Illness|2773,2778|false|false|false|C0545082|Visit|visit
Event|Event|History of Present Illness|2786,2792|false|false|false|||clinic
Event|Event|History of Present Illness|2802,2807|false|false|false|||noted
Attribute|Clinical Attribute|History of Present Illness|2817,2823|false|false|false|C0944911||weight
Event|Event|History of Present Illness|2817,2823|false|false|false|||weight
Finding|Finding|History of Present Illness|2817,2823|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|History of Present Illness|2817,2823|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|History of Present Illness|2817,2823|false|false|false|C1305866|Weighing patient|weight
Procedure|Laboratory Procedure|History of Present Illness|2837,2840|false|false|false|C3161851|liquid-based cytology (procedure)|lbs
Finding|Idea or Concept|History of Present Illness|2862,2866|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|History of Present Illness|2862,2866|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|History of Present Illness|2862,2866|false|false|false|C1553498|home health encounter|home
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2867,2872|false|false|false|C0222045|Integumentary scale|scale
Event|Activity|History of Present Illness|2867,2872|false|false|false|C1947916|Scaling|scale
Event|Event|History of Present Illness|2867,2872|false|false|false|||scale
Finding|Conceptual Entity|History of Present Illness|2867,2872|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Finding|Intellectual Product|History of Present Illness|2867,2872|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Event|Event|History of Present Illness|2882,2890|false|false|false|||reported
Event|Event|History of Present Illness|2891,2900|false|false|false|||decreased
Finding|Sign or Symptom|History of Present Illness|2891,2909|false|false|false|C0232462|Decrease in appetite|decreased appetite
Event|Event|History of Present Illness|2901,2909|false|false|false|||appetite
Finding|Organism Function|History of Present Illness|2901,2909|false|false|false|C0003618|Desire for food|appetite
Event|Event|History of Present Illness|2918,2928|false|false|false|||attributes
Event|Event|History of Present Illness|2932,2938|false|false|false|||eating
Drug|Food|History of Present Illness|2951,2955|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|History of Present Illness|2951,2955|false|false|false|||diet
Finding|Functional Concept|History of Present Illness|2951,2955|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|History of Present Illness|2951,2955|false|false|false|C0012159|Diet therapy|diet
Event|Activity|History of Present Illness|2981,2985|false|false|false|C1947933|care activity|care
Event|Event|History of Present Illness|2981,2985|false|false|false|||care
Finding|Finding|History of Present Illness|2981,2985|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|History of Present Illness|2981,2985|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Event|Event|History of Present Illness|2997,3002|false|false|false|||makes
Drug|Food|History of Present Illness|3007,3011|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Drug|Immunologic Factor|History of Present Illness|3007,3011|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Drug|Pharmacologic Substance|History of Present Illness|3007,3011|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Event|Event|History of Present Illness|3007,3011|false|false|false|||food
Event|Event|History of Present Illness|3021,3029|false|false|false|||adhering
Finding|Finding|History of Present Illness|3035,3038|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|History of Present Illness|3035,3038|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Finding|History of Present Illness|3035,3045|false|false|false|C0860871|Sodium decreased|low sodium
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|3035,3045|false|false|false|C0012169|Low sodium diet|low sodium
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|3035,3050|false|false|false|C0012169|Low sodium diet|low sodium diet
Drug|Biologically Active Substance|History of Present Illness|3039,3045|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|History of Present Illness|3039,3045|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|History of Present Illness|3039,3045|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Event|Event|History of Present Illness|3039,3045|false|false|false|||sodium
Finding|Physiologic Function|History of Present Illness|3039,3045|false|false|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|History of Present Illness|3039,3045|false|false|false|C0337443|Sodium measurement|sodium
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|3039,3050|false|false|false|C0301592|Sodium diet|sodium diet
Drug|Food|History of Present Illness|3046,3050|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|History of Present Illness|3046,3050|false|false|false|||diet
Finding|Functional Concept|History of Present Illness|3046,3050|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|History of Present Illness|3046,3050|false|false|false|C0012159|Diet therapy|diet
Event|Event|History of Present Illness|3069,3073|true|false|false|||like
Finding|Finding|History of Present Illness|3077,3081|true|false|false|C4281574|Much|much
Finding|Daily or Recreational Activity|History of Present Illness|3089,3101|true|false|false|C0184625||regular diet
Drug|Food|History of Present Illness|3097,3101|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|History of Present Illness|3097,3101|false|false|false|||diet
Finding|Functional Concept|History of Present Illness|3097,3101|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|History of Present Illness|3097,3101|false|false|false|C0012159|Diet therapy|diet
Event|Event|History of Present Illness|3106,3112|false|false|false|||drinks
Event|Event|History of Present Illness|3117,3124|false|false|false|||glasses
Drug|Inorganic Chemical|History of Present Illness|3128,3133|false|false|false|C0043047;C1550678|Water Specimen;water|water
Drug|Pharmacologic Substance|History of Present Illness|3128,3133|false|false|false|C0043047;C1550678|Water Specimen;water|water
Event|Event|History of Present Illness|3128,3133|false|false|false|||water
Finding|Intellectual Product|History of Present Illness|3128,3133|false|false|false|C1547961|Water - Specimen Source Codes|water
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|3128,3133|false|false|false|C0020311|Hydrotherapy|water
Drug|Food|History of Present Illness|3137,3142|false|false|false|C1268568|Juice|juice
Event|Event|History of Present Illness|3137,3142|false|false|false|||juice
Event|Event|History of Present Illness|3157,3163|false|false|false|||taking
Drug|Organic Chemical|History of Present Illness|3164,3173|false|false|false|C0076840|torsemide|torsemide
Drug|Pharmacologic Substance|History of Present Illness|3164,3173|false|false|false|C0076840|torsemide|torsemide
Event|Event|History of Present Illness|3164,3173|false|false|false|||torsemide
Event|Event|History of Present Illness|3195,3204|false|false|false|||decreased
Finding|Finding|History of Present Illness|3220,3232|false|false|false|C3845714|Several days|several days
Finding|Gene or Genome|History of Present Illness|3233,3236|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|History of Present Illness|3243,3247|false|false|false|||felt
Event|Event|History of Present Illness|3255,3264|false|false|false|||urinating
Event|Event|History of Present Illness|3289,3292|false|false|false|||ran
Drug|Organic Chemical|History of Present Illness|3300,3310|false|false|false|C0257343|tamsulosin|tamsulosin
Drug|Pharmacologic Substance|History of Present Illness|3300,3310|false|false|false|C0257343|tamsulosin|tamsulosin
Event|Event|History of Present Illness|3300,3310|false|false|false|||tamsulosin
Finding|Finding|History of Present Illness|3311,3323|false|false|false|C3845714|Several days|several days
Finding|Gene or Genome|History of Present Illness|3324,3327|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|History of Present Illness|3331,3338|false|false|false|||stopped
Event|Event|History of Present Illness|3339,3345|false|false|false|||taking
Finding|Finding|History of Present Illness|3367,3371|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|History of Present Illness|3367,3371|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|History of Present Illness|3367,3371|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|History of Present Illness|3376,3381|false|false|false|||noted
Event|Event|History of Present Illness|3382,3390|false|false|false|||becoming
Finding|Body Substance|History of Present Illness|3401,3407|false|false|false|C0225386|Breath|breath
Event|Event|History of Present Illness|3414,3420|false|false|false|||taking
Event|Event|History of Present Illness|3424,3429|false|false|false|||steps
Finding|Conceptual Entity|History of Present Illness|3424,3429|false|false|false|C1261552|Step (specific stage)|steps
Procedure|Health Care Activity|History of Present Illness|3424,3429|false|false|false|C4722257|STEPS to Enhance Physical Activity|steps
Event|Event|History of Present Illness|3450,3456|false|false|false|||volume
Finding|Intellectual Product|History of Present Illness|3450,3456|false|false|false|C1705102|Volume (publication)|volume
Event|Event|History of Present Illness|3468,3473|false|false|false|||noted
Event|Event|History of Present Illness|3477,3481|false|false|false|||exam
Finding|Functional Concept|History of Present Illness|3477,3481|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|History of Present Illness|3477,3481|false|false|false|C0582103|Medical Examination|exam
Event|Event|History of Present Illness|3489,3500|false|false|false|||recommended
Event|Event|History of Present Illness|3505,3514|false|false|false|||admission
Procedure|Health Care Activity|History of Present Illness|3505,3514|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|History of Present Illness|3529,3537|false|false|false|||diuresis
Finding|Organ or Tissue Function|History of Present Illness|3529,3537|false|false|false|C0012797|Diuresis|diuresis
Anatomy|Anatomical Structure|History of Present Illness|3546,3551|false|false|false|C3714591|Floor (anatomic)|floor
Event|Event|History of Present Illness|3556,3564|false|false|false|||endorses
Finding|Idea or Concept|History of Present Illness|3569,3574|false|false|false|C1552828|Table Frame - above|above
Event|Event|History of Present Illness|3575,3582|false|false|false|||history
Finding|Conceptual Entity|History of Present Illness|3575,3582|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|3575,3582|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|3575,3582|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Event|Event|History of Present Illness|3587,3592|false|false|false|||noted
Event|Event|History of Present Illness|3602,3605|false|false|false|||SOB
Finding|Sign or Symptom|History of Present Illness|3602,3605|false|false|false|C0013404|Dyspnea|SOB
Finding|Functional Concept|History of Present Illness|3610,3621|false|false|false|C0205329|Progressive|progressive
Event|Event|History of Present Illness|3622,3628|false|false|false|||gotten
Event|Event|History of Present Illness|3629,3634|false|false|false|||worse
Finding|Finding|History of Present Illness|3629,3634|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Idea or Concept|History of Present Illness|3629,3634|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Idea or Concept|History of Present Illness|3636,3642|false|false|false|C0750554|MOSTLY|Mostly
Event|Event|History of Present Illness|3643,3649|false|false|false|||occurs
Event|Activity|History of Present Illness|3655,3663|false|false|false|C0441655|Activities|activity
Event|Event|History of Present Illness|3655,3663|false|false|false|||activity
Finding|Daily or Recreational Activity|History of Present Illness|3655,3663|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Finding|Finding|History of Present Illness|3655,3663|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Event|Event|History of Present Illness|3665,3669|false|false|false|||None
Finding|Functional Concept|History of Present Illness|3670,3677|true|false|false|C0443144|At rest (qualifier value)|at rest
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|3673,3677|true|false|false|C1742913|REST protein, human|rest
Drug|Biologically Active Substance|History of Present Illness|3673,3677|true|false|false|C1742913|REST protein, human|rest
Finding|Daily or Recreational Activity|History of Present Illness|3673,3677|true|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Gene or Genome|History of Present Illness|3673,3677|true|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Molecular Function|History of Present Illness|3673,3677|true|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Event|Event|History of Present Illness|3682,3687|false|false|false|||noted
Attribute|Clinical Attribute|History of Present Illness|3697,3703|false|false|false|C0944911||weight
Event|Event|History of Present Illness|3697,3703|false|false|false|||weight
Finding|Finding|History of Present Illness|3697,3703|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|History of Present Illness|3697,3703|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|History of Present Illness|3697,3703|false|false|false|C1305866|Weighing patient|weight
Event|Event|History of Present Illness|3721,3731|false|false|false|||decreasing
Disorder|Disease or Syndrome|History of Present Illness|3736,3752|false|false|false|C0003123|Anorexia|lack of appetite
Finding|Finding|History of Present Illness|3736,3752|false|false|false|C1971624|Loss of appetite (finding)|lack of appetite
Event|Event|History of Present Illness|3744,3752|false|false|false|||appetite
Finding|Organism Function|History of Present Illness|3744,3752|false|false|false|C0003618|Desire for food|appetite
Finding|Idea or Concept|History of Present Illness|3785,3789|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|History of Present Illness|3785,3789|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|History of Present Illness|3785,3789|false|false|false|C1553498|home health encounter|home
Procedure|Health Care Activity|History of Present Illness|3785,3796|false|false|false|C1553498|home health encounter|home health
Event|Event|History of Present Illness|3790,3796|false|false|false|||health
Finding|Idea or Concept|History of Present Illness|3790,3796|false|false|false|C0018684|Health|health
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|3797,3800|false|false|false|C1454018|AICDA protein, human|aid
Drug|Enzyme|History of Present Illness|3797,3800|false|false|false|C1454018|AICDA protein, human|aid
Event|Event|History of Present Illness|3797,3800|false|false|false|||aid
Finding|Gene or Genome|History of Present Illness|3797,3800|false|false|false|C1421876;C3540469|AICDA gene;AICDA wt Allele|aid
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|3797,3800|false|false|false|C0021588;C0280108|AID - Artificial insemination by donor;dacarbazine/doxorubicin/ifosfamide protocol|aid
Event|Event|History of Present Illness|3801,3809|false|false|false|||everyday
Event|Event|History of Present Illness|3829,3834|false|false|false|||helps
Disorder|Disease or Syndrome|History of Present Illness|3844,3847|false|false|false|C5443983|VISCERAL LEIOMYOPATHY, AFRICAN DEGENERATIVE|ADL
Event|Event|History of Present Illness|3844,3847|false|false|false|||ADL
Finding|Daily or Recreational Activity|History of Present Illness|3844,3847|false|false|false|C0001288;C1420005;C5960776|Activity of daily living (function);SGCA gene;SGCA wt Allele|ADL
Finding|Gene or Genome|History of Present Illness|3844,3847|false|false|false|C0001288;C1420005;C5960776|Activity of daily living (function);SGCA gene;SGCA wt Allele|ADL
Anatomy|Body Location or Region|History of Present Illness|3862,3871|false|false|false|C0000726|Abdomen|abdominal
Event|Event|History of Present Illness|3872,3880|false|false|false|||bloading
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|3884,3891|false|false|false|C0018787|Heart|Cardiac
Finding|Intellectual Product|History of Present Illness|3884,3891|false|false|false|C1314974|Cardiac attachment|Cardiac
Event|Event|History of Present Illness|3892,3898|false|false|false|||review
Finding|Idea or Concept|History of Present Illness|3892,3898|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Intellectual Product|History of Present Illness|3892,3898|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Functional Concept|History of Present Illness|3892,3901|false|false|false|C0699752|Review of|review of
Attribute|Clinical Attribute|History of Present Illness|3892,3909|false|false|false|C0488564;C0488565||review of systems
Procedure|Health Care Activity|History of Present Illness|3892,3909|false|false|false|C0489633|Review of systems (procedure)|review of systems
Event|Event|History of Present Illness|3902,3909|false|false|false|||systems
Finding|Functional Concept|History of Present Illness|3902,3909|false|false|false|C0449913|System|systems
Event|Event|History of Present Illness|3913,3920|false|false|false|||notable
Disorder|Anatomical Abnormality|History of Present Illness|3925,3932|false|false|false|C1689985|Absence (morphologic abnormality)|absence
Event|Event|History of Present Illness|3925,3932|false|false|false|||absence
Finding|Functional Concept|History of Present Illness|3925,3932|false|false|false|C0332197|Absent|absence
Finding|Functional Concept|History of Present Illness|3925,3935|false|false|false|C0332197|Absent|absence of
Anatomy|Body Location or Region|History of Present Illness|3936,3941|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|3936,3941|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|3936,3946|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|3936,3946|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|3942,3946|false|true|false|C2598155||pain
Event|Event|History of Present Illness|3942,3946|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|3942,3946|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|3942,3946|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Disorder|Disease or Syndrome|History of Present Illness|3948,3976|false|false|false|C1956415|Paroxysmal nocturnal dyspnea|paroxysmal nocturnal dyspnea
Event|Event|History of Present Illness|3969,3976|false|false|false|||dyspnea
Finding|Finding|History of Present Illness|3969,3976|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|History of Present Illness|3969,3976|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Event|Event|History of Present Illness|3978,3987|false|false|false|||orthopnea
Finding|Finding|History of Present Illness|3978,3987|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Finding|Sign or Symptom|History of Present Illness|3978,3987|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Event|Event|History of Present Illness|3989,4001|false|false|false|||palpitations
Finding|Finding|History of Present Illness|3989,4001|false|false|false|C0030252|Palpitations|palpitations
Event|Event|History of Present Illness|4003,4010|false|false|false|||syncope
Finding|Sign or Symptom|History of Present Illness|4003,4010|false|false|false|C0039070|Syncope|syncope
Event|Event|History of Present Illness|4015,4025|false|false|false|||presyncope
Finding|Sign or Symptom|History of Present Illness|4015,4025|false|false|false|C0700200|Presyncope|presyncope
Anatomy|Body Space or Junction|History of Present Illness|4028,4031|false|false|false|C0262327|rostral sulcus|ROS
Drug|Biologically Active Substance|History of Present Illness|4028,4031|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Element, Ion, or Isotope|History of Present Illness|4028,4031|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Organic Chemical|History of Present Illness|4028,4031|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Pharmacologic Substance|History of Present Illness|4028,4031|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Event|Event|History of Present Illness|4028,4031|false|false|false|||ROS
Finding|Gene or Genome|History of Present Illness|4028,4031|false|false|false|C0812281;C1709820|ROS1 gene;ROS1 wt Allele|ROS
Procedure|Health Care Activity|History of Present Illness|4028,4031|false|false|false|C0489633|Review of systems (procedure)|ROS
Event|Event|History of Present Illness|4042,4050|false|false|false|||negative
Finding|Classification|History of Present Illness|4042,4050|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|History of Present Illness|4042,4050|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|History of Present Illness|4042,4050|false|false|false|C5237010|Expression Negative|negative
Event|Event|History of Present Illness|4069,4074|false|false|false|||noted
Finding|Idea or Concept|History of Present Illness|4075,4080|false|false|false|C1552828|Table Frame - above|above
Finding|Finding|Past Medical History|4139,4147|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|MODERATE
Finding|Intellectual Product|Past Medical History|4139,4147|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|MODERATE
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|4148,4155|false|false|false|C0007272|Carotid Arteries|CAROTID
Disorder|Disease or Syndrome|Past Medical History|4148,4163|false|false|false|C0741975|carotid disease|CAROTID DISEASE
Disorder|Disease or Syndrome|Past Medical History|4156,4163|false|false|false|C0012634|Disease|DISEASE
Event|Event|Past Medical History|4156,4163|false|false|false|||DISEASE
Event|Event|Past Medical History|4180,4187|false|false|false|||FAILURE
Finding|Functional Concept|Past Medical History|4180,4187|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|FAILURE
Finding|Idea or Concept|Past Medical History|4180,4187|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|FAILURE
Finding|Individual Behavior|Past Medical History|4180,4187|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|FAILURE
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|4189,4197|false|false|false|C0018787|Heart|CORONARY
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|4189,4204|false|false|false|C0205042|Coronary artery|CORONARY ARTERY
Disorder|Disease or Syndrome|Past Medical History|4189,4212|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|CORONARY ARTERY DISEASE
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|4198,4204|false|false|false|C0003842;C0226004|Arterial system;Arteries|ARTERY
Anatomy|Body System|Past Medical History|4198,4204|false|false|false|C0003842;C0226004|Arterial system;Arteries|ARTERY
Disorder|Disease or Syndrome|Past Medical History|4198,4212|false|false|false|C0852949|Arteriopathic disease|ARTERY DISEASE
Disorder|Disease or Syndrome|Past Medical History|4205,4212|false|false|false|C0012634|Disease|DISEASE
Event|Event|Past Medical History|4205,4212|false|false|false|||DISEASE
Anatomy|Body Location or Region|Past Medical History|4214,4230|false|false|false|C0744316|gastroesophageal|GASTROESOPHAGEAL
Disorder|Disease or Syndrome|Past Medical History|4214,4237|false|false|false|C0017168|Gastroesophageal reflux disease|GASTROESOPHAGEAL REFLUX
Finding|Finding|Past Medical History|4214,4237|false|false|false|C3813607;C4317146|Acid reflux;Infantile Gastroesophageal Reflux|GASTROESOPHAGEAL REFLUX
Event|Event|Past Medical History|4231,4237|false|false|false|||REFLUX
Finding|Pathologic Function|Past Medical History|4231,4237|false|false|false|C0232483|Reflux|REFLUX
Disorder|Disease or Syndrome|Past Medical History|4239,4251|false|false|false|C0020538|Hypertensive disease|HYPERTENSION
Event|Event|Past Medical History|4239,4251|false|false|false|||HYPERTENSION
Finding|Finding|Past Medical History|4253,4259|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|SEVERE
Finding|Intellectual Product|Past Medical History|4253,4259|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|SEVERE
Disorder|Disease or Syndrome|Past Medical History|4260,4269|false|false|false|C0034067|Pulmonary Emphysema|EMPHYSEMA
Event|Event|Past Medical History|4260,4269|false|false|false|||EMPHYSEMA
Finding|Pathologic Function|Past Medical History|4260,4269|false|false|false|C0013990|Pathological accumulation of air in tissues|EMPHYSEMA
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|4271,4280|false|false|false|C0024109|Lung|PULMONARY
Attribute|Clinical Attribute|Past Medical History|4271,4280|false|false|false|C2707265||PULMONARY
Finding|Finding|Past Medical History|4271,4280|false|false|false|C4522268|Pulmonary (intended site)|PULMONARY
Finding|Pathologic Function|Past Medical History|4271,4293|false|false|false|C0020542|Pulmonary Hypertension|PULMONARY HYPERTENSION
Disorder|Disease or Syndrome|Past Medical History|4281,4293|false|false|false|C0020538|Hypertensive disease|HYPERTENSION
Event|Event|Past Medical History|4281,4293|false|false|false|||HYPERTENSION
Finding|Functional Concept|Past Medical History|4295,4300|false|false|false|C1552823|Table Cell Horizontal Align - right|RIGHT
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|4295,4314|false|false|false|C0225916|Structure of right branch of atrioventricular bundle|RIGHT BUNDLE BRANCH
Disorder|Disease or Syndrome|Past Medical History|4295,4320|false|false|false|C0085615|Right bundle branch block|RIGHT BUNDLE BRANCH BLOCK
Finding|Finding|Past Medical History|4295,4320|false|false|false|C0344421||RIGHT BUNDLE BRANCH BLOCK
Disorder|Disease or Syndrome|Past Medical History|4301,4320|false|false|false|C0006384;C1879286|Bundle-Branch Block;Hereditary bundle branch system defect|BUNDLE BRANCH BLOCK
Drug|Chemical Viewed Structurally|Past Medical History|4308,4314|false|false|false|C1881507|Macromolecular Branch|BRANCH
Drug|Biomedical or Dental Material|Past Medical History|4315,4320|false|false|false|C1706085|Block Dosage Form|BLOCK
Event|Event|Past Medical History|4315,4320|false|false|false|||BLOCK
Finding|Body Substance|Past Medical History|4315,4320|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|BLOCK
Finding|Finding|Past Medical History|4315,4320|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|BLOCK
Finding|Functional Concept|Past Medical History|4315,4320|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|BLOCK
Finding|Pathologic Function|Past Medical History|4322,4350|false|false|false|C1704272|Benign Prostatic Hyperplasia|BENIGN PROSTATIC HYPERTROPHY
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|4329,4338|false|false|false|C0033572|Prostate|PROSTATIC
Disorder|Disease or Syndrome|Past Medical History|4329,4350|false|false|false|C1739363|Prostatic Hypertrophy|PROSTATIC HYPERTROPHY
Finding|Pathologic Function|Past Medical History|4329,4350|false|false|false|C1704272;C2937421|Benign Prostatic Hyperplasia;Prostatic Hyperplasia|PROSTATIC HYPERTROPHY
Event|Event|Past Medical History|4339,4350|false|false|false|||HYPERTROPHY
Finding|Pathologic Function|Past Medical History|4339,4350|false|false|false|C0020564|Hypertrophy|HYPERTROPHY
Disorder|Disease or Syndrome|Past Medical History|4352,4366|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|HYPERLIPIDEMIA
Event|Event|Past Medical History|4352,4366|false|false|false|||HYPERLIPIDEMIA
Finding|Finding|Past Medical History|4352,4366|false|false|false|C0428465|Serum lipids high (finding)|HYPERLIPIDEMIA
Event|Event|Past Medical History|4368,4378|false|false|false|||PAROXYSMAL
Disorder|Disease or Syndrome|Past Medical History|4368,4398|false|false|false|C0235480|Paroxysmal atrial fibrillation|PAROXYSMAL ATRIAL FIBRILLATION
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|4379,4385|false|false|false|C0018792|Heart Atrium|ATRIAL
Attribute|Clinical Attribute|Past Medical History|4379,4398|false|false|false|C2926591||ATRIAL FIBRILLATION
Disorder|Disease or Syndrome|Past Medical History|4379,4398|false|false|false|C0004238|Atrial Fibrillation|ATRIAL FIBRILLATION
Lab|Laboratory or Test Result|Past Medical History|4379,4398|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|ATRIAL FIBRILLATION
Disorder|Disease or Syndrome|Past Medical History|4386,4398|false|false|false|C0232197|Fibrillation|FIBRILLATION
Event|Event|Past Medical History|4386,4398|false|false|false|||FIBRILLATION
Event|Event|Past Surgical History|4445,4458|false|false|false|||CARDIOVERSION
Procedure|Therapeutic or Preventive Procedure|Past Surgical History|4445,4458|false|false|false|C0013778|Electric Countershock|CARDIOVERSION
Finding|Functional Concept|Past Surgical History|4464,4469|false|false|false|C1552823|Table Cell Horizontal Align - right|RIGHT
Anatomy|Body Part, Organ, or Organ Component|Past Surgical History|4464,4480|false|false|false|C1261075|Structure of right lower lobe of lung|RIGHT LOWER LOBE
Anatomy|Body Location or Region|Past Surgical History|4470,4475|false|false|false|C1548802|Body Site Modifier - Lower|LOWER
Event|Activity|Past Surgical History|4470,4475|false|false|false|C2003888|Lower (action)|LOWER
Anatomy|Body Part, Organ, or Organ Component|Past Surgical History|4470,4480|false|false|false|C0225758|Structure of lower lobe of lung|LOWER LOBE
Anatomy|Body Part, Organ, or Organ Component|Past Surgical History|4476,4480|false|false|false|C0796494|lobe|LOBE
Finding|Gene or Genome|Past Surgical History|4476,4480|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|LOBE
Event|Event|Past Surgical History|4481,4490|false|false|false|||LOBECTOMY
Procedure|Therapeutic or Preventive Procedure|Past Surgical History|4481,4490|false|true|false|C0023928|Lobectomy|LOBECTOMY
Anatomy|Body Part, Organ, or Organ Component|Past Surgical History|4496,4504|false|false|false|C0018787|Heart|CORONARY
Procedure|Therapeutic or Preventive Procedure|Past Surgical History|4496,4511|false|false|false|C0010055|Coronary Artery Bypass Surgery|CORONARY BYPASS
Procedure|Therapeutic or Preventive Procedure|Past Surgical History|4496,4519|false|false|false|C0010055|Coronary Artery Bypass Surgery|CORONARY BYPASS SURGERY
Event|Event|Past Surgical History|4505,4511|false|false|false|||BYPASS
Procedure|Therapeutic or Preventive Procedure|Past Surgical History|4505,4511|false|false|false|C0813207|Creation of shunt|BYPASS
Procedure|Therapeutic or Preventive Procedure|Past Surgical History|4505,4519|false|false|false|C1536078|Bypass surgery|BYPASS SURGERY
Event|Event|Past Surgical History|4512,4519|false|false|false|||SURGERY
Finding|Finding|Past Surgical History|4512,4519|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Finding|Functional Concept|Past Surgical History|4512,4519|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Finding|Idea or Concept|Past Surgical History|4512,4519|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Procedure|Therapeutic or Preventive Procedure|Past Surgical History|4512,4519|false|false|false|C0543467|Operative Surgical Procedures|SURGERY
Procedure|Health Care Activity|General Exam|4598,4607|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Finding|Finding|General Exam|4608,4616|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|General Exam|4608,4616|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|General Exam|4608,4616|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|General Exam|4608,4628|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAMINATION
Procedure|Health Care Activity|General Exam|4608,4628|false|false|false|C0031809|Physical Examination|PHYSICAL EXAMINATION
Event|Activity|General Exam|4617,4628|false|false|false|C4321457|Examination|EXAMINATION
Event|Event|General Exam|4617,4628|false|false|false|||EXAMINATION
Procedure|Health Care Activity|General Exam|4617,4628|false|false|false|C0031809;C0582103|Medical Examination;Physical Examination|EXAMINATION
Event|Event|General Exam|4668,4672|false|false|false|||Data
Finding|Idea or Concept|General Exam|4668,4672|false|false|false|C1511726|Data|Data
Event|Event|General Exam|4679,4686|false|false|false|||updated
Event|Event|General Exam|4703,4707|false|false|false|||Temp
Finding|Gene or Genome|General Exam|4703,4707|false|false|false|C1823816|C1orf210 gene|Temp
Procedure|Therapeutic or Preventive Procedure|General Exam|4703,4707|false|false|false|C0279848|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Temp
Event|Event|General Exam|4769,4777|false|false|false|||delivery
Finding|Finding|General Exam|4769,4777|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Finding|Functional Concept|General Exam|4769,4777|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Finding|Organism Function|General Exam|4769,4777|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Procedure|Therapeutic or Preventive Procedure|General Exam|4769,4777|false|false|false|C0011209|Obstetric Delivery|delivery
Event|Event|General Exam|4808,4815|false|false|false|||GENERAL
Finding|Classification|General Exam|4808,4815|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|General Exam|4808,4815|false|false|false|C3812897|General medical service|GENERAL
Finding|Finding|General Exam|4817,4821|false|false|false|C5575035|Well (answer to question)|Well
Event|Event|General Exam|4822,4831|false|false|false|||developed
Finding|Finding|General Exam|4833,4837|false|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|4838,4847|false|false|false|||nourished
Event|Event|General Exam|4848,4852|false|false|false|||male
Finding|Finding|General Exam|4848,4852|false|false|false|C1706180|Male Gender|male
Disorder|Disease or Syndrome|General Exam|4856,4859|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|4856,4859|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|4856,4859|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|4856,4859|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|4856,4859|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|General Exam|4856,4859|false|false|false|||NAD
Finding|Finding|General Exam|4856,4859|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Finding|Finding|General Exam|4861,4869|false|false|false|C1961028|Oriented to place|Oriented
Attribute|Clinical Attribute|General Exam|4875,4879|false|false|false|C2713234||Mood
Event|Event|General Exam|4875,4879|false|false|false|||Mood
Finding|Conceptual Entity|General Exam|4875,4879|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Finding|Finding|General Exam|4875,4879|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Finding|Mental Process|General Exam|4875,4879|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Event|Event|General Exam|4881,4887|false|false|false|||affect
Event|Event|General Exam|4888,4899|false|false|false|||appropriate
Anatomy|Body Location or Region|General Exam|4903,4908|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|General Exam|4910,4915|false|false|false|C0036270|Scalp structure|Scalp
Disorder|Injury or Poisoning|General Exam|4910,4926|false|false|false|C0240937|Scalp laceration|Scalp laceration
Disorder|Injury or Poisoning|General Exam|4916,4926|false|false|false|C0043246|Laceration|laceration
Event|Event|General Exam|4916,4926|false|false|false|||laceration
Event|Event|General Exam|4927,4932|false|false|false|||noted
Anatomy|Body Part, Organ, or Organ Component|General Exam|4934,4940|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|General Exam|4934,4940|false|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|General Exam|4934,4940|false|false|false|||Sclera
Procedure|Health Care Activity|General Exam|4934,4940|false|false|false|C2228481|examination of sclera|Sclera
Event|Event|General Exam|4950,4957|false|false|false|||icteric
Finding|Sign or Symptom|General Exam|4950,4957|false|false|false|C0022346|Icterus|icteric
Event|Event|General Exam|4959,4964|false|false|false|||PERRL
Finding|Finding|General Exam|4959,4964|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Event|Event|General Exam|4966,4970|false|false|false|||EOMI
Anatomy|Body Part, Organ, or Organ Component|General Exam|4972,4983|false|false|false|C0009758;C0229274|Structure of palpebral conjunctiva;conjunctiva|Conjunctiva
Disorder|Disease or Syndrome|General Exam|4972,4983|false|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|Conjunctiva
Disorder|Neoplastic Process|General Exam|4972,4983|false|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|Conjunctiva
Event|Event|General Exam|4972,4983|false|false|false|||Conjunctiva
Finding|Body Substance|General Exam|4972,4983|false|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|Conjunctiva
Finding|Intellectual Product|General Exam|4972,4983|false|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|Conjunctiva
Procedure|Health Care Activity|General Exam|4972,4983|false|false|false|C0872390;C2228431|Procedure on conjunctiva;examination of conjunctiva|Conjunctiva
Event|Event|General Exam|4989,4993|false|false|false|||pink
Event|Event|General Exam|4998,5004|true|false|false|||pallor
Finding|Finding|General Exam|4998,5004|true|false|false|C0241137|Pallor of skin|pallor
Event|Event|General Exam|5008,5016|true|false|false|||cyanosis
Finding|Sign or Symptom|General Exam|5008,5016|true|false|false|C0010520|Cyanosis|cyanosis
Anatomy|Body Space or Junction|General Exam|5024,5028|true|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|General Exam|5024,5028|true|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|General Exam|5024,5028|true|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|General Exam|5024,5028|true|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Anatomy|Tissue|General Exam|5029,5035|false|false|false|C0026724|Mucous Membrane|mucosa
Finding|Intellectual Product|General Exam|5029,5035|false|false|false|C1561514||mucosa
Disorder|Disease or Syndrome|General Exam|5040,5051|true|false|false|C0155210;C0302314|Eyelid Xanthoma;Xanthoma|xanthelasma
Event|Event|General Exam|5040,5051|true|false|false|||xanthelasma
Anatomy|Body Location or Region|General Exam|5055,5059|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|General Exam|5055,5059|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|General Exam|5055,5059|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|General Exam|5061,5067|false|false|false|||Supple
Finding|Functional Concept|General Exam|5061,5067|false|false|false|C0332254|Supple|Supple
Event|Event|General Exam|5069,5072|false|false|false|||JVP
Finding|Finding|General Exam|5069,5072|false|false|false|C0428897|Jugular venous pressure|JVP
Disorder|Cell or Molecular Dysfunction|General Exam|5086,5094|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Event|Event|General Exam|5086,5094|false|false|false|||positive
Finding|Classification|General Exam|5086,5094|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|General Exam|5086,5094|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|General Exam|5095,5115|false|false|false|C5784512|Hepatojugular Reflex|hepatojugular reflex
Event|Event|General Exam|5109,5115|false|false|false|||reflex
Finding|Finding|General Exam|5109,5115|false|false|false|C0034929;C0439840;C0596002|Observation of reflex;Reflex action;Reflex motion descriptor|reflex
Finding|Organ or Tissue Function|General Exam|5109,5115|false|false|false|C0034929;C0439840;C0596002|Observation of reflex;Reflex action;Reflex motion descriptor|reflex
Anatomy|Body Part, Organ, or Organ Component|General Exam|5118,5125|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|General Exam|5118,5125|false|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Activity|General Exam|5135,5139|false|false|false|C0871208|Rating (action)|rate
Event|Event|General Exam|5135,5139|false|false|false|||rate
Finding|Idea or Concept|General Exam|5135,5139|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|General Exam|5144,5150|false|false|false|||rhythm
Finding|Finding|General Exam|5144,5150|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|General Exam|5144,5150|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Event|Event|General Exam|5185,5191|false|false|false|||murmur
Finding|Finding|General Exam|5185,5191|false|false|false|C0018808|Heart murmur|murmur
Anatomy|Cell Component|General Exam|5212,5216|true|false|false|C3890171|dinoflagellate apex|apex
Drug|Amino Acid, Peptide, or Protein|General Exam|5212,5216|true|false|false|C0140145|APEX1 protein, human|apex
Drug|Enzyme|General Exam|5212,5216|true|false|false|C0140145|APEX1 protein, human|apex
Finding|Gene or Genome|General Exam|5212,5216|true|false|false|C1332102|APEX1 gene|apex
Event|Event|General Exam|5221,5225|true|false|false|||rubs
Finding|Finding|General Exam|5221,5225|true|false|false|C0232267|Pericardial friction rub|rubs
Event|Event|General Exam|5230,5237|true|false|false|||gallops
Event|Event|General Exam|5242,5249|true|false|false|||thrills
Finding|Finding|General Exam|5242,5249|true|false|false|C0232269|Cardiac thrill (finding)|thrills
Event|Event|General Exam|5253,5258|true|false|false|||lifts
Anatomy|Body Part, Organ, or Organ Component|General Exam|5262,5267|false|false|false|C0024109|Lung|LUNGS
Anatomy|Body Location or Region|General Exam|5272,5277|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|General Exam|5272,5277|true|false|false|C0741025|Chest problem|chest
Anatomy|Body Location or Region|General Exam|5272,5282|true|false|false|C0205076;C4266615|Chest wall structure;Chest>Chest wall|chest wall
Anatomy|Body Part, Organ, or Organ Component|General Exam|5272,5282|true|false|false|C0205076;C4266615|Chest wall structure;Chest>Chest wall|chest wall
Disorder|Anatomical Abnormality|General Exam|5272,5294|true|false|false|C3164427|Deformity of chest wall|chest wall deformities
Disorder|Congenital Abnormality|General Exam|5283,5294|true|false|false|C0000768|Congenital Abnormality|deformities
Event|Event|General Exam|5283,5294|true|false|false|||deformities
Event|Event|General Exam|5298,5308|true|false|false|||tenderness
Finding|Mental Process|General Exam|5298,5308|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|General Exam|5298,5308|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Cell Function|General Exam|5310,5321|true|false|false|C0035203;C0282636|Cell Respiration;Respiration|Respiration
Finding|Physiologic Function|General Exam|5310,5321|true|false|false|C0035203;C0282636|Cell Respiration;Respiration|Respiration
Phenomenon|Biologic Function|General Exam|5310,5321|true|false|false|C1160636|respiratory system process|Respiration
Event|Event|General Exam|5325,5334|true|false|false|||unlabored
Finding|Functional Concept|General Exam|5325,5334|true|false|false|C2983702|Unlabored|unlabored
Disorder|Congenital Abnormality|General Exam|5343,5359|true|false|false|C0158784|Accessory skeletal muscle|accessory muscle
Finding|Finding|General Exam|5343,5363|true|false|false|C1821466|Use of accessory muscles|accessory muscle use
Anatomy|Body Part, Organ, or Organ Component|General Exam|5353,5359|true|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|General Exam|5353,5359|true|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Event|Event|General Exam|5360,5363|true|false|false|||use
Finding|Functional Concept|General Exam|5360,5363|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|General Exam|5360,5363|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Event|Event|General Exam|5375,5383|false|false|false|||crackles
Finding|Finding|General Exam|5375,5383|false|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Anatomy|Body Location or Region|General Exam|5385,5392|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|General Exam|5385,5392|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|General Exam|5385,5392|false|false|false|||ABDOMEN
Finding|Finding|General Exam|5385,5392|false|false|false|C0941288|Abdomen problem|ABDOMEN
Event|Event|General Exam|5401,5410|false|false|false|||distended
Finding|Finding|General Exam|5401,5410|false|false|false|C0700124|Dilated|distended
Anatomy|Body Part, Organ, or Organ Component|General Exam|5424,5429|false|false|false|C0021853|Intestines|bowel
Finding|Finding|General Exam|5424,5436|false|false|false|C0232693|Bowel sounds|bowel sounds
Event|Event|General Exam|5430,5436|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|General Exam|5430,5436|false|false|false|C0037709||sounds
Disorder|Disease or Syndrome|General Exam|5438,5442|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|General Exam|5438,5442|false|false|false|||soft
Event|Event|General Exam|5447,5457|false|false|false|||non-tender
Event|Event|General Exam|5461,5470|false|false|false|||palpation
Procedure|Diagnostic Procedure|General Exam|5461,5470|false|false|false|C0030247|Palpation|palpation
Event|Event|General Exam|5496,5508|true|false|false|||organomegaly
Finding|Finding|General Exam|5496,5508|true|false|false|C4054315|Organomegaly|organomegaly
Event|Event|General Exam|5512,5516|true|false|false|||mass
Finding|Finding|General Exam|5512,5516|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|General Exam|5512,5516|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|General Exam|5512,5516|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Anatomy|Body Part, Organ, or Organ Component|General Exam|5517,5528|true|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Phenomenon|Natural Phenomenon or Process|General Exam|5530,5534|false|false|false|C0678568||Cool
Finding|Finding|General Exam|5536,5552|false|false|false|C1720243|1+ pitting edema|1+ pitting edema
Finding|Functional Concept|General Exam|5539,5546|false|false|false|C0205323|Pitting|pitting
Finding|Finding|General Exam|5539,5552|false|false|false|C0333243|Pitting edema|pitting edema
Attribute|Clinical Attribute|General Exam|5547,5552|false|false|false|C1717255||edema
Event|Event|General Exam|5547,5552|false|false|false|||edema
Finding|Pathologic Function|General Exam|5547,5552|false|false|false|C0013604|Edema|edema
Anatomy|Body Location or Region|General Exam|5556,5560|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Part, Organ, or Organ Component|General Exam|5556,5560|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Space or Junction|General Exam|5556,5560|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Procedure|Diagnostic Procedure|General Exam|5556,5560|false|false|false|C0562271|Examination of knee joint|knee
Anatomy|Body Part, Organ, or Organ Component|General Exam|5556,5565|false|false|false|C0030647|Patella|knee caps
Disorder|Disease or Syndrome|General Exam|5561,5565|false|false|false|C2316212;C3662487|Catastrophic antiphospholipid syndrome;Cryopyrin-Associated Periodic Syndromes|caps
Drug|Biomedical or Dental Material|General Exam|5561,5565|false|false|false|C0006935|capsule (pharmacologic)|caps
Event|Event|General Exam|5561,5565|false|false|false|||caps
Finding|Gene or Genome|General Exam|5561,5565|false|false|false|C1413079;C1413120|CADPS gene;CAPS gene|caps
Attribute|Clinical Attribute|General Exam|5577,5583|false|false|false|C5889824||status
Finding|Idea or Concept|General Exam|5577,5583|false|false|false|C1546481|What subject filter - Status|status
Disorder|Disease or Syndrome|General Exam|5584,5594|false|false|false|C0011603|Dermatitis|dermatitis
Event|Event|General Exam|5584,5594|false|false|false|||dermatitis
Anatomy|Body System|General Exam|5597,5601|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|General Exam|5597,5601|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|General Exam|5597,5601|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|General Exam|5597,5601|false|false|false|||SKIN
Finding|Body Substance|General Exam|5597,5601|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|General Exam|5597,5601|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Event|Event|General Exam|5603,5612|false|false|false|||Eccymosis
Event|Event|General Exam|5613,5618|false|false|false|||noted
Finding|Functional Concept|General Exam|5622,5626|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|General Exam|5622,5631|false|false|false|C0230371|Structure of left hand|left hand
Anatomy|Body Part, Organ, or Organ Component|General Exam|5627,5631|false|false|false|C0018563;C4285005|Hand;Upper extremity>Hand|hand
Finding|Finding|General Exam|5627,5631|false|false|false|C0741992|Hand problem|hand
Procedure|Diagnostic Procedure|General Exam|5642,5653|false|false|false|C0184922||open biopsy
Event|Event|General Exam|5647,5653|false|false|false|||biopsy
Finding|Finding|General Exam|5647,5653|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Finding|Intellectual Product|General Exam|5647,5653|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Procedure|Diagnostic Procedure|General Exam|5647,5653|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Procedure|Health Care Activity|General Exam|5647,5653|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Event|Event|General Exam|5655,5663|false|false|false|||excision
Procedure|Therapeutic or Preventive Procedure|General Exam|5655,5663|false|false|false|C0015252;C0728940|Excision;removal technique|excision
Finding|Functional Concept|General Exam|5673,5677|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|General Exam|5673,5682|false|false|false|C0817700|Anterior part of left leg|left shin
Anatomy|Body Location or Region|General Exam|5678,5682|false|false|false|C0230444|Shin|shin
Finding|Functional Concept|General Exam|5687,5692|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|General Exam|5687,5697|false|false|false|C0489801|Posterior part of right leg|right calf
Anatomy|Body Location or Region|General Exam|5693,5697|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|General Exam|5693,5697|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Drug|Food|General Exam|5698,5704|false|false|false|C5890763||PULSES
Event|Event|General Exam|5698,5704|false|false|false|||PULSES
Finding|Physiologic Function|General Exam|5698,5704|false|false|false|C0391850|Physiologic pulse|PULSES
Procedure|Health Care Activity|General Exam|5698,5704|false|false|false|C0034107|Pulse taking|PULSES
Attribute|Clinical Attribute|General Exam|5706,5712|false|false|false|C4522154|Distal Resection Margin|Distal
Drug|Food|General Exam|5713,5719|false|false|false|C5890763||pulses
Event|Event|General Exam|5713,5719|false|false|false|||pulses
Finding|Physiologic Function|General Exam|5713,5719|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|5713,5719|false|false|false|C0034107|Pulse taking|pulses
Event|Event|General Exam|5733,5742|false|false|false|||symmetric
Finding|Conceptual Entity|General Exam|5733,5742|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|General Exam|5733,5742|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Event|Event|General Exam|5746,5755|false|false|false|||Discharge
Finding|Body Substance|General Exam|5746,5755|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|General Exam|5746,5755|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|General Exam|5746,5755|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|General Exam|5746,5755|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|General Exam|5756,5764|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|General Exam|5756,5764|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|General Exam|5756,5764|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|General Exam|5756,5769|false|false|false|C1509143|physical examination (physical finding)|Physical exam
Procedure|Health Care Activity|General Exam|5756,5769|false|false|false|C0031809|Physical Examination|Physical exam
Event|Event|General Exam|5765,5769|false|false|false|||exam
Finding|Functional Concept|General Exam|5765,5769|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|General Exam|5765,5769|false|false|false|C0582103|Medical Examination|exam
Event|Event|General Exam|5800,5804|false|false|false|||Data
Finding|Idea or Concept|General Exam|5800,5804|false|false|false|C1511726|Data|Data
Event|Event|General Exam|5811,5818|false|false|false|||updated
Event|Event|General Exam|5834,5838|false|false|false|||Temp
Finding|Gene or Genome|General Exam|5834,5838|false|false|false|C1823816|C1orf210 gene|Temp
Procedure|Therapeutic or Preventive Procedure|General Exam|5834,5838|false|false|false|C0279848|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Temp
Event|Event|General Exam|5938,5946|false|false|false|||delivery
Finding|Finding|General Exam|5938,5946|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Finding|Functional Concept|General Exam|5938,5946|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Finding|Organism Function|General Exam|5938,5946|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Procedure|Therapeutic or Preventive Procedure|General Exam|5938,5946|false|false|false|C0011209|Obstetric Delivery|delivery
Event|Event|General Exam|5954,5961|false|false|false|||General
Finding|Classification|General Exam|5954,5961|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|General Exam|5954,5961|false|false|false|C3812897|General medical service|General
Event|Event|General Exam|5971,5980|false|false|false|||gentleman
Disorder|Disease or Syndrome|General Exam|5984,5987|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|5984,5987|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|5984,5987|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|5984,5987|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|5984,5987|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|General Exam|5984,5987|false|false|false|||NAD
Finding|Finding|General Exam|5984,5987|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|General Exam|5988,5993|false|false|false|C1512338|HEENT|HEENT
Drug|Biomedical or Dental Material|General Exam|5995,6003|false|false|false|C1705365|Dressing Dosage Form|dressing
Event|Event|General Exam|5995,6003|false|false|false|||dressing
Finding|Daily or Recreational Activity|General Exam|5995,6003|false|false|false|C0518459;C1305428|Ability to dress|dressing
Finding|Finding|General Exam|5995,6003|false|false|false|C0518459;C1305428|Ability to dress|dressing
Procedure|Health Care Activity|General Exam|5995,6003|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Procedure|Therapeutic or Preventive Procedure|General Exam|5995,6003|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Event|Activity|General Exam|6007,6012|false|false|false|C1882509|put - instruction imperative|place
Event|Event|General Exam|6007,6012|false|false|false|||place
Finding|Functional Concept|General Exam|6007,6012|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|General Exam|6007,6012|false|false|false|C1533810||place
Anatomy|Body Part, Organ, or Organ Component|General Exam|6016,6021|false|false|false|C0036270|Scalp structure|scalp
Event|Event|General Exam|6034,6038|false|false|false|||fall
Finding|Finding|General Exam|6034,6038|false|false|false|C0085639|Falls|fall
Anatomy|Body Part, Organ, or Organ Component|General Exam|6039,6044|false|false|false|C0036270|Scalp structure|scalp
Disorder|Injury or Poisoning|General Exam|6045,6055|false|false|false|C0043246|Laceration|laceration
Event|Event|General Exam|6045,6055|false|false|false|||laceration
Anatomy|Body Part, Organ, or Organ Component|General Exam|6063,6069|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|General Exam|6063,6069|false|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|General Exam|6063,6069|false|false|false|||Sclera
Procedure|Health Care Activity|General Exam|6063,6069|false|false|false|C2228481|examination of sclera|Sclera
Event|Event|General Exam|6077,6084|false|false|false|||icteric
Finding|Sign or Symptom|General Exam|6077,6084|false|false|false|C0022346|Icterus|icteric
Anatomy|Body Part, Organ, or Organ Component|General Exam|6086,6092|false|false|false|C0034121|Pupil|pupils
Anatomy|Body Part, Organ, or Organ Component|General Exam|6108,6111|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|General Exam|6108,6111|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Location or Region|General Exam|6113,6117|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|General Exam|6113,6117|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|General Exam|6113,6117|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|General Exam|6119,6122|false|false|false|||JVP
Finding|Finding|General Exam|6119,6122|false|false|false|C0428897|Jugular venous pressure|JVP
Disorder|Cell or Molecular Dysfunction|General Exam|6134,6142|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Event|Event|General Exam|6134,6142|false|false|false|||positive
Finding|Classification|General Exam|6134,6142|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|General Exam|6134,6142|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|General Exam|6143,6163|false|false|false|C5784512|Hepatojugular Reflex|hepatojugular reflex
Event|Event|General Exam|6157,6163|false|false|false|||reflex
Finding|Finding|General Exam|6157,6163|false|false|false|C0034929;C0439840;C0596002|Observation of reflex;Reflex action;Reflex motion descriptor|reflex
Finding|Organ or Tissue Function|General Exam|6157,6163|false|false|false|C0034929;C0439840;C0596002|Observation of reflex;Reflex action;Reflex motion descriptor|reflex
Event|Event|General Exam|6181,6190|false|false|false|||irregular
Anatomy|Body Location or Region|General Exam|6197,6207|true|false|false|C0230134|Structure of precordium|precordium
Event|Event|General Exam|6211,6216|true|false|false|||quiet
Event|Event|General Exam|6225,6227|true|false|false|||RV
Disorder|Disease or Syndrome|General Exam|6228,6233|true|false|false|C3714496|Chronic obstructive pulmonary disease of horses|heave
Event|Event|General Exam|6228,6233|true|false|false|||heave
Finding|Functional Concept|General Exam|6256,6261|false|false|false|C1534709|Splitting|split
Finding|Finding|General Exam|6256,6264|false|false|false|C0425619|Second heart sound split|split S2
Disorder|Disease or Syndrome|General Exam|6277,6281|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|General Exam|6277,6281|false|false|false|||soft
Event|Event|General Exam|6299,6305|false|false|false|||murmur
Finding|Finding|General Exam|6299,6305|false|false|false|C0018808|Heart murmur|murmur
Anatomy|Cell Component|General Exam|6326,6330|false|false|false|C3890171|dinoflagellate apex|apex
Drug|Amino Acid, Peptide, or Protein|General Exam|6326,6330|false|false|false|C0140145|APEX1 protein, human|apex
Drug|Enzyme|General Exam|6326,6330|false|false|false|C0140145|APEX1 protein, human|apex
Finding|Gene or Genome|General Exam|6326,6330|false|false|false|C1332102|APEX1 gene|apex
Anatomy|Body Part, Organ, or Organ Component|General Exam|6332,6337|false|false|false|C0024109|Lung|LUNGS
Event|Event|General Exam|6346,6352|false|false|false|||effort
Finding|Organism Function|General Exam|6346,6352|false|false|false|C0015264|Exertion|effort
Event|Event|General Exam|6369,6377|false|false|false|||crackles
Finding|Finding|General Exam|6369,6377|false|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Anatomy|Body Location or Region|General Exam|6378,6381|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|Abd
Disorder|Cell or Molecular Dysfunction|General Exam|6378,6381|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|Abd
Disorder|Disease or Syndrome|General Exam|6383,6387|true|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|General Exam|6383,6387|true|false|false|||soft
Event|Event|General Exam|6395,6404|true|false|false|||distended
Finding|Finding|General Exam|6395,6404|true|false|false|C0700124|Dilated|distended
Event|Event|General Exam|6409,6417|true|false|false|||guarding
Finding|Finding|General Exam|6409,6417|true|false|false|C0427198|Protective muscle spasm|guarding
Disorder|Congenital Abnormality|General Exam|6430,6433|false|false|false|C0015306|Hereditary Multiple Exostoses|EXT
Event|Event|General Exam|6430,6433|false|false|false|||EXT
Finding|Gene or Genome|General Exam|6430,6433|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|EXT
Finding|Finding|General Exam|6436,6452|false|false|false|C1720243|1+ pitting edema|1+ pitting edema
Finding|Functional Concept|General Exam|6439,6446|false|false|false|C0205323|Pitting|pitting
Finding|Finding|General Exam|6439,6452|false|false|false|C0333243|Pitting edema|pitting edema
Attribute|Clinical Attribute|General Exam|6447,6452|false|false|false|C1717255||edema
Event|Event|General Exam|6447,6452|false|false|false|||edema
Finding|Pathologic Function|General Exam|6447,6452|false|false|false|C0013604|Edema|edema
Anatomy|Body Part, Organ, or Organ Component|General Exam|6471,6474|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Anatomy|Body Part, Organ, or Organ Component|General Exam|6479,6482|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Anatomy|Body System|General Exam|6483,6487|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|General Exam|6483,6487|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|General Exam|6483,6487|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|General Exam|6483,6487|false|false|false|||SKIN
Finding|Body Substance|General Exam|6483,6487|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|General Exam|6483,6487|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Procedure|Therapeutic or Preventive Procedure|General Exam|6499,6507|false|false|false|C0015252;C0728940|Excision;removal technique|excision
Procedure|Diagnostic Procedure|General Exam|6499,6514|false|false|false|C0184921|Excision biopsy|excision biopsy
Event|Event|General Exam|6508,6514|false|false|false|||biopsy
Finding|Finding|General Exam|6508,6514|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Finding|Intellectual Product|General Exam|6508,6514|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Procedure|Diagnostic Procedure|General Exam|6508,6514|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Procedure|Health Care Activity|General Exam|6508,6514|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Disorder|Injury or Poisoning|General Exam|6515,6521|false|false|false|C0043250|Traumatic Wound|wounds
Event|Event|General Exam|6515,6521|false|false|false|||wounds
Anatomy|Body Part, Organ, or Organ Component|General Exam|6525,6529|false|false|false|C1140621|Leg|legs
Attribute|Clinical Attribute|General Exam|6525,6529|false|false|false|C5781420||legs
Event|Event|General Exam|6531,6538|false|false|false|||covered
Drug|Biomedical or Dental Material|General Exam|6544,6552|false|false|false|C1705365|Dressing Dosage Form|dressing
Event|Event|General Exam|6544,6552|false|false|false|||dressing
Finding|Daily or Recreational Activity|General Exam|6544,6552|false|false|false|C0518459;C1305428|Ability to dress|dressing
Finding|Finding|General Exam|6544,6552|false|false|false|C0518459;C1305428|Ability to dress|dressing
Procedure|Health Care Activity|General Exam|6544,6552|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Procedure|Therapeutic or Preventive Procedure|General Exam|6544,6552|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Event|Event|General Exam|6567,6573|false|false|false|||Speech
Finding|Organism Function|General Exam|6567,6573|false|false|false|C0037817|Speech|Speech
Procedure|Diagnostic Procedure|General Exam|6567,6573|false|false|false|C0846595|Speech assessment|Speech
Event|Event|General Exam|6582,6590|false|false|false|||strength
Finding|Idea or Concept|General Exam|6582,6590|false|false|false|C0808080|Strength (attribute)|strength
Event|Event|General Exam|6599,6605|false|false|false|||intact
Finding|Finding|General Exam|6599,6605|false|false|false|C1554187|Gender Status - Intact|intact
Disorder|Neoplastic Process|General Exam|6647,6650|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|General Exam|6647,6650|false|false|false|||PTT
Procedure|Laboratory Procedure|General Exam|6647,6650|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Event|Event|General Exam|6674,6677|false|false|false|||PLT
Procedure|Laboratory Procedure|General Exam|6674,6677|false|false|false|C0201617|Primed lymphocyte test|PLT
Event|Event|General Exam|6702,6707|false|false|false|||NEUTS
Finding|Body Substance|General Exam|6714,6720|false|false|false|C0024202|Lymph|LYMPHS
Drug|Antibiotic|General Exam|6726,6731|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Biomedical or Dental Material|General Exam|6726,6731|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Organic Chemical|General Exam|6726,6731|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Disorder|Disease or Syndrome|General Exam|6737,6740|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|EOS
Event|Event|General Exam|6737,6740|false|false|false|||EOS
Finding|Gene or Genome|General Exam|6737,6740|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|EOS
Anatomy|Cell|General Exam|6845,6848|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|6853,6856|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|6853,6856|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|6853,6856|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|6863,6866|false|false|false|C0019046|Hemoglobin|HGB
Drug|Biologically Active Substance|General Exam|6863,6866|false|false|false|C0019046|Hemoglobin|HGB
Event|Event|General Exam|6863,6866|false|false|false|||HGB
Finding|Gene or Genome|General Exam|6863,6866|false|false|false|C1424337|CYGB gene|HGB
Lab|Laboratory or Test Result|General Exam|6863,6866|false|false|false|C0019029|Hemoglobin concentration|HGB
Event|Event|General Exam|6872,6875|false|false|false|||HCT
Procedure|Laboratory Procedure|General Exam|6872,6875|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|General Exam|6872,6875|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Disorder|Virus|General Exam|6882,6885|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|General Exam|6882,6885|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|6882,6885|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|6882,6885|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|6892,6895|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|6892,6895|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|6892,6895|false|false|false|||MCH
Finding|Gene or Genome|General Exam|6892,6895|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|6892,6895|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|6892,6895|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|6901,6905|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|6901,6905|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Drug|Amino Acid, Peptide, or Protein|General Exam|6960,6968|false|false|false|C0015879|Ferritin|FERRITIN
Drug|Biologically Active Substance|General Exam|6960,6968|false|false|false|C0015879|Ferritin|FERRITIN
Drug|Pharmacologic Substance|General Exam|6960,6968|false|false|false|C0015879|Ferritin|FERRITIN
Event|Event|General Exam|6960,6968|false|false|false|||FERRITIN
Procedure|Laboratory Procedure|General Exam|6960,6968|false|false|false|C0373607|Ferritin measurement|FERRITIN
Drug|Amino Acid, Peptide, or Protein|General Exam|6973,6976|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Biologically Active Substance|General Exam|6973,6976|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Hormone|General Exam|6973,6976|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Pharmacologic Substance|General Exam|6973,6976|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Event|Event|General Exam|6973,6976|false|false|false|||TRF
Finding|Gene or Genome|General Exam|6973,6976|false|false|false|C1334121;C1336604;C1705002|IL5 gene;TERF1 gene;TERF1 wt Allele|TRF
Drug|Biologically Active Substance|General Exam|6995,7002|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Element, Ion, or Isotope|General Exam|6995,7002|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Inorganic Chemical|General Exam|6995,7002|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Pharmacologic Substance|General Exam|6995,7002|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Vitamin|General Exam|6995,7002|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Event|Event|General Exam|6995,7002|false|false|false|||CALCIUM
Finding|Physiologic Function|General Exam|6995,7002|false|false|false|C4553026|Calcium metabolic function|CALCIUM
Procedure|Laboratory Procedure|General Exam|6995,7002|false|false|false|C0201925|Calcium measurement|CALCIUM
Drug|Element, Ion, or Isotope|General Exam|7007,7016|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Drug|Inorganic Chemical|General Exam|7007,7016|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Drug|Pharmacologic Substance|General Exam|7007,7016|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Procedure|Laboratory Procedure|General Exam|7007,7016|false|false|false|C0523826|Phosphate measurement|PHOSPHATE
Drug|Biologically Active Substance|General Exam|7021,7030|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Element, Ion, or Isotope|General Exam|7021,7030|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Inorganic Chemical|General Exam|7021,7030|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Pharmacologic Substance|General Exam|7021,7030|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Procedure|Laboratory Procedure|General Exam|7021,7030|false|false|false|C0373675|Magnesium measurement|MAGNESIUM
Drug|Biologically Active Substance|General Exam|7037,7041|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|IRON
Drug|Element, Ion, or Isotope|General Exam|7037,7041|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|IRON
Drug|Pharmacologic Substance|General Exam|7037,7041|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|IRON
Event|Event|General Exam|7037,7041|false|false|false|||IRON
Procedure|Laboratory Procedure|General Exam|7037,7041|false|false|false|C0337439|Iron measurement|IRON
Drug|Amino Acid, Peptide, or Protein|General Exam|7059,7064|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|General Exam|7059,7064|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|General Exam|7059,7064|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|General Exam|7059,7064|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Disorder|Neoplastic Process|General Exam|7098,7101|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|7098,7101|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|General Exam|7098,7101|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|General Exam|7098,7101|false|false|false|||ALT
Finding|Gene or Genome|General Exam|7098,7101|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|General Exam|7098,7101|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|General Exam|7098,7101|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|General Exam|7098,7101|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|7102,7106|false|false|false|C0376147|SGPT - Glutamate pyruvate transaminase|SGPT
Drug|Enzyme|General Exam|7102,7106|false|false|false|C0376147|SGPT - Glutamate pyruvate transaminase|SGPT
Event|Event|General Exam|7102,7106|false|false|false|||SGPT
Finding|Gene or Genome|General Exam|7102,7106|false|false|false|C1415274|GPT gene|SGPT
Procedure|Laboratory Procedure|General Exam|7102,7106|false|false|false|C0036828|Serum Alanine Transaminase Test|SGPT
Anatomy|Body Space or Junction|General Exam|7112,7115|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|General Exam|7112,7115|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|7112,7115|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|General Exam|7112,7115|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|General Exam|7112,7115|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|General Exam|7112,7115|false|false|false|||AST
Finding|Gene or Genome|General Exam|7112,7115|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|7116,7120|false|false|false|C0242192|SGOT - Glutamate oxaloacetate transaminase|SGOT
Drug|Enzyme|General Exam|7116,7120|false|false|false|C0242192|SGOT - Glutamate oxaloacetate transaminase|SGOT
Event|Event|General Exam|7116,7120|false|false|false|||SGOT
Finding|Gene or Genome|General Exam|7116,7120|false|false|false|C1415181|GOT1 gene|SGOT
Procedure|Laboratory Procedure|General Exam|7116,7120|false|false|false|C0201899|Aspartate aminotransferase measurement|SGOT
Drug|Amino Acid, Peptide, or Protein|General Exam|7129,7132|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Drug|Enzyme|General Exam|7129,7132|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Event|Event|General Exam|7129,7132|false|false|false|||LDH
Finding|Finding|General Exam|7129,7132|false|false|false|C0851148|Lifetime Drinking History|LDH
Procedure|Laboratory Procedure|General Exam|7129,7132|false|false|false|C0202113|Lactate dehydrogenase measurement|LDH
Drug|Amino Acid, Peptide, or Protein|General Exam|7139,7142|false|false|false|C1663627|ALK protein, human|ALK
Drug|Enzyme|General Exam|7139,7142|false|false|false|C1663627|ALK protein, human|ALK
Event|Event|General Exam|7139,7142|false|false|false|||ALK
Finding|Gene or Genome|General Exam|7139,7142|false|false|false|C1332080;C1663627;C1704943|ALK gene;ALK protein, human;ALK wt Allele|ALK
Finding|Receptor|General Exam|7139,7142|false|false|false|C1332080;C1663627;C1704943|ALK gene;ALK protein, human;ALK wt Allele|ALK
Event|Event|General Exam|7158,7162|false|false|false|||BILI
Drug|Biologically Active Substance|General Exam|7213,7220|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|General Exam|7213,7220|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|General Exam|7213,7220|false|false|false|C0017725|glucose|GLUCOSE
Event|Event|General Exam|7213,7220|false|false|false|||GLUCOSE
Lab|Laboratory or Test Result|General Exam|7213,7220|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|General Exam|7213,7220|false|false|false|C0337438|Glucose measurement|GLUCOSE
Drug|Biologically Active Substance|General Exam|7225,7229|false|false|false|C0041942|urea|UREA
Drug|Organic Chemical|General Exam|7225,7229|false|false|false|C0041942|urea|UREA
Drug|Pharmacologic Substance|General Exam|7225,7229|false|false|false|C0041942|urea|UREA
Event|Event|General Exam|7225,7229|false|false|false|||UREA
Procedure|Laboratory Procedure|General Exam|7225,7229|false|false|false|C0523961|Urea measurement|UREA
Drug|Biologically Active Substance|General Exam|7247,7253|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Element, Ion, or Isotope|General Exam|7247,7253|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Pharmacologic Substance|General Exam|7247,7253|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Event|Event|General Exam|7247,7253|false|false|false|||SODIUM
Finding|Physiologic Function|General Exam|7247,7253|false|false|false|C4553025|Sodium metabolic function|SODIUM
Procedure|Laboratory Procedure|General Exam|7247,7253|false|false|false|C0337443|Sodium measurement|SODIUM
Drug|Biologically Active Substance|General Exam|7259,7268|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Element, Ion, or Isotope|General Exam|7259,7268|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Food|General Exam|7259,7268|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Inorganic Chemical|General Exam|7259,7268|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Pharmacologic Substance|General Exam|7259,7268|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Event|Event|General Exam|7259,7268|false|false|false|||POTASSIUM
Finding|Physiologic Function|General Exam|7259,7268|false|false|false|C4553027|Potassium metabolic function|POTASSIUM
Procedure|Laboratory Procedure|General Exam|7259,7268|false|false|false|C0202194|Potassium measurement|POTASSIUM
Drug|Element, Ion, or Isotope|General Exam|7273,7281|false|false|false|C0008203;C0596019|Chlorides;chloride ion|CHLORIDE
Event|Event|General Exam|7273,7281|false|false|false|||CHLORIDE
Finding|Physiologic Function|General Exam|7273,7281|false|false|false|C4553021|Chloride metabolic function|CHLORIDE
Procedure|Laboratory Procedure|General Exam|7273,7281|false|false|false|C0201952|Chloride measurement|CHLORIDE
Drug|Biologically Active Substance|General Exam|7292,7295|false|false|false|C0007012|carbon dioxide|CO2
Drug|Inorganic Chemical|General Exam|7292,7295|false|false|false|C0007012|carbon dioxide|CO2
Event|Event|General Exam|7292,7295|false|false|false|||CO2
Finding|Finding|General Exam|7292,7295|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Finding|Gene or Genome|General Exam|7292,7295|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Drug|Element, Ion, or Isotope|General Exam|7299,7304|false|false|false|C0003075|Anions|ANION
Attribute|Clinical Attribute|General Exam|7299,7308|false|false|false|C0003074|Anion Gap|ANION GAP
Lab|Laboratory or Test Result|General Exam|7299,7308|false|false|false|C1509129|Anion gap result|ANION GAP
Procedure|Laboratory Procedure|General Exam|7299,7308|false|false|false|C0201889;C2189246|Anion gap measurement;blood anion gap (lab test)|ANION GAP
Drug|Amino Acid, Peptide, or Protein|General Exam|7305,7308|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Drug|Biologically Active Substance|General Exam|7305,7308|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Event|Event|General Exam|7305,7308|false|false|false|||GAP
Finding|Gene or Genome|General Exam|7305,7308|false|false|false|C1419277;C2984552|RASA1 gene;RASA1 wt Allele|GAP
Finding|Body Substance|General Exam|7324,7329|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|7324,7329|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|7324,7329|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Body Substance|General Exam|7331,7338|false|false|false|C0020191|Hyalin Substance|HYALINE
Finding|Body Substance|General Exam|7354,7359|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|7354,7359|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|7354,7359|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Lab|Laboratory or Test Result|General Exam|7354,7364|false|false|false|C0221752;C2188659|Red blood cells urine positive|URINE  RBC
Anatomy|Cell|General Exam|7361,7364|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|7361,7364|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|7361,7364|false|false|false|C0014792|Erythrocytes|RBC
Anatomy|Cell|General Exam|7367,7370|true|false|false|C0023516|Leukocytes|WBC
Finding|Functional Concept|General Exam|7374,7382|true|false|false|C1510439|bacteria aspects|BACTERIA
Drug|Food|General Exam|7388,7393|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Immunologic Factor|General Exam|7388,7393|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|7388,7393|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Pharmacologic Substance|General Exam|7388,7393|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Event|Event|General Exam|7388,7393|true|false|false|||YEAST
Event|Event|General Exam|7394,7398|true|false|false|||NONE
Disorder|Disease or Syndrome|General Exam|7400,7403|true|false|false|C0267963|Exocrine pancreatic insufficiency|EPI
Drug|Amino Acid, Peptide, or Protein|General Exam|7400,7403|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Biologically Active Substance|General Exam|7400,7403|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Hormone|General Exam|7400,7403|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Organic Chemical|General Exam|7400,7403|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Pharmacologic Substance|General Exam|7400,7403|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Event|Event|General Exam|7400,7403|true|false|false|||EPI
Finding|Gene or Genome|General Exam|7400,7403|true|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|EPI
Finding|Intellectual Product|General Exam|7400,7403|true|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|EPI
Procedure|Diagnostic Procedure|General Exam|7400,7403|true|false|false|C0162734;C3641909|Echo-Planar Imaging;Electronic Portal Imaging|EPI
Finding|Body Substance|General Exam|7419,7424|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|7419,7424|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|7419,7424|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Disorder|Disease or Syndrome|General Exam|7419,7431|false|false|false|C0018965|Hematuria|URINE  BLOOD
Disorder|Disease or Syndrome|General Exam|7426,7431|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|7426,7431|false|false|false|||BLOOD
Finding|Body Substance|General Exam|7426,7431|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Event|General Exam|7432,7435|false|false|false|||NEG
Finding|Finding|General Exam|7432,7435|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|General Exam|7436,7443|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Drug|Inorganic Chemical|General Exam|7436,7443|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Drug|Pharmacologic Substance|General Exam|7436,7443|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Finding|Finding|General Exam|7444,7447|false|false|false|C5848551|Neg - answer|NEG
Drug|Amino Acid, Peptide, or Protein|General Exam|7448,7455|false|false|false|C0033684|Proteins|PROTEIN
Drug|Biologically Active Substance|General Exam|7448,7455|false|false|false|C0033684|Proteins|PROTEIN
Event|Event|General Exam|7448,7455|false|false|false|||PROTEIN
Finding|Conceptual Entity|General Exam|7448,7455|false|false|false|C1521746|Protein Info|PROTEIN
Procedure|Laboratory Procedure|General Exam|7448,7455|false|false|false|C0202202|Protein measurement|PROTEIN
Drug|Biologically Active Substance|General Exam|7461,7468|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|General Exam|7461,7468|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|General Exam|7461,7468|false|false|false|C0017725|glucose|GLUCOSE
Event|Event|General Exam|7461,7468|false|false|false|||GLUCOSE
Lab|Laboratory or Test Result|General Exam|7461,7468|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|General Exam|7461,7468|false|false|false|C0337438|Glucose measurement|GLUCOSE
Event|Event|General Exam|7469,7472|false|false|false|||NEG
Finding|Finding|General Exam|7469,7472|false|false|false|C5848551|Neg - answer|NEG
Drug|Organic Chemical|General Exam|7473,7479|false|false|false|C0022634|Ketones|KETONE
Event|Event|General Exam|7480,7483|false|false|false|||NEG
Finding|Finding|General Exam|7480,7483|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|General Exam|7484,7493|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Drug|Organic Chemical|General Exam|7484,7493|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Drug|Pharmacologic Substance|General Exam|7484,7493|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Procedure|Laboratory Procedure|General Exam|7484,7493|false|false|false|C0201913;C0863174|Bilirubin, total measurement;blood bilirubin level test|BILIRUBIN
Event|Event|General Exam|7494,7497|false|false|false|||NEG
Finding|Finding|General Exam|7494,7497|false|false|false|C5848551|Neg - answer|NEG
Event|Event|General Exam|7508,7511|false|false|false|||NEG
Finding|Finding|General Exam|7508,7511|false|false|false|C5848551|Neg - answer|NEG
Event|Event|General Exam|7525,7528|false|false|false|||NEG
Finding|Finding|General Exam|7525,7528|false|false|false|C5848551|Neg - answer|NEG
Finding|Body Substance|General Exam|7541,7546|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|7541,7546|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|7541,7546|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Finding|General Exam|7541,7553|false|false|false|C0278030|Color of urine|URINE  COLOR
Drug|Biomedical or Dental Material|General Exam|7548,7553|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|COLOR
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|7548,7553|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|COLOR
Event|Event|General Exam|7548,7553|false|false|false|||COLOR
Drug|Organic Chemical|General Exam|7554,7559|false|false|false|C4047917|Cereal plant straw|Straw
Event|Event|General Exam|7567,7572|false|false|false|||Clear
Finding|Idea or Concept|General Exam|7567,7572|false|false|false|C1550016|Remote control command - Clear|Clear
Disorder|Disease or Syndrome|General Exam|7592,7597|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|7592,7597|false|false|false|||BLOOD
Finding|Body Substance|General Exam|7592,7597|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|7598,7601|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|7606,7609|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|7606,7609|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|7606,7609|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|7616,7619|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|7616,7619|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|7616,7619|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|7616,7619|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|7625,7628|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|7625,7628|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|7636,7639|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|7636,7639|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|7636,7639|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|7636,7639|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|7636,7639|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|7643,7646|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|7643,7646|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|7643,7646|false|false|false|||MCH
Finding|Gene or Genome|General Exam|7643,7646|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|7643,7646|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|7643,7646|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|7652,7656|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|7652,7656|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|7685,7688|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|7705,7710|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|7705,7710|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|7711,7714|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|7731,7736|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|7731,7736|false|false|false|||BLOOD
Finding|Body Substance|General Exam|7731,7736|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|7731,7744|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|7731,7744|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|7731,7744|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|7737,7744|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|7737,7744|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|7737,7744|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|7737,7744|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|7737,7744|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|7737,7744|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|7792,7796|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|7792,7796|false|false|false|C0005367|Bicarbonates|HCO3
Event|Event|General Exam|7792,7796|false|false|false|||HCO3
Procedure|Laboratory Procedure|General Exam|7792,7796|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|7818,7823|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|7818,7823|false|false|false|||BLOOD
Finding|Body Substance|General Exam|7818,7823|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|7824,7827|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|7824,7827|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|General Exam|7824,7827|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|General Exam|7824,7827|false|false|false|||ALT
Finding|Gene or Genome|General Exam|7824,7827|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|General Exam|7824,7827|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|General Exam|7824,7827|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|General Exam|7824,7827|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|General Exam|7832,7835|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|General Exam|7832,7835|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|7832,7835|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|General Exam|7832,7835|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|General Exam|7832,7835|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|General Exam|7832,7835|false|false|false|||AST
Finding|Gene or Genome|General Exam|7832,7835|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|7840,7847|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|General Exam|7840,7847|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|General Exam|7876,7881|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|7876,7881|false|false|false|||BLOOD
Finding|Body Substance|General Exam|7876,7881|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|7876,7889|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|General Exam|7882,7889|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|7882,7889|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|7882,7889|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|7882,7889|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|7882,7889|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|General Exam|7882,7889|false|false|false|||Calcium
Finding|Physiologic Function|General Exam|7882,7889|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|7882,7889|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|General Exam|7922,7927|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|7922,7927|false|false|false|||BLOOD
Finding|Body Substance|General Exam|7922,7927|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|7952,7955|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Biologically Active Substance|General Exam|7952,7955|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Hormone|General Exam|7952,7955|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Pharmacologic Substance|General Exam|7952,7955|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Event|Event|General Exam|7952,7955|false|false|false|||TRF
Finding|Gene or Genome|General Exam|7952,7955|false|false|false|C1334121;C1336604;C1705002|IL5 gene;TERF1 gene;TERF1 wt Allele|TRF
Finding|Idea or Concept|Hospital Course|7985,7997|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Finding|Body Substance|Hospital Course|8028,8037|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|Hospital Course|8028,8037|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|Hospital Course|8028,8037|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|Hospital Course|8028,8037|false|false|false|C0030685|Patient Discharge|DISCHARGE
Attribute|Clinical Attribute|Hospital Course|8038,8044|false|false|false|C0944911||WEIGHT
Event|Event|Hospital Course|8038,8044|false|false|false|||WEIGHT
Finding|Finding|Hospital Course|8038,8044|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|WEIGHT
Finding|Sign or Symptom|Hospital Course|8038,8044|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|WEIGHT
Procedure|Health Care Activity|Hospital Course|8038,8044|false|false|false|C1305866|Weighing patient|WEIGHT
Finding|Body Substance|Hospital Course|8067,8076|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|Hospital Course|8067,8076|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|Hospital Course|8067,8076|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|Hospital Course|8067,8076|false|false|false|C0030685|Patient Discharge|DISCHARGE
Drug|Biologically Active Substance|Hospital Course|8080,8083|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Drug|Inorganic Chemical|Hospital Course|8080,8083|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Event|Event|Hospital Course|8080,8083|false|false|false|||BUN
Procedure|Laboratory Procedure|Hospital Course|8080,8083|false|false|false|C0005845|Blood urea nitrogen measurement|BUN
Drug|Biologically Active Substance|Hospital Course|8093,8096|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Drug|Inorganic Chemical|Hospital Course|8093,8096|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Event|Event|Hospital Course|8093,8096|false|false|false|||BUN
Procedure|Laboratory Procedure|Hospital Course|8093,8096|false|false|false|C0005845|Blood urea nitrogen measurement|BUN
Finding|Body Substance|Hospital Course|8100,8109|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|Hospital Course|8100,8109|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|Hospital Course|8100,8109|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|Hospital Course|8100,8109|false|false|false|C0030685|Patient Discharge|DISCHARGE
Drug|Pharmacologic Substance|Hospital Course|8110,8118|false|false|false|C0012798;C5399719|Diuretic [APC];Diuretics|DIURETIC
Event|Event|Hospital Course|8110,8118|false|false|false|||DIURETIC
Drug|Organic Chemical|Hospital Course|8123,8132|false|false|false|C0076840|torsemide|Torsemide
Drug|Pharmacologic Substance|Hospital Course|8123,8132|false|false|false|C0076840|torsemide|Torsemide
Drug|Pharmacologic Substance|Hospital Course|8139,8149|false|false|false|C0013227|Pharmaceutical Preparations|MEDICATION
Event|Event|Hospital Course|8139,8149|false|false|false|||MEDICATION
Finding|Intellectual Product|Hospital Course|8139,8149|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|MEDICATION
Event|Event|Hospital Course|8150,8157|false|false|false|||CHANGES
Finding|Functional Concept|Hospital Course|8150,8157|false|false|false|C0392747|Changing|CHANGES
Event|Event|Hospital Course|8159,8168|false|false|false|||Decreased
Drug|Biologically Active Substance|Hospital Course|8175,8184|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Element, Ion, or Isotope|Hospital Course|8175,8184|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Food|Hospital Course|8175,8184|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Inorganic Chemical|Hospital Course|8175,8184|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Pharmacologic Substance|Hospital Course|8175,8184|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Event|Event|Hospital Course|8175,8184|false|false|false|||potassium
Finding|Physiologic Function|Hospital Course|8175,8184|false|false|false|C4553027|Potassium metabolic function|potassium
Procedure|Laboratory Procedure|Hospital Course|8175,8184|false|false|false|C0202194|Potassium measurement|potassium
Finding|Functional Concept|Hospital Course|8247,8253|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Event|Event|Hospital Course|8254,8260|false|false|false|||Chem10
Drug|Inorganic Chemical|Hospital Course|8303,8314|false|false|false|C0013832;C3536863|Electrolyte [EPC];Electrolytes|electrolyte
Drug|Pharmacologic Substance|Hospital Course|8303,8314|false|false|false|C0013832;C3536863|Electrolyte [EPC];Electrolytes|electrolyte
Event|Event|Hospital Course|8315,8324|false|false|false|||repletion
Event|Event|Hospital Course|8348,8354|false|false|false|||follow
Attribute|Clinical Attribute|Hospital Course|8358,8364|false|false|false|C0944911||weight
Event|Event|Hospital Course|8358,8364|false|false|false|||weight
Finding|Finding|Hospital Course|8358,8364|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|Hospital Course|8358,8364|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|Hospital Course|8358,8364|false|false|false|C1305866|Weighing patient|weight
Finding|Intellectual Product|Hospital Course|8369,8375|false|false|false|C1705102|Volume (publication)|volume
Attribute|Clinical Attribute|Hospital Course|8376,8382|false|false|false|C5889824||status
Event|Event|Hospital Course|8376,8382|false|false|false|||status
Finding|Idea or Concept|Hospital Course|8376,8382|false|false|false|C1546481|What subject filter - Status|status
Event|Event|Hospital Course|8387,8393|false|false|false|||adjust
Drug|Organic Chemical|Hospital Course|8395,8404|false|false|false|C0076840|torsemide|torsemide
Drug|Pharmacologic Substance|Hospital Course|8395,8404|false|false|false|C0076840|torsemide|torsemide
Event|Event|Hospital Course|8395,8404|false|false|false|||torsemide
Event|Event|Hospital Course|8421,8425|false|false|false|||CODE
Event|Occupational Activity|Hospital Course|8421,8425|false|false|false|C0009219|Coding|CODE
Finding|Intellectual Product|Hospital Course|8421,8425|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|CODE
Procedure|Health Care Activity|Hospital Course|8421,8432|false|false|false|C0742531|CODE STATUS|CODE STATUS
Attribute|Clinical Attribute|Hospital Course|8426,8432|false|false|false|C5889824||STATUS
Event|Event|Hospital Course|8426,8432|false|false|false|||STATUS
Finding|Idea or Concept|Hospital Course|8426,8432|false|false|false|C1546481|What subject filter - Status|STATUS
Finding|Idea or Concept|Hospital Course|8448,8454|false|false|false|C0018684|Health|Health
Procedure|Health Care Activity|Hospital Course|8448,8459|false|false|false|C0086388|Health Care|Health care
Event|Activity|Hospital Course|8455,8459|false|false|false|C1947933|care activity|care
Event|Event|Hospital Course|8455,8459|false|false|false|||care
Finding|Finding|Hospital Course|8455,8459|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Hospital Course|8455,8459|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Hospital Course|8460,8465|false|false|false|C3897813|Advance Directive - Proxy|proxy
Event|Event|Hospital Course|8466,8472|false|false|false|||chosen
Finding|Finding|Hospital Course|8474,8477|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Gene or Genome|Hospital Course|8474,8477|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Idea or Concept|Hospital Course|8474,8477|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Intellectual Product|Hospital Course|8474,8477|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Event|Event|Hospital Course|8479,8483|false|false|false|||Name
Finding|Intellectual Product|Hospital Course|8479,8483|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Finding|Idea or Concept|Hospital Course|8487,8493|false|false|false|C0018684|Health|health
Procedure|Health Care Activity|Hospital Course|8487,8498|false|false|false|C0086388|Health Care|health care
Event|Activity|Hospital Course|8494,8498|false|false|false|C1947933|care activity|care
Event|Event|Hospital Course|8494,8498|false|false|false|||care
Finding|Finding|Hospital Course|8494,8498|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Hospital Course|8494,8498|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Hospital Course|8499,8504|false|false|false|C3897813|Advance Directive - Proxy|proxy
Finding|Gene or Genome|Hospital Course|8516,8519|false|false|false|C1420310|SON gene|son
Finding|Idea or Concept|Hospital Course|8521,8526|false|false|false|C1515258;C1547567;C1548343;C1576870|Authorization Mode - Phone;MDFAttributeType - Phone;Telephone Number;Visit User Code - Phone|Phone
Finding|Intellectual Product|Hospital Course|8521,8526|false|false|false|C1515258;C1547567;C1548343;C1576870|Authorization Mode - Phone;MDFAttributeType - Phone;Telephone Number;Visit User Code - Phone|Phone
Finding|Intellectual Product|Hospital Course|8521,8533|false|false|false|C1515258|Telephone Number|Phone number
Event|Event|Hospital Course|8527,8533|false|false|false|||number
Finding|Idea or Concept|Hospital Course|8527,8533|false|false|false|C1554106|MDF AttributeType - Number|number
Finding|Body Substance|Hospital Course|8563,8570|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|PATIENT
Finding|Idea or Concept|Hospital Course|8563,8570|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|PATIENT
Finding|Intellectual Product|Hospital Course|8563,8570|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|PATIENT
Finding|Intellectual Product|Hospital Course|8563,8578|false|false|false|C2964278|Patient summary|PATIENT SUMMARY
Finding|Intellectual Product|Hospital Course|8571,8578|false|false|false|C1552616;C1706244|Summary (document);summary - ActRelationshipSubset|SUMMARY
Event|Event|Hospital Course|8635,8639|false|false|false|||PMHx
Disorder|Disease or Syndrome|Hospital Course|8643,8646|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8643,8646|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|8643,8646|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Hospital Course|8643,8646|false|false|false|||CAD
Finding|Gene or Genome|Hospital Course|8643,8646|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|8643,8646|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|8643,8646|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8643,8646|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|Hospital Course|8652,8656|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8652,8656|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8672,8675|false|false|false|C2713669|SERPINA5 protein, human|PCI
Drug|Biologically Active Substance|Hospital Course|8672,8675|false|false|false|C2713669|SERPINA5 protein, human|PCI
Event|Event|Hospital Course|8672,8675|false|false|false|||PCI
Finding|Gene or Genome|Hospital Course|8672,8675|false|false|false|C1418370;C1705930;C4049621|Peritoneal Cancer Index;SERPINA5 gene;SERPINA5 wt Allele|PCI
Finding|Intellectual Product|Hospital Course|8672,8675|false|false|false|C1418370;C1705930;C4049621|Peritoneal Cancer Index;SERPINA5 gene;SERPINA5 wt Allele|PCI
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8672,8675|false|false|false|C1514496;C1532338;C4724254|Percutaneous Coronary Intervention;Prophylactic Cranial Irradiation;photochemical internalization|PCI
Finding|Finding|Hospital Course|8693,8701|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|Hospital Course|8693,8701|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Event|Event|Hospital Course|8702,8711|false|false|false|||tricuspid
Event|Event|Hospital Course|8712,8725|false|false|false|||regurgitation
Finding|Finding|Hospital Course|8712,8725|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|Hospital Course|8712,8725|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|Hospital Course|8712,8725|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Finding|Functional Concept|Hospital Course|8727,8732|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Finding|Pathologic Function|Hospital Course|8727,8756|false|false|false|C0242707|Right Ventricular Dysfunction|right ventricular dysfunction
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8733,8744|false|false|false|C0018827|Heart Ventricle|ventricular
Finding|Pathologic Function|Hospital Course|8733,8756|false|false|false|C0242973|Ventricular Dysfunction|ventricular dysfunction
Disorder|Disease or Syndrome|Hospital Course|8745,8756|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Event|Event|Hospital Course|8745,8756|false|false|false|||dysfunction
Finding|Conceptual Entity|Hospital Course|8745,8756|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|Hospital Course|8745,8756|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|Hospital Course|8745,8756|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Finding|Hospital Course|8758,8766|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|Hospital Course|8758,8766|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8767,8776|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Hospital Course|8767,8776|false|false|false|C2707265||pulmonary
Finding|Finding|Hospital Course|8767,8776|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Disorder|Disease or Syndrome|Hospital Course|8777,8789|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|Hospital Course|8777,8789|false|false|false|||hypertension
Disorder|Disease or Syndrome|Hospital Course|8795,8825|false|false|false|C0235480|Paroxysmal atrial fibrillation|paroxysmal atrial fibrillation
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8806,8812|false|false|false|C0018792|Heart Atrium|atrial
Attribute|Clinical Attribute|Hospital Course|8806,8825|false|false|false|C2926591||atrial fibrillation
Disorder|Disease or Syndrome|Hospital Course|8806,8825|false|false|false|C0004238|Atrial Fibrillation|atrial fibrillation
Lab|Laboratory or Test Result|Hospital Course|8806,8825|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|atrial fibrillation
Disorder|Disease or Syndrome|Hospital Course|8813,8825|false|false|false|C0232197|Fibrillation|fibrillation
Event|Event|Hospital Course|8813,8825|false|false|false|||fibrillation
Drug|Organic Chemical|Hospital Course|8829,8837|false|false|false|C1831808|apixaban|apixaban
Drug|Pharmacologic Substance|Hospital Course|8829,8837|false|false|false|C1831808|apixaban|apixaban
Event|Event|Hospital Course|8829,8837|false|false|false|||apixaban
Attribute|Clinical Attribute|Hospital Course|8839,8844|false|false|false|C1300072|Tumor stage|stage
Event|Event|Hospital Course|8849,8856|false|false|false|||chronic
Finding|Intellectual Product|Hospital Course|8849,8856|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Hospital Course|8849,8856|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|Hospital Course|8849,8871|false|false|false|C1561643|Chronic Kidney Diseases|chronic kidney disease
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8857,8863|false|false|false|C0022646;C0227665|Both kidneys;Kidney|kidney
Disorder|Neoplastic Process|Hospital Course|8857,8863|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|kidney
Finding|Sign or Symptom|Hospital Course|8857,8863|false|false|false|C0812426|Kidney problem|kidney
Procedure|Diagnostic Procedure|Hospital Course|8857,8863|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8857,8863|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Disorder|Disease or Syndrome|Hospital Course|8857,8871|false|false|false|C0022658|Kidney Diseases|kidney disease
Disorder|Disease or Syndrome|Hospital Course|8864,8871|false|false|false|C0012634|Disease|disease
Event|Event|Hospital Course|8864,8871|false|false|false|||disease
Drug|Biomedical or Dental Material|Hospital Course|8873,8881|false|false|false|C0168634|BaseLine dental cement|Baseline
Finding|Idea or Concept|Hospital Course|8873,8881|false|false|false|C1552824|baseline - TableCellVerticalAlign|Baseline
Disorder|Disease or Syndrome|Hospital Course|8895,8918|false|false|false|C0007820|Cerebrovascular Disorders|cerebrovascular disease
Disorder|Disease or Syndrome|Hospital Course|8911,8918|false|false|false|C0012634|Disease|disease
Event|Event|Hospital Course|8911,8918|false|false|false|||disease
Finding|Functional Concept|Hospital Course|8924,8934|false|false|false|C0036525;C1522484|Metastatic to;metastatic qualifier|metastatic
Disorder|Neoplastic Process|Hospital Course|8924,8943|false|false|false|C0278883|Metastatic melanoma|metastatic melanoma
Disorder|Neoplastic Process|Hospital Course|8935,8943|false|true|false|C0025202|melanoma|melanoma
Drug|Immunologic Factor|Hospital Course|8935,8943|false|true|false|C0796561|Melanoma vaccine|melanoma
Drug|Pharmacologic Substance|Hospital Course|8935,8943|false|true|false|C0796561|Melanoma vaccine|melanoma
Event|Event|Hospital Course|8935,8943|false|false|false|||melanoma
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8947,8954|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Immunologic Factor|Hospital Course|8947,8954|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Pharmacologic Substance|Hospital Course|8947,8954|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Event|Event|Hospital Course|8947,8954|false|false|false|||unknown
Finding|Finding|Hospital Course|8947,8954|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Functional Concept|Hospital Course|8947,8954|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Idea or Concept|Hospital Course|8947,8954|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Intellectual Product|Hospital Course|8947,8954|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Cell Function|Hospital Course|8966,8976|false|false|false|C1155874|Cell Cycle Checkpoints|checkpoint
Drug|Biologically Active Substance|Hospital Course|8977,8986|false|false|false|C1999216|Inhibitor|inhibitor
Event|Event|Hospital Course|8977,8986|false|false|false|||inhibitor
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8987,9000|false|false|false|C3658706|pembrolizumab|pembrolizumab
Drug|Immunologic Factor|Hospital Course|8987,9000|false|false|false|C3658706|pembrolizumab|pembrolizumab
Drug|Pharmacologic Substance|Hospital Course|8987,9000|false|false|false|C3658706|pembrolizumab|pembrolizumab
Event|Event|Hospital Course|8987,9000|false|false|false|||pembrolizumab
Event|Event|Hospital Course|9009,9014|false|false|false|||found
Event|Event|Hospital Course|9015,9021|false|false|false|||volume
Finding|Intellectual Product|Hospital Course|9015,9021|false|false|false|C1705102|Volume (publication)|volume
Event|Event|Hospital Course|9022,9032|false|false|false|||overloaded
Finding|Finding|Hospital Course|9038,9047|false|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Functional Concept|Hospital Course|9038,9047|false|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Event|Event|Hospital Course|9048,9051|false|false|false|||DOE
Finding|Sign or Symptom|Hospital Course|9048,9051|false|false|false|C0231807|Dyspnea on exertion|DOE
Event|Event|Hospital Course|9053,9061|false|false|false|||admitted
Finding|Intellectual Product|Hospital Course|9065,9070|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|Hospital Course|9076,9083|false|false|false|||failure
Finding|Functional Concept|Hospital Course|9076,9083|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|Hospital Course|9076,9083|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|Hospital Course|9076,9083|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|Hospital Course|9091,9099|false|false|false|||diuresis
Finding|Organ or Tissue Function|Hospital Course|9091,9099|false|false|false|C0012797|Diuresis|diuresis
Event|Event|Hospital Course|9105,9117|false|false|false|||transitioned
Anatomy|Body Space or Junction|Hospital Course|9121,9125|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|9121,9125|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|9121,9125|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|9121,9125|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|Hospital Course|9126,9135|false|false|false|||duiretics
Event|Event|Hospital Course|9141,9151|false|false|false|||CORONARIES
Finding|Functional Concept|Hospital Course|9153,9157|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Disorder|Disease or Syndrome|Hospital Course|9167,9194|false|false|false|C0581375|Double coronary vessel disease|two vessel coronary disease
Anatomy|Body Location or Region|Hospital Course|9171,9177|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9171,9177|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9171,9186|false|false|false|C0010075|Coronary Vessels|vessel coronary
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9178,9186|false|false|false|C0018787|Heart|coronary
Disorder|Disease or Syndrome|Hospital Course|9178,9194|false|false|false|C0010068;C1956346|Coronary Artery Disease;Coronary heart disease|coronary disease
Disorder|Disease or Syndrome|Hospital Course|9187,9194|false|false|false|C0012634|Disease|disease
Event|Event|Hospital Course|9187,9194|false|false|false|||disease
Event|Event|Hospital Course|9204,9208|false|false|false|||PUMP
Finding|Molecular Function|Hospital Course|9204,9208|false|false|false|C1150186|matrix metalloproteinase 7 activity|PUMP
Event|Event|Hospital Course|9221,9227|false|false|false|||RHYTHM
Finding|Finding|Hospital Course|9221,9227|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|RHYTHM
Finding|Physiologic Function|Hospital Course|9221,9227|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|RHYTHM
Anatomy|Tissue|Hospital Course|9229,9236|false|false|false|C4050503|Ectopic Graft|Ectopic
Disorder|Disease or Syndrome|Hospital Course|9229,9243|false|false|false|C1399226|Ectopic rhythm|Ectopic rhythm
Event|Event|Hospital Course|9237,9243|false|false|false|||rhythm
Finding|Finding|Hospital Course|9237,9243|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|Hospital Course|9237,9243|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Finding|Hospital Course|9245,9260|false|false|false|C0600125|Prolonged PR interval|PR prolongation
Event|Event|Hospital Course|9248,9260|false|false|false|||prolongation
Finding|Functional Concept|Hospital Course|9262,9266|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Finding|Hospital Course|9262,9281|false|false|false|C0232297|Left axis deviation|left axis deviation
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9267,9271|false|false|false|C0004457|Axis vertebra|axis
Disorder|Injury or Poisoning|Hospital Course|9267,9271|false|false|false|C0349013|Fracture of second cervical vertebra|axis
Finding|Finding|Hospital Course|9267,9281|false|false|false|C0262387|axis deviation|axis deviation
Event|Event|Hospital Course|9272,9281|false|false|false|||deviation
Finding|Finding|Hospital Course|9272,9281|false|false|false|C1705236|Protocol Deviation|deviation
Disorder|Disease or Syndrome|Hospital Course|9284,9288|false|false|false|C0085615|Right bundle branch block|RBBB
Event|Event|Hospital Course|9284,9288|false|false|false|||RBBB
Finding|Finding|Hospital Course|9284,9288|false|false|false|C0344421||RBBB
Event|Event|Hospital Course|9297,9303|false|false|false|||ISSUES
Finding|Functional Concept|Hospital Course|9328,9335|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|Failure
Finding|Idea or Concept|Hospital Course|9328,9335|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|Failure
Finding|Individual Behavior|Hospital Course|9328,9335|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|Failure
Finding|Finding|Hospital Course|9341,9366|false|false|false|C4022792|Reduced left ventricular ejection fraction|reduced ejection fraction
Attribute|Clinical Attribute|Hospital Course|9349,9357|false|false|false|C0812388|Ejection time|ejection
Finding|Daily or Recreational Activity|Hospital Course|9349,9357|false|false|false|C0336969|Ejection as a Sports activity|ejection
Phenomenon|Phenomenon or Process|Hospital Course|9349,9357|false|false|false|C0302131|Ejection as a Circumstance of Injury|ejection
Finding|Finding|Hospital Course|9349,9366|false|false|false|C2020641;C2700378|Ejection fraction;stress echo measurements ejection fraction|ejection fraction
Procedure|Diagnostic Procedure|Hospital Course|9349,9366|false|false|false|C0489482|Ejection fraction (procedure)|ejection fraction
Event|Event|Hospital Course|9358,9366|false|false|false|||fraction
Finding|Intellectual Product|Hospital Course|9358,9366|false|false|false|C1554103|MDFAttributeType - Fraction|fraction
Finding|Functional Concept|Hospital Course|9369,9374|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Finding|Pathologic Function|Hospital Course|9369,9398|false|false|false|C0242707|Right Ventricular Dysfunction|Right ventricular dysfunction
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9375,9386|false|false|false|C0018827|Heart Ventricle|ventricular
Finding|Pathologic Function|Hospital Course|9375,9398|false|false|false|C0242973|Ventricular Dysfunction|ventricular dysfunction
Disorder|Disease or Syndrome|Hospital Course|9387,9398|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Event|Event|Hospital Course|9387,9398|false|false|false|||dysfunction
Finding|Conceptual Entity|Hospital Course|9387,9398|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|Hospital Course|9387,9398|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|Hospital Course|9387,9398|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Procedure|Health Care Activity|Hospital Course|9404,9408|false|false|false|C1315068|Pulmonary ventilator management|pulm
Disorder|Disease or Syndrome|Hospital Course|9409,9412|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|Hospital Course|9409,9412|false|false|false|||HTN
Finding|Intellectual Product|Hospital Course|9415,9421|false|false|false|C1705102|Volume (publication)|Volume
Finding|Pathologic Function|Hospital Course|9415,9430|false|false|false|C0546817|Hypervolemia (finding)|Volume overload
Event|Event|Hospital Course|9422,9430|false|false|false|||overload
Finding|Functional Concept|Hospital Course|9439,9446|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|Hospital Course|9439,9446|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|Hospital Course|9439,9446|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|Hospital Course|9447,9459|false|false|false|||exacerbation
Finding|Finding|Hospital Course|9447,9459|false|false|false|C4086268|Exacerbation|exacerbation
Finding|Finding|Hospital Course|9463,9469|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|9463,9469|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Disorder|Neoplastic Process|Hospital Course|9470,9479|false|false|false|C0027627|Neoplasm Metastasis|secondary
Event|Event|Hospital Course|9470,9479|false|false|false|||secondary
Finding|Functional Concept|Hospital Course|9470,9479|false|false|false|C1522484|metastatic qualifier|secondary
Event|Event|Hospital Course|9494,9508|false|false|false|||administration
Event|Occupational Activity|Hospital Course|9494,9508|false|false|false|C0001554|Administration occupational activities|administration
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9494,9508|false|false|false|C1533734|Administration (procedure)|administration
Drug|Substance|Hospital Course|9515,9521|false|false|false|C0302908|Liquid substance|fluids
Event|Event|Hospital Course|9515,9521|false|false|false|||fluids
Finding|Body Substance|Hospital Course|9515,9521|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9515,9521|false|false|false|C0016286|Fluid Therapy|fluids
Finding|Functional Concept|Hospital Course|9522,9536|false|false|false|C0332287|In addition to|in addition to
Event|Event|Hospital Course|9525,9533|false|false|false|||addition
Finding|Functional Concept|Hospital Course|9525,9533|false|false|false|C0332287;C1883712|Add - instruction imperative;In addition to|addition
Event|Event|Hospital Course|9541,9545|false|false|false|||self
Finding|Idea or Concept|Hospital Course|9541,9545|false|false|false|C0036588;C1551994|Self;subscriber - self|self
Finding|Intellectual Product|Hospital Course|9541,9545|false|false|false|C0036588;C1551994|Self;subscriber - self|self
Event|Event|Hospital Course|9551,9560|false|false|false|||titration
Procedure|Laboratory Procedure|Hospital Course|9551,9560|false|false|false|C0162621|Titration Method|titration
Drug|Organic Chemical|Hospital Course|9568,9577|false|false|false|C0076840|torsemide|torsemide
Drug|Pharmacologic Substance|Hospital Course|9568,9577|false|false|false|C0076840|torsemide|torsemide
Event|Event|Hospital Course|9568,9577|false|false|false|||torsemide
Finding|Intellectual Product|Hospital Course|9592,9596|false|false|false|C1561540|Transaction counts and value totals - week|week
Finding|Functional Concept|Hospital Course|9601,9609|false|false|false|C0332287;C1883712|Add - instruction imperative;In addition to|addition
Event|Event|Hospital Course|9623,9629|true|false|false|||follow
Finding|Functional Concept|Hospital Course|9632,9642|true|false|false|C0443288;C1548390;C1549594;C1610594|Confidentiality - restricted;Confidentiality code - Restricted;Document Confidentiality Status - Restricted;Restricted|restricted
Finding|Idea or Concept|Hospital Course|9632,9642|true|false|false|C0443288;C1548390;C1549594;C1610594|Confidentiality - restricted;Confidentiality code - Restricted;Document Confidentiality Status - Restricted;Restricted|restricted
Finding|Intellectual Product|Hospital Course|9632,9642|true|false|false|C0443288;C1548390;C1549594;C1610594|Confidentiality - restricted;Confidentiality code - Restricted;Document Confidentiality Status - Restricted;Restricted|restricted
Drug|Substance|Hospital Course|9643,9648|true|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|9643,9648|true|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|Hospital Course|9649,9655|true|false|false|||intake
Finding|Functional Concept|Hospital Course|9649,9655|true|false|false|C1512806|Intake|intake
Procedure|Health Care Activity|Hospital Course|9649,9655|true|false|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|intake
Event|Event|Hospital Course|9660,9666|true|false|false|||drinks
Event|Event|Hospital Course|9671,9678|false|false|false|||glasses
Drug|Inorganic Chemical|Hospital Course|9682,9687|false|false|false|C0043047;C1550678|Water Specimen;water|water
Drug|Pharmacologic Substance|Hospital Course|9682,9687|false|false|false|C0043047;C1550678|Water Specimen;water|water
Event|Event|Hospital Course|9682,9687|false|false|false|||water
Finding|Intellectual Product|Hospital Course|9682,9687|false|false|false|C1547961|Water - Specimen Source Codes|water
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9682,9687|false|false|false|C0020311|Hydrotherapy|water
Drug|Food|Hospital Course|9691,9696|false|false|false|C1268568|Juice|juice
Event|Event|Hospital Course|9691,9696|false|false|false|||juice
Event|Event|Hospital Course|9728,9737|true|false|false|||tolerated
Event|Event|Hospital Course|9738,9747|true|false|false|||guideline
Finding|Intellectual Product|Hospital Course|9738,9747|true|false|false|C0162791;C0282423|Guideline (Publication Type);Guidelines|guideline
Event|Event|Hospital Course|9748,9756|true|false|false|||directed
Finding|Functional Concept|Hospital Course|9757,9764|true|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|Hospital Course|9757,9764|true|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|Hospital Course|9757,9764|true|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|Hospital Course|9757,9764|true|false|false|C0199168|Medical service|medical
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9757,9772|true|false|false|C0418981;C2069680|Medical therapy;disposition medical therapy|medical therapy
Event|Event|Hospital Course|9765,9772|true|false|false|||therapy
Finding|Finding|Hospital Course|9765,9772|true|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|Hospital Course|9765,9772|true|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9765,9772|true|false|false|C0087111|Therapeutic procedure|therapy
Event|Event|Hospital Course|9790,9796|false|false|false|||issues
Finding|Intellectual Product|Hospital Course|9802,9807|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Disease or Syndrome|Hospital Course|9802,9821|false|false|false|C0022660;C2609414|Acute kidney injury;Kidney Failure, Acute|acute kidney injury
Disorder|Injury or Poisoning|Hospital Course|9802,9821|false|false|false|C0022660;C2609414|Acute kidney injury;Kidney Failure, Acute|acute kidney injury
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9808,9814|false|false|false|C0022646;C0227665|Both kidneys;Kidney|kidney
Disorder|Neoplastic Process|Hospital Course|9808,9814|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|kidney
Event|Event|Hospital Course|9808,9814|false|false|false|||kidney
Finding|Sign or Symptom|Hospital Course|9808,9814|false|false|false|C0812426|Kidney problem|kidney
Procedure|Diagnostic Procedure|Hospital Course|9808,9814|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9808,9814|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Disorder|Injury or Poisoning|Hospital Course|9808,9821|false|false|false|C0160420|Injury of kidney|kidney injury
Disorder|Injury or Poisoning|Hospital Course|9815,9821|false|false|false|C3263722;C3263723|Traumatic AND/OR non-traumatic injury;Traumatic injury|injury
Event|Event|Hospital Course|9815,9821|false|false|false|||injury
Event|Event|Hospital Course|9835,9848|false|false|false|||transaminitis
Finding|Finding|Hospital Course|9835,9848|false|false|false|C2242708|Hypertransaminasaemia|transaminitis
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9858,9871|false|false|false|C3658706|pembrolizumab|pembrolizumab
Drug|Immunologic Factor|Hospital Course|9858,9871|false|false|false|C3658706|pembrolizumab|pembrolizumab
Drug|Pharmacologic Substance|Hospital Course|9858,9871|false|false|false|C3658706|pembrolizumab|pembrolizumab
Event|Event|Hospital Course|9872,9879|false|false|false|||therapy
Finding|Finding|Hospital Course|9872,9879|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|Hospital Course|9872,9879|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9872,9879|false|false|false|C0087111|Therapeutic procedure|therapy
Event|Event|Hospital Course|9899,9905|false|false|false|||volume
Finding|Intellectual Product|Hospital Course|9899,9905|false|false|false|C1705102|Volume (publication)|volume
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9931,9934|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Hormone|Hospital Course|9931,9934|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Pharmacologic Substance|Hospital Course|9931,9934|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Event|Event|Hospital Course|9931,9934|false|false|false|||BNP
Finding|Gene or Genome|Hospital Course|9931,9934|false|false|false|C1417808;C2982014|NPPB gene;NPPB wt Allele|BNP
Procedure|Laboratory Procedure|Hospital Course|9931,9934|false|false|false|C1095989|Brain natriuretic peptide measurement|BNP
Event|Event|Hospital Course|9945,9954|false|false|false|||initiated
Drug|Organic Chemical|Hospital Course|9958,9963|false|false|false|C0699992|Lasix|lasix
Drug|Pharmacologic Substance|Hospital Course|9958,9963|false|false|false|C0699992|Lasix|lasix
Event|Event|Hospital Course|9958,9963|false|false|false|||lasix
Event|Event|Hospital Course|9968,9973|false|false|false|||bolus
Finding|Body Substance|Hospital Course|9968,9973|false|false|false|C1186706;C1550436|Bolus of ingested food;Response Modality - Bolus|bolus
Finding|Intellectual Product|Hospital Course|9968,9973|false|false|false|C1186706;C1550436|Bolus of ingested food;Response Modality - Bolus|bolus
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9968,9973|false|false|false|C1511237|bolus infusion|bolus
Drug|Organic Chemical|Hospital Course|9992,9997|false|false|false|C0699992|Lasix|lasix
Drug|Pharmacologic Substance|Hospital Course|9992,9997|false|false|false|C0699992|Lasix|lasix
Disorder|Neoplastic Process|Hospital Course|9998,10001|false|false|false|C1135868|Gestational Trophoblastic Neoplasms|gtt
Drug|Biomedical or Dental Material|Hospital Course|9998,10001|false|false|false|C0991568|Drops - Drug Form|gtt
Event|Event|Hospital Course|9998,10001|false|false|false|||gtt
Procedure|Laboratory Procedure|Hospital Course|9998,10001|false|false|false|C0017741|Glucose tolerance test|gtt
Finding|Idea or Concept|Hospital Course|10007,10011|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Finding|Finding|Hospital Course|10007,10020|false|false|false|C5453003|Good response|good response
Event|Event|Hospital Course|10012,10020|false|false|false|||response
Finding|Finding|Hospital Course|10012,10020|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Intellectual Product|Hospital Course|10012,10020|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Mental Process|Hospital Course|10012,10020|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Event|Event|Hospital Course|10040,10049|false|false|false|||increased
Event|Event|Hospital Course|10075,10083|false|false|false|||improved
Disorder|Cell or Molecular Dysfunction|Hospital Course|10089,10099|false|false|false|C0599156|Transition Mutation|transition
Event|Activity|Hospital Course|10089,10099|false|false|false|C2700061|Transition (action)|transition
Event|Event|Hospital Course|10089,10099|false|false|false|||transition
Drug|Organic Chemical|Hospital Course|10106,10115|false|false|false|C0076840|torsemide|Torsemide
Drug|Pharmacologic Substance|Hospital Course|10106,10115|false|false|false|C0076840|torsemide|Torsemide
Event|Event|Hospital Course|10106,10115|false|false|false|||Torsemide
Event|Event|Hospital Course|10133,10142|false|false|false|||monitored
Event|Event|Hospital Course|10160,10168|false|false|false|||repleted
Drug|Biologically Active Substance|Hospital Course|10174,10183|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Element, Ion, or Isotope|Hospital Course|10174,10183|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Food|Hospital Course|10174,10183|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Inorganic Chemical|Hospital Course|10174,10183|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Pharmacologic Substance|Hospital Course|10174,10183|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Event|Event|Hospital Course|10174,10183|false|false|false|||potassium
Finding|Physiologic Function|Hospital Course|10174,10183|false|false|false|C4553027|Potassium metabolic function|potassium
Procedure|Laboratory Procedure|Hospital Course|10174,10183|false|false|false|C0202194|Potassium measurement|potassium
Event|Event|Hospital Course|10198,10207|true|false|false|||reduction
Finding|Finding|Hospital Course|10198,10207|true|false|false|C0392756|Reduced|reduction
Phenomenon|Natural Phenomenon or Process|Hospital Course|10198,10207|true|false|false|C0301630|Reduction (chemical)|reduction
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10198,10207|true|false|false|C1293152;C4551656|Reduction procedure;Surgical reduction|reduction
Event|Event|Hospital Course|10211,10217|true|false|false|||neural
Finding|Functional Concept|Hospital Course|10211,10217|true|false|false|C3714606|Neural|neural
Drug|Element, Ion, or Isotope|Hospital Course|10227,10235|true|false|false|C3540676|Blockade|blockade
Drug|Pharmacologic Substance|Hospital Course|10227,10235|true|false|false|C3540676|Blockade|blockade
Event|Event|Hospital Course|10227,10235|true|false|false|||blockade
Finding|Functional Concept|Hospital Course|10227,10235|true|false|false|C0332206|Blocking|blockade
Event|Event|Hospital Course|10241,10246|false|false|false|||added
Finding|Intellectual Product|Hospital Course|10251,10258|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|Hospital Course|10251,10258|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Disorder|Disease or Syndrome|Hospital Course|10251,10273|false|false|false|C1561643|Chronic Kidney Diseases|Chronic Kidney Disease
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10259,10265|false|false|false|C0022646;C0227665|Both kidneys;Kidney|Kidney
Disorder|Neoplastic Process|Hospital Course|10259,10265|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|Kidney
Event|Event|Hospital Course|10259,10265|false|false|false|||Kidney
Finding|Sign or Symptom|Hospital Course|10259,10265|false|false|false|C0812426|Kidney problem|Kidney
Procedure|Diagnostic Procedure|Hospital Course|10259,10265|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|Kidney
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10259,10265|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|Kidney
Disorder|Disease or Syndrome|Hospital Course|10259,10273|false|false|false|C0022658|Kidney Diseases|Kidney Disease
Disorder|Disease or Syndrome|Hospital Course|10266,10273|false|false|false|C0012634|Disease|Disease
Drug|Biomedical or Dental Material|Hospital Course|10275,10283|false|false|false|C0168634|BaseLine dental cement|Baseline
Event|Event|Hospital Course|10275,10283|false|false|false|||Baseline
Finding|Idea or Concept|Hospital Course|10275,10283|false|false|false|C1552824|baseline - TableCellVerticalAlign|Baseline
Event|Event|Hospital Course|10305,10314|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|10305,10314|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|Hospital Course|10315,10321|false|false|false|||Stable
Finding|Intellectual Product|Hospital Course|10315,10321|false|false|false|C1547311|Patient Condition Code - Stable|Stable
Event|Event|Hospital Course|10331,10340|false|false|false|||discharge
Finding|Body Substance|Hospital Course|10331,10340|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|10331,10340|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|10331,10340|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|10331,10340|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|Hospital Course|10358,10367|false|false|false|||uptrended
Drug|Biomedical or Dental Material|Hospital Course|10374,10382|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|Hospital Course|10374,10382|false|false|false|||baseline
Finding|Idea or Concept|Hospital Course|10374,10382|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Finding|Hospital Course|10407,10413|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|10407,10413|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Drug|Pharmacologic Substance|Hospital Course|10431,10439|false|false|false|C0012798;C5399719|Diuretic [APC];Diuretics|diuretic
Finding|Finding|Hospital Course|10431,10445|false|false|false|C0239192|DIURETIC USAGE|diuretic usage
Event|Event|Hospital Course|10440,10445|false|false|false|||usage
Finding|Functional Concept|Hospital Course|10440,10445|false|false|false|C0457083|Usage|usage
Event|Event|Hospital Course|10452,10460|false|false|false|||improved
Drug|Pharmacologic Substance|Hospital Course|10476,10485|false|false|false|C0012798|Diuretics|diuretics
Event|Event|Hospital Course|10476,10485|false|false|false|||diuretics
Finding|Finding|Hospital Course|10492,10498|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|10492,10498|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Disorder|Disease or Syndrome|Hospital Course|10499,10519|false|true|false|C2242703|Cardio-Renal Syndrome|cardiorenal syndrome
Disorder|Disease or Syndrome|Hospital Course|10511,10519|false|true|false|C0039082|Syndrome|syndrome
Event|Event|Hospital Course|10511,10519|false|false|false|||syndrome
Event|Event|Hospital Course|10525,10533|false|false|false|||addition
Finding|Functional Concept|Hospital Course|10525,10533|false|false|false|C0332287;C1883712|Add - instruction imperative;In addition to|addition
Event|Event|Hospital Course|10534,10541|false|false|false|||patient
Finding|Body Substance|Hospital Course|10534,10541|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|10534,10541|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|10534,10541|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|10555,10559|false|false|false|||seen
Finding|Functional Concept|Hospital Course|10563,10569|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|Hospital Course|10563,10569|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|Hospital Course|10563,10572|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|Hospital Course|10563,10572|false|false|false|C1522577|follow-up|follow-up
Event|Event|Hospital Course|10594,10598|false|false|false|||felt
Disorder|Disease or Syndrome|Hospital Course|10603,10606|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Event|Event|Hospital Course|10603,10606|false|false|false|||CKD
Event|Event|Hospital Course|10616,10622|false|false|false|||likely
Finding|Finding|Hospital Course|10616,10622|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|10616,10622|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Drug|Organic Chemical|Hospital Course|10629,10636|false|true|false|C0163712|Relate - vinyl resin|related
Event|Event|Hospital Course|10629,10636|false|false|false|||related
Finding|Finding|Hospital Course|10629,10636|false|true|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|Hospital Course|10629,10636|false|true|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10640,10653|false|true|false|C3658706|pembrolizumab|pembrolizumab
Drug|Immunologic Factor|Hospital Course|10640,10653|false|true|false|C3658706|pembrolizumab|pembrolizumab
Drug|Pharmacologic Substance|Hospital Course|10640,10653|false|true|false|C3658706|pembrolizumab|pembrolizumab
Event|Event|Hospital Course|10640,10653|false|false|false|||pembrolizumab
Finding|Finding|Hospital Course|10664,10670|true|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|10664,10670|true|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Drug|Organic Chemical|Hospital Course|10671,10678|true|true|false|C0163712|Relate - vinyl resin|related
Event|Event|Hospital Course|10671,10678|true|false|false|||related
Finding|Finding|Hospital Course|10671,10678|true|true|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|Hospital Course|10671,10678|true|true|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Attribute|Clinical Attribute|Hospital Course|10682,10685|true|true|false|C1114365||age
Drug|Biologically Active Substance|Hospital Course|10682,10685|true|true|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|Hospital Course|10682,10685|true|true|false|C0162574|Glycation End Products, Advanced|age
Event|Event|Hospital Course|10682,10685|true|false|false|||age
Drug|Organic Chemical|Hospital Course|10686,10693|true|true|false|C0163712|Relate - vinyl resin|related
Event|Event|Hospital Course|10686,10693|true|false|false|||related
Finding|Finding|Hospital Course|10686,10693|true|true|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|Hospital Course|10686,10693|true|true|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Event|Event|Hospital Course|10694,10701|false|false|false|||decline
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10705,10710|true|false|false|C0022646|Kidney|renal
Disorder|Disease or Syndrome|Hospital Course|10705,10710|true|false|false|C0042075|Urologic Diseases|renal
Event|Event|Hospital Course|10712,10720|true|false|false|||function
Finding|Finding|Hospital Course|10712,10720|true|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|Hospital Course|10712,10720|true|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|Hospital Course|10712,10720|true|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|Hospital Course|10712,10720|true|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Drug|Biologically Active Substance|Hospital Course|10722,10732|false|false|false|C0010294|creatinine|Creatinine
Drug|Organic Chemical|Hospital Course|10722,10732|false|false|false|C0010294|creatinine|Creatinine
Event|Event|Hospital Course|10722,10732|false|false|false|||Creatinine
Finding|Physiologic Function|Hospital Course|10722,10732|false|false|false|C4551889|Creatinine metabolic function|Creatinine
Procedure|Laboratory Procedure|Hospital Course|10722,10732|false|false|false|C0201975|Creatinine measurement|Creatinine
Event|Event|Hospital Course|10740,10749|false|false|false|||discharge
Finding|Body Substance|Hospital Course|10740,10749|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|10740,10749|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|10740,10749|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|10740,10749|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|Hospital Course|10751,10757|false|false|false|||stable
Finding|Intellectual Product|Hospital Course|10751,10757|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Functional Concept|Hospital Course|10763,10773|false|false|false|C0036525;C1522484|Metastatic to;metastatic qualifier|Metastatic
Disorder|Neoplastic Process|Hospital Course|10763,10782|false|false|false|C0278883|Metastatic melanoma|Metastatic Melanoma
Disorder|Neoplastic Process|Hospital Course|10774,10782|false|false|false|C0025202|melanoma|Melanoma
Drug|Immunologic Factor|Hospital Course|10774,10782|false|false|false|C0796561|Melanoma vaccine|Melanoma
Drug|Pharmacologic Substance|Hospital Course|10774,10782|false|false|false|C0796561|Melanoma vaccine|Melanoma
Event|Event|Hospital Course|10774,10782|false|false|false|||Melanoma
Event|Event|Hospital Course|10790,10798|false|false|false|||followed
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10832,10845|false|false|false|C3658706|pembrolizumab|Pembrolizumab
Drug|Immunologic Factor|Hospital Course|10832,10845|false|false|false|C3658706|pembrolizumab|Pembrolizumab
Drug|Pharmacologic Substance|Hospital Course|10832,10845|false|false|false|C3658706|pembrolizumab|Pembrolizumab
Event|Event|Hospital Course|10856,10860|false|false|false|||held
Event|Event|Hospital Course|10865,10873|false|false|false|||diarrhea
Finding|Finding|Hospital Course|10865,10873|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|Hospital Course|10865,10873|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Event|Event|Hospital Course|10884,10888|false|false|false|||LFTs
Event|Event|Hospital Course|10893,10902|false|false|false|||worsening
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10903,10909|false|false|false|C0022646;C0227665|Both kidneys;Kidney|kidney
Disorder|Neoplastic Process|Hospital Course|10903,10909|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|kidney
Event|Event|Hospital Course|10903,10909|false|false|false|||kidney
Finding|Sign or Symptom|Hospital Course|10903,10909|false|false|false|C0812426|Kidney problem|kidney
Procedure|Diagnostic Procedure|Hospital Course|10903,10909|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10903,10909|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Finding|Organ or Tissue Function|Hospital Course|10903,10918|false|false|false|C0232804|Renal function|kidney function
Event|Event|Hospital Course|10910,10918|false|false|false|||function
Finding|Finding|Hospital Course|10910,10918|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|Hospital Course|10910,10918|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|Hospital Course|10910,10918|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|Hospital Course|10910,10918|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Classification|Hospital Course|10920,10928|true|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Finding|Finding|Hospital Course|10920,10928|true|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Lab|Laboratory or Test Result|Hospital Course|10920,10928|true|false|false|C5237010|Expression Negative|Negative
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10929,10937|true|false|false|C0041199|Troponin|troponin
Drug|Biologically Active Substance|Hospital Course|10929,10937|true|false|false|C0041199|Troponin|troponin
Event|Event|Hospital Course|10929,10937|true|false|false|||troponin
Procedure|Laboratory Procedure|Hospital Course|10929,10937|true|false|false|C0523952|Troponin measurement|troponin
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10942,10947|true|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK MB
Drug|Enzyme|Hospital Course|10942,10947|true|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK MB
Procedure|Laboratory Procedure|Hospital Course|10942,10947|true|false|false|C0523584|Creatine kinase MB measurement|CK MB
Event|Event|Hospital Course|10945,10947|true|false|false|||MB
Event|Event|Hospital Course|10953,10960|true|false|false|||concern
Finding|Idea or Concept|Hospital Course|10953,10960|true|false|false|C2699424|Concern|concern
Drug|Pharmacologic Substance|Hospital Course|10965,10969|true|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|drug
Finding|Finding|Hospital Course|10965,10969|true|false|false|C0740721|Drug problem|drug
Disorder|Disease or Syndrome|Hospital Course|10978,10989|false|false|false|C0027059|Myocarditis|myocarditis
Event|Event|Hospital Course|10978,10989|false|false|false|||myocarditis
Event|Event|Hospital Course|11005,11013|false|false|false|||Followup
Procedure|Health Care Activity|Hospital Course|11005,11013|false|false|false|C1522577|follow-up|Followup
Event|Event|Hospital Course|11045,11054|false|false|false|||discharge
Finding|Body Substance|Hospital Course|11045,11054|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|11045,11054|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|11045,11054|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|11045,11054|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|Hospital Course|11067,11081|false|false|false|||transaminiatis
Event|Event|Hospital Course|11082,11088|false|false|false|||Stable
Finding|Intellectual Product|Hospital Course|11082,11088|false|false|false|C1547311|Patient Condition Code - Stable|Stable
Drug|Organic Chemical|Hospital Course|11090,11096|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Statin
Drug|Pharmacologic Substance|Hospital Course|11090,11096|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Statin
Event|Event|Hospital Course|11090,11096|false|false|false|||Statin
Finding|Gene or Genome|Hospital Course|11090,11096|false|false|false|C1414273|EEF1A2 gene|Statin
Event|Event|Hospital Course|11125,11129|false|false|false|||held
Event|Event|Hospital Course|11134,11141|true|false|false|||changes
Finding|Functional Concept|Hospital Course|11134,11141|true|false|false|C0392747|Changing|changes
Event|Event|Hospital Course|11142,11146|true|false|false|||made
Event|Event|Hospital Course|11155,11164|true|false|false|||admission
Procedure|Health Care Activity|Hospital Course|11155,11164|true|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11170,11177|false|false|false|C0042027|Urinary tract|Urinary
Finding|Finding|Hospital Course|11170,11187|false|false|false|C0042023|Increased frequency of micturition|Urinary frequency
Event|Event|Hospital Course|11178,11187|false|false|false|||frequency
Finding|Intellectual Product|Hospital Course|11178,11187|false|false|false|C3898838;C4321352|Frequency;How Often|frequency
Event|Event|Hospital Course|11188,11194|false|false|false|||Likely
Finding|Finding|Hospital Course|11188,11194|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Idea or Concept|Hospital Course|11188,11194|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Drug|Pharmacologic Substance|Hospital Course|11202,11210|false|true|false|C0012798;C5399719|Diuretic [APC];Diuretics|diuretic
Event|Event|Hospital Course|11211,11214|false|false|false|||use
Finding|Functional Concept|Hospital Course|11211,11214|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|Hospital Course|11211,11214|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Event|Event|Hospital Course|11216,11224|false|false|false|||Afebrile
Finding|Finding|Hospital Course|11216,11224|false|false|false|C0277797|Apyrexial|Afebrile
Finding|Idea or Concept|Hospital Course|11254,11258|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|11254,11258|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|11254,11258|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|11259,11269|false|false|false|C0257343|tamsulosin|tamsulosin
Drug|Pharmacologic Substance|Hospital Course|11259,11269|false|false|false|C0257343|tamsulosin|tamsulosin
Event|Event|Hospital Course|11259,11269|false|false|false|||tamsulosin
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11273,11281|false|false|false|C0018787|Heart|Coronary
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11273,11288|false|false|false|C0205042|Coronary artery|Coronary artery
Disorder|Disease or Syndrome|Hospital Course|11273,11296|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|Coronary artery disease
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11282,11288|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|Hospital Course|11282,11288|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Disorder|Disease or Syndrome|Hospital Course|11282,11296|false|false|false|C0852949|Arteriopathic disease|artery disease
Disorder|Disease or Syndrome|Hospital Course|11289,11296|false|false|false|C0012634|Disease|disease
Event|Event|Hospital Course|11289,11296|false|false|false|||disease
Event|Event|Hospital Course|11302,11306|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11302,11306|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11311,11314|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|Hospital Course|11311,11314|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|Hospital Course|11311,11314|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11315,11318|false|false|false|C2713669|SERPINA5 protein, human|PCI
Drug|Biologically Active Substance|Hospital Course|11315,11318|false|false|false|C2713669|SERPINA5 protein, human|PCI
Event|Event|Hospital Course|11315,11318|false|false|false|||PCI
Finding|Gene or Genome|Hospital Course|11315,11318|false|false|false|C1418370;C1705930;C4049621|Peritoneal Cancer Index;SERPINA5 gene;SERPINA5 wt Allele|PCI
Finding|Intellectual Product|Hospital Course|11315,11318|false|false|false|C1418370;C1705930;C4049621|Peritoneal Cancer Index;SERPINA5 gene;SERPINA5 wt Allele|PCI
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11315,11318|false|false|false|C1514496;C1532338;C4724254|Percutaneous Coronary Intervention;Prophylactic Cranial Irradiation;photochemical internalization|PCI
Event|Event|Hospital Course|11321,11330|false|false|false|||Continued
Drug|Organic Chemical|Hospital Course|11331,11338|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|Hospital Course|11331,11338|false|false|false|C0004057|aspirin|aspirin
Event|Event|Hospital Course|11331,11338|false|false|false|||aspirin
Drug|Organic Chemical|Hospital Course|11352,11358|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Statin
Drug|Pharmacologic Substance|Hospital Course|11352,11358|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Statin
Event|Event|Hospital Course|11352,11358|false|false|false|||Statin
Finding|Gene or Genome|Hospital Course|11352,11358|false|false|false|C1414273|EEF1A2 gene|Statin
Event|Event|Hospital Course|11359,11366|false|false|false|||stopped
Event|Event|Hospital Course|11376,11385|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|11376,11385|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|Hospital Course|11402,11406|false|false|false|||LFTs
Event|Event|Hospital Course|11419,11426|false|false|false|||holding
Event|Event|Hospital Course|11430,11437|false|false|false|||CHRONIC
Finding|Intellectual Product|Hospital Course|11430,11437|false|false|false|C1547296|Chronic - Admission Level of Care Code|CHRONIC
Procedure|Health Care Activity|Hospital Course|11430,11437|false|false|false|C1555457|Provision of recurring care for chronic illness|CHRONIC
Disorder|Disease or Syndrome|Hospital Course|11466,11496|false|false|false|C0235480|Paroxysmal atrial fibrillation|Paroxysmal Atrial fibrillation
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11477,11483|false|false|false|C0018792|Heart Atrium|Atrial
Attribute|Clinical Attribute|Hospital Course|11477,11496|false|false|false|C2926591||Atrial fibrillation
Disorder|Disease or Syndrome|Hospital Course|11477,11496|false|false|false|C0004238|Atrial Fibrillation|Atrial fibrillation
Lab|Laboratory or Test Result|Hospital Course|11477,11496|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Atrial fibrillation
Disorder|Disease or Syndrome|Hospital Course|11484,11496|false|false|false|C0232197|Fibrillation|fibrillation
Event|Event|Hospital Course|11484,11496|false|false|false|||fibrillation
Event|Event|Hospital Course|11505,11513|false|false|false|||Continue
Drug|Organic Chemical|Hospital Course|11514,11524|false|false|false|C0002598|amiodarone|amiodarone
Drug|Pharmacologic Substance|Hospital Course|11514,11524|false|false|false|C0002598|amiodarone|amiodarone
Event|Event|Hospital Course|11514,11524|false|false|false|||amiodarone
Procedure|Laboratory Procedure|Hospital Course|11514,11524|false|false|false|C5399868|Drug assay amiodarone|amiodarone
Event|Event|Hospital Course|11525,11530|false|false|false|||200mg
Finding|Finding|Hospital Course|11535,11541|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|Hospital Course|11535,11541|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Drug|Organic Chemical|Hospital Course|11542,11549|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|Hospital Course|11542,11549|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|Hospital Course|11542,11549|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Event|Event|Hospital Course|11542,11549|false|false|false|||control
Finding|Conceptual Entity|Hospital Course|11542,11549|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|Hospital Course|11542,11549|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|Hospital Course|11542,11549|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Event|Event|Hospital Course|11550,11558|false|false|false|||strategy
Finding|Mental Process|Hospital Course|11550,11558|false|false|false|C0679199|Strategy|strategy
Event|Activity|Hospital Course|11560,11570|false|false|false|C1283169||monitoring
Procedure|Health Care Activity|Hospital Course|11560,11570|false|false|false|C0150369|Preventive monitoring|monitoring
Phenomenon|Human-caused Phenomenon or Process|Hospital Course|11571,11577|false|false|false|C0036043|Safety|safety
Lab|Laboratory or Test Result|Hospital Course|11578,11582|false|false|false|C0587081|Laboratory test finding|labs
Event|Event|Hospital Course|11595,11610|false|false|false|||anticoagulation
Finding|Finding|Hospital Course|11595,11610|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|Hospital Course|11595,11610|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11595,11610|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Drug|Organic Chemical|Hospital Course|11616,11624|false|false|false|C1831808|apixaban|apixaban
Drug|Pharmacologic Substance|Hospital Course|11616,11624|false|false|false|C1831808|apixaban|apixaban
Event|Event|Hospital Course|11616,11624|false|false|false|||apixaban
Disorder|Disease or Syndrome|Hospital Course|11646,11658|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|Hospital Course|11646,11658|false|false|false|||Hypertension
Event|Event|Hospital Course|11660,11666|false|false|false|||Stable
Finding|Intellectual Product|Hospital Course|11660,11666|false|false|false|C1547311|Patient Condition Code - Stable|Stable
Attribute|Clinical Attribute|Hospital Course|11671,11682|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|11671,11682|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|11671,11682|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|11671,11682|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|11671,11695|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|11686,11695|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|11686,11695|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|Hospital Course|11714,11724|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Hospital Course|11714,11724|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|Hospital Course|11714,11729|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|Hospital Course|11725,11729|false|false|false|||list
Finding|Intellectual Product|Hospital Course|11725,11729|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|Hospital Course|11737,11747|false|false|false|||inaccurate
Event|Event|Hospital Course|11752,11760|false|false|false|||requires
Event|Event|Hospital Course|11770,11783|false|false|false|||investigation
Finding|Intellectual Product|Hospital Course|11770,11783|false|false|false|C1552578|Act Class - investigation|investigation
Procedure|Health Care Activity|Hospital Course|11770,11783|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|investigation
Drug|Organic Chemical|Hospital Course|11788,11798|false|false|false|C0002598|amiodarone|Amiodarone
Drug|Pharmacologic Substance|Hospital Course|11788,11798|false|false|false|C0002598|amiodarone|Amiodarone
Event|Event|Hospital Course|11788,11798|false|false|false|||Amiodarone
Procedure|Laboratory Procedure|Hospital Course|11788,11798|false|false|false|C5399868|Drug assay amiodarone|Amiodarone
Drug|Organic Chemical|Hospital Course|11819,11826|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Hospital Course|11819,11826|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|Hospital Course|11846,11854|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|11846,11854|false|false|false|C1692318|docusate|Docusate
Event|Event|Hospital Course|11846,11854|false|false|false|||Docusate
Drug|Organic Chemical|Hospital Course|11846,11861|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|Hospital Course|11846,11861|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|Hospital Course|11855,11861|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|11855,11861|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|11855,11861|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|11855,11861|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|11855,11861|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|11855,11861|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|Hospital Course|11872,11875|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11872,11875|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|11872,11875|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|11872,11875|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|11872,11875|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|11880,11885|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|Hospital Course|11880,11885|false|false|false|C3489575|sennosides, USP|Senna
Drug|Organic Chemical|Hospital Course|11904,11911|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|11904,11911|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|11904,11911|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|Hospital Course|11904,11913|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|Hospital Course|11904,11913|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|Hospital Course|11904,11913|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|Hospital Course|11904,11913|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|Hospital Course|11904,11913|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|Hospital Course|11912,11913|false|false|false|||D
Event|Event|Hospital Course|11919,11923|false|false|false|||UNIT
Drug|Organic Chemical|Hospital Course|11937,11942|false|false|false|C2369992|Align|Align
Drug|Pharmacologic Substance|Hospital Course|11937,11942|false|false|false|C2369992|Align|Align
Drug|Pharmacologic Substance|Hospital Course|11944,11968|false|false|false|C4019097|herbal medicines bifidobacterium infantis|bifidobacterium infantis
Event|Event|Hospital Course|11960,11968|false|false|false|||infantis
Anatomy|Body Space or Junction|Hospital Course|11975,11979|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|11975,11979|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|11975,11979|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|11975,11979|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|Hospital Course|11980,11985|false|false|false|||DAILY
Drug|Biologically Active Substance|Hospital Course|11990,11998|false|false|false|C0009235|Coenzymes|coenzyme
Drug|Organic Chemical|Hospital Course|11990,11998|false|false|false|C0009235|Coenzymes|coenzyme
Event|Event|Hospital Course|11990,11998|false|false|false|||coenzyme
Drug|Biologically Active Substance|Hospital Course|11990,12002|false|false|false|C0041536|ubidecarenone|coenzyme Q10
Drug|Organic Chemical|Hospital Course|11990,12002|false|false|false|C0041536|ubidecarenone|coenzyme Q10
Drug|Pharmacologic Substance|Hospital Course|11990,12002|false|false|false|C0041536|ubidecarenone|coenzyme Q10
Event|Event|Hospital Course|11999,12002|false|false|false|||Q10
Finding|Gene or Genome|Hospital Course|11999,12002|false|false|false|C1414333;C2827473|AGO2 gene;AGO2 wt Allele|Q10
Anatomy|Body Space or Junction|Hospital Course|12010,12014|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|12010,12014|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|12010,12014|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|12010,12014|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|Hospital Course|12015,12020|false|false|false|||DAILY
Drug|Organic Chemical|Hospital Course|12025,12035|false|false|false|C0257343|tamsulosin|Tamsulosin
Drug|Pharmacologic Substance|Hospital Course|12025,12035|false|false|false|C0257343|tamsulosin|Tamsulosin
Event|Event|Hospital Course|12046,12049|false|false|false|||QHS
Drug|Organic Chemical|Hospital Course|12054,12063|false|false|false|C0076840|torsemide|Torsemide
Drug|Pharmacologic Substance|Hospital Course|12054,12063|false|false|false|C0076840|torsemide|Torsemide
Drug|Element, Ion, or Isotope|Hospital Course|12084,12091|false|false|false|C2346592|Ferrous|Ferrous
Drug|Inorganic Chemical|Hospital Course|12084,12099|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Pharmacologic Substance|Hospital Course|12084,12099|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Element, Ion, or Isotope|Hospital Course|12092,12099|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Inorganic Chemical|Hospital Course|12092,12099|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Pharmacologic Substance|Hospital Course|12092,12099|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Event|Event|Hospital Course|12092,12099|false|false|false|||Sulfate
Drug|Organic Chemical|Hospital Course|12121,12131|false|false|false|C0074393|sertraline|Sertraline
Drug|Pharmacologic Substance|Hospital Course|12121,12131|false|false|false|C0074393|sertraline|Sertraline
Drug|Biologically Active Substance|Hospital Course|12152,12161|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|Hospital Course|12152,12161|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|Hospital Course|12152,12161|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|Hospital Course|12152,12161|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|Hospital Course|12152,12161|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Event|Event|Hospital Course|12152,12161|false|false|false|||Potassium
Finding|Physiologic Function|Hospital Course|12152,12161|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|Hospital Course|12152,12161|false|false|false|C0202194|Potassium measurement|Potassium
Drug|Inorganic Chemical|Hospital Course|12152,12170|false|false|false|C0032825|potassium chloride|Potassium Chloride
Drug|Pharmacologic Substance|Hospital Course|12152,12170|false|false|false|C0032825|potassium chloride|Potassium Chloride
Drug|Element, Ion, or Isotope|Hospital Course|12162,12170|false|false|false|C0008203;C0596019|Chlorides;chloride ion|Chloride
Event|Event|Hospital Course|12162,12170|false|false|false|||Chloride
Finding|Physiologic Function|Hospital Course|12162,12170|false|false|false|C4553021|Chloride metabolic function|Chloride
Procedure|Laboratory Procedure|Hospital Course|12162,12170|false|false|false|C0201952|Chloride measurement|Chloride
Event|Event|Hospital Course|12174,12177|false|false|false|||mEq
Disorder|Mental or Behavioral Dysfunction|Hospital Course|12181,12184|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12181,12184|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|12181,12184|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|12181,12184|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|12181,12184|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|12190,12198|false|false|false|C1831808|apixaban|Apixaban
Drug|Pharmacologic Substance|Hospital Course|12190,12198|false|false|false|C1831808|apixaban|Apixaban
Disorder|Mental or Behavioral Dysfunction|Hospital Course|12209,12212|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12209,12212|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|12209,12212|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|12209,12212|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|12209,12212|false|false|false|C1332410|BID gene|BID
Drug|Antibiotic|Hospital Course|12218,12228|false|false|false|C0007716|cephalexin|Cephalexin
Drug|Organic Chemical|Hospital Course|12218,12228|false|false|false|C0007716|cephalexin|Cephalexin
Event|Event|Hospital Course|12247,12256|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|12247,12256|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|12247,12256|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|12247,12256|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|12247,12256|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|12247,12268|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|12257,12268|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|12257,12268|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|12257,12268|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|12257,12268|false|false|false|C4284232|Medications|Medications
Drug|Biologically Active Substance|Hospital Course|12274,12283|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|Hospital Course|12274,12283|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|Hospital Course|12274,12283|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|Hospital Course|12274,12283|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|Hospital Course|12274,12283|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Event|Event|Hospital Course|12274,12283|false|false|false|||Potassium
Finding|Physiologic Function|Hospital Course|12274,12283|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|Hospital Course|12274,12283|false|false|false|C0202194|Potassium measurement|Potassium
Drug|Inorganic Chemical|Hospital Course|12274,12292|false|false|false|C0032825|potassium chloride|Potassium Chloride
Drug|Pharmacologic Substance|Hospital Course|12274,12292|false|false|false|C0032825|potassium chloride|Potassium Chloride
Drug|Element, Ion, or Isotope|Hospital Course|12284,12292|false|false|false|C0008203;C0596019|Chlorides;chloride ion|Chloride
Event|Event|Hospital Course|12284,12292|false|false|false|||Chloride
Finding|Physiologic Function|Hospital Course|12284,12292|false|false|false|C4553021|Chloride metabolic function|Chloride
Procedure|Laboratory Procedure|Hospital Course|12284,12292|false|false|false|C0201952|Chloride measurement|Chloride
Event|Event|Hospital Course|12296,12299|false|false|false|||mEq
Drug|Biologically Active Substance|Hospital Course|12314,12323|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Element, Ion, or Isotope|Hospital Course|12314,12323|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Food|Hospital Course|12314,12323|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Inorganic Chemical|Hospital Course|12314,12323|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Pharmacologic Substance|Hospital Course|12314,12323|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Event|Event|Hospital Course|12314,12323|false|false|false|||potassium
Finding|Physiologic Function|Hospital Course|12314,12323|false|false|false|C4553027|Potassium metabolic function|potassium
Procedure|Laboratory Procedure|Hospital Course|12314,12323|false|false|false|C0202194|Potassium measurement|potassium
Drug|Inorganic Chemical|Hospital Course|12314,12332|false|false|false|C0032825|potassium chloride|potassium chloride
Drug|Pharmacologic Substance|Hospital Course|12314,12332|false|false|false|C0032825|potassium chloride|potassium chloride
Drug|Element, Ion, or Isotope|Hospital Course|12324,12332|false|false|false|C0008203;C0596019|Chlorides;chloride ion|chloride
Event|Event|Hospital Course|12324,12332|false|false|false|||chloride
Finding|Physiologic Function|Hospital Course|12324,12332|false|false|false|C4553021|Chloride metabolic function|chloride
Procedure|Laboratory Procedure|Hospital Course|12324,12332|false|false|false|C0201952|Chloride measurement|chloride
Finding|Functional Concept|Hospital Course|12352,12360|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|12355,12360|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|12355,12360|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Intellectual Product|Hospital Course|12361,12365|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|12361,12371|false|false|false|C3537736|Once A Day|once a day
Event|Event|Hospital Course|12368,12371|false|false|false|||day
Finding|Idea or Concept|Hospital Course|12368,12371|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|12368,12371|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biomedical or Dental Material|Hospital Course|12383,12389|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|12390,12397|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|12390,12397|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|12406,12411|false|false|false|C2369992|Align|Align
Drug|Pharmacologic Substance|Hospital Course|12406,12411|false|false|false|C2369992|Align|Align
Drug|Pharmacologic Substance|Hospital Course|12413,12437|false|false|false|C4019097|herbal medicines bifidobacterium infantis|bifidobacterium infantis
Event|Event|Hospital Course|12429,12437|false|false|false|||infantis
Anatomy|Body Space or Junction|Hospital Course|12444,12448|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|12444,12448|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|12444,12448|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|12444,12448|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|Hospital Course|12449,12454|false|false|false|||DAILY
Drug|Organic Chemical|Hospital Course|12461,12471|false|false|false|C0002598|amiodarone|Amiodarone
Drug|Pharmacologic Substance|Hospital Course|12461,12471|false|false|false|C0002598|amiodarone|Amiodarone
Event|Event|Hospital Course|12461,12471|false|false|false|||Amiodarone
Procedure|Laboratory Procedure|Hospital Course|12461,12471|false|false|false|C5399868|Drug assay amiodarone|Amiodarone
Drug|Organic Chemical|Hospital Course|12494,12502|false|false|false|C1831808|apixaban|Apixaban
Drug|Pharmacologic Substance|Hospital Course|12494,12502|false|false|false|C1831808|apixaban|Apixaban
Disorder|Mental or Behavioral Dysfunction|Hospital Course|12513,12516|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12513,12516|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|12513,12516|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|12513,12516|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|12513,12516|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|12523,12530|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Hospital Course|12523,12530|false|false|false|C0004057|aspirin|Aspirin
Drug|Biologically Active Substance|Hospital Course|12552,12560|false|false|false|C0009235|Coenzymes|coenzyme
Drug|Organic Chemical|Hospital Course|12552,12560|false|false|false|C0009235|Coenzymes|coenzyme
Event|Event|Hospital Course|12552,12560|false|false|false|||coenzyme
Drug|Biologically Active Substance|Hospital Course|12552,12564|false|false|false|C0041536|ubidecarenone|coenzyme Q10
Drug|Organic Chemical|Hospital Course|12552,12564|false|false|false|C0041536|ubidecarenone|coenzyme Q10
Drug|Pharmacologic Substance|Hospital Course|12552,12564|false|false|false|C0041536|ubidecarenone|coenzyme Q10
Event|Event|Hospital Course|12561,12564|false|false|false|||Q10
Finding|Gene or Genome|Hospital Course|12561,12564|false|false|false|C1414333;C2827473|AGO2 gene;AGO2 wt Allele|Q10
Anatomy|Body Space or Junction|Hospital Course|12572,12576|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|12572,12576|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|12572,12576|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|12572,12576|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|Hospital Course|12577,12582|false|false|false|||DAILY
Drug|Organic Chemical|Hospital Course|12589,12597|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|12589,12597|false|false|false|C1692318|docusate|Docusate
Event|Event|Hospital Course|12589,12597|false|false|false|||Docusate
Drug|Organic Chemical|Hospital Course|12589,12604|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|Hospital Course|12589,12604|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|Hospital Course|12598,12604|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|12598,12604|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|12598,12604|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|12598,12604|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|12598,12604|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|12598,12604|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|Hospital Course|12615,12618|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12615,12618|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|12615,12618|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|12615,12618|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|12615,12618|false|false|false|C1332410|BID gene|BID
Drug|Element, Ion, or Isotope|Hospital Course|12625,12632|false|false|false|C2346592|Ferrous|Ferrous
Drug|Inorganic Chemical|Hospital Course|12625,12640|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Pharmacologic Substance|Hospital Course|12625,12640|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Element, Ion, or Isotope|Hospital Course|12633,12640|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Inorganic Chemical|Hospital Course|12633,12640|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Pharmacologic Substance|Hospital Course|12633,12640|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Event|Event|Hospital Course|12633,12640|false|false|false|||Sulfate
Drug|Organic Chemical|Hospital Course|12663,12668|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|Hospital Course|12663,12668|false|false|false|C3489575|sennosides, USP|Senna
Drug|Organic Chemical|Hospital Course|12690,12700|false|false|false|C0074393|sertraline|Sertraline
Drug|Pharmacologic Substance|Hospital Course|12690,12700|false|false|false|C0074393|sertraline|Sertraline
Drug|Organic Chemical|Hospital Course|12723,12733|false|false|false|C0257343|tamsulosin|Tamsulosin
Drug|Pharmacologic Substance|Hospital Course|12723,12733|false|false|false|C0257343|tamsulosin|Tamsulosin
Drug|Organic Chemical|Hospital Course|12753,12763|false|false|false|C0257343|tamsulosin|tamsulosin
Drug|Pharmacologic Substance|Hospital Course|12753,12763|false|false|false|C0257343|tamsulosin|tamsulosin
Event|Event|Hospital Course|12753,12763|false|false|false|||tamsulosin
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12773,12780|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|Hospital Course|12773,12780|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|Hospital Course|12773,12780|false|false|false|C0006935|capsule (pharmacologic)|capsule
Finding|Functional Concept|Hospital Course|12784,12792|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|12787,12792|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|12787,12792|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12812,12819|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|12812,12819|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|12812,12819|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Event|Event|Hospital Course|12820,12827|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|12820,12827|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|12837,12846|false|false|false|C0076840|torsemide|Torsemide
Drug|Pharmacologic Substance|Hospital Course|12837,12846|false|false|false|C0076840|torsemide|Torsemide
Drug|Organic Chemical|Hospital Course|12869,12876|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|12869,12876|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|12869,12876|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|Hospital Course|12869,12878|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|Hospital Course|12869,12878|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|Hospital Course|12869,12878|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|Hospital Course|12869,12878|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|Hospital Course|12869,12878|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|Hospital Course|12884,12888|false|false|false|||UNIT
Event|Event|Hospital Course|12903,12912|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|12903,12912|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|12903,12912|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|12903,12912|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|12903,12912|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|12903,12924|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|12903,12924|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|12913,12924|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|12913,12924|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|12913,12924|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|Hospital Course|12926,12930|false|false|false|||Home
Finding|Idea or Concept|Hospital Course|12926,12930|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|12926,12930|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|12926,12930|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|Hospital Course|12936,12943|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|Hospital Course|12936,12943|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|Hospital Course|12946,12954|false|false|false|||Facility
Finding|Intellectual Product|Hospital Course|12946,12954|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|Hospital Course|12962,12971|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|12962,12971|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|12962,12971|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|12962,12971|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|12962,12971|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|12962,12981|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|12972,12981|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|12972,12981|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|12972,12981|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|12972,12981|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|12972,12981|false|false|false|C0011900|Diagnosis|Diagnosis
Event|Event|Principle Diagnosis|13025,13039|false|false|false|||excerterbation
Disorder|Neoplastic Process|Principle Diagnosis|13041,13050|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Finding|Functional Concept|Principle Diagnosis|13041,13050|false|false|false|C1522484|metastatic qualifier|Secondary
Attribute|Clinical Attribute|Principle Diagnosis|13041,13060|false|false|false|C4255018||Secondary diagnosis
Finding|Finding|Principle Diagnosis|13041,13060|false|false|false|C0332138|Secondary diagnosis|Secondary diagnosis
Attribute|Clinical Attribute|Principle Diagnosis|13051,13060|false|false|false|C0945731||diagnosis
Event|Event|Principle Diagnosis|13051,13060|false|false|false|||diagnosis
Finding|Classification|Principle Diagnosis|13051,13060|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|Principle Diagnosis|13051,13060|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|Principle Diagnosis|13051,13060|false|false|false|C0011900|Diagnosis|diagnosis
Event|Event|Principle Diagnosis|13081,13094|false|false|false|||Transaminitis
Finding|Finding|Principle Diagnosis|13081,13094|false|false|false|C2242708|Hypertransaminasaemia|Transaminitis
Finding|Functional Concept|Principle Diagnosis|13095,13105|false|false|false|C0036525;C1522484|Metastatic to;metastatic qualifier|Metastatic
Disorder|Neoplastic Process|Principle Diagnosis|13095,13114|false|false|false|C0278883|Metastatic melanoma|Metastatic melanoma
Disorder|Neoplastic Process|Principle Diagnosis|13106,13114|false|false|false|C0025202|melanoma|melanoma
Drug|Immunologic Factor|Principle Diagnosis|13106,13114|false|false|false|C0796561|Melanoma vaccine|melanoma
Drug|Pharmacologic Substance|Principle Diagnosis|13106,13114|false|false|false|C0796561|Melanoma vaccine|melanoma
Event|Event|Principle Diagnosis|13106,13114|false|false|false|||melanoma
Disorder|Disease or Syndrome|Principle Diagnosis|13115,13118|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Event|Event|Principle Diagnosis|13115,13118|false|false|false|||CKD
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|13119,13127|false|false|false|C0018787|Heart|Coronary
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|13119,13134|false|false|false|C0205042|Coronary artery|Coronary artery
Disorder|Disease or Syndrome|Principle Diagnosis|13119,13142|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|Coronary artery disease
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|13128,13134|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|Principle Diagnosis|13128,13134|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Disorder|Disease or Syndrome|Principle Diagnosis|13128,13142|false|false|false|C0852949|Arteriopathic disease|artery disease
Disorder|Disease or Syndrome|Principle Diagnosis|13135,13142|false|false|false|C0012634|Disease|disease
Event|Event|Principle Diagnosis|13135,13142|false|false|false|||disease
Event|Event|Principle Diagnosis|13148,13152|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|Principle Diagnosis|13148,13152|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|13157,13160|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|Principle Diagnosis|13157,13160|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|Principle Diagnosis|13157,13160|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Drug|Amino Acid, Peptide, or Protein|Principle Diagnosis|13161,13164|false|false|false|C2713669|SERPINA5 protein, human|PCI
Drug|Biologically Active Substance|Principle Diagnosis|13161,13164|false|false|false|C2713669|SERPINA5 protein, human|PCI
Event|Event|Principle Diagnosis|13161,13164|false|false|false|||PCI
Finding|Gene or Genome|Principle Diagnosis|13161,13164|false|false|false|C1418370;C1705930;C4049621|Peritoneal Cancer Index;SERPINA5 gene;SERPINA5 wt Allele|PCI
Finding|Intellectual Product|Principle Diagnosis|13161,13164|false|false|false|C1418370;C1705930;C4049621|Peritoneal Cancer Index;SERPINA5 gene;SERPINA5 wt Allele|PCI
Procedure|Therapeutic or Preventive Procedure|Principle Diagnosis|13161,13164|false|false|false|C1514496;C1532338;C4724254|Percutaneous Coronary Intervention;Prophylactic Cranial Irradiation;photochemical internalization|PCI
Finding|Mental Process|Discharge Condition|13189,13195|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|13189,13202|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|13189,13202|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|13196,13202|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|13196,13202|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|13204,13209|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|13204,13209|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|13214,13222|false|false|false|||coherent
Finding|Finding|Discharge Condition|13214,13222|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|13224,13229|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|13224,13246|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|13224,13246|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|13233,13246|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|13233,13246|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|13233,13246|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|13248,13253|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|13248,13253|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|13248,13253|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|13248,13253|false|false|false|||Alert
Finding|Finding|Discharge Condition|13248,13253|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|13248,13253|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|13248,13253|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|13258,13269|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|13258,13269|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|13271,13279|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|13271,13279|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|13271,13279|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|13280,13286|false|false|false|C5889824||Status
Event|Event|Discharge Condition|13280,13286|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|13280,13286|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|Discharge Condition|13288,13298|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|13288,13298|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|13288,13298|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|13288,13298|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|13301,13309|false|false|false|||requires
Event|Event|Discharge Condition|13310,13320|false|false|false|||assistance
Finding|Social Behavior|Discharge Condition|13310,13320|false|false|false|C0018896|Helping Behavior|assistance
Drug|Amino Acid, Peptide, or Protein|Discharge Condition|13324,13327|false|false|false|C1454018|AICDA protein, human|aid
Drug|Enzyme|Discharge Condition|13324,13327|false|false|false|C1454018|AICDA protein, human|aid
Event|Event|Discharge Condition|13324,13327|false|false|false|||aid
Finding|Gene or Genome|Discharge Condition|13324,13327|false|false|false|C1421876;C3540469|AICDA gene;AICDA wt Allele|aid
Procedure|Therapeutic or Preventive Procedure|Discharge Condition|13324,13327|false|false|false|C0021588;C0280108|AID - Artificial insemination by donor;dacarbazine/doxorubicin/ifosfamide protocol|aid
Event|Event|Discharge Condition|13329,13335|false|false|false|||walker
Finding|Gene or Genome|Discharge Instructions|13457,13461|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|Discharge Instructions|13484,13492|false|false|false|||pleasure
Finding|Intellectual Product|Discharge Instructions|13484,13492|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|Discharge Instructions|13484,13492|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|Discharge Instructions|13500,13504|false|false|false|C1947933|care activity|care
Event|Event|Discharge Instructions|13500,13504|false|false|false|||care
Finding|Finding|Discharge Instructions|13500,13504|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|13500,13504|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|13500,13507|false|false|false|C1555558|care of - AddressPartType|care of
Event|Event|Discharge Instructions|13532,13535|false|false|false|||WAS
Event|Event|Discharge Instructions|13538,13546|false|false|false|||ADMITTED
Event|Event|Discharge Instructions|13554,13562|false|false|false|||HOSPITAL
Finding|Idea or Concept|Discharge Instructions|13554,13562|false|false|false|C1547192|Organization unit type - Hospital|HOSPITAL
Event|Event|Discharge Instructions|13575,13582|false|false|false|||feeling
Finding|Sign or Symptom|Discharge Instructions|13583,13598|false|false|false|C0013404|Dyspnea|short of breath
Event|Event|Discharge Instructions|13592,13598|false|false|false|||breath
Finding|Body Substance|Discharge Instructions|13592,13598|false|false|false|C0225386|Breath|breath
Drug|Substance|Discharge Instructions|13615,13620|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|Discharge Instructions|13615,13620|false|false|false|||fluid
Finding|Intellectual Product|Discharge Instructions|13615,13620|false|false|false|C1546638|Fluid Specimen Code|fluid
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|13630,13635|false|false|false|C0024109|Lung|lungs
Event|Event|Discharge Instructions|13646,13652|false|false|false|||caused
Attribute|Clinical Attribute|Discharge Instructions|13658,13667|false|false|false|C3864998||condition
Disorder|Disease or Syndrome|Discharge Instructions|13658,13667|false|false|false|C0012634|Disease|condition
Event|Event|Discharge Instructions|13658,13667|false|false|false|||condition
Finding|Conceptual Entity|Discharge Instructions|13658,13667|false|false|false|C1705253|Logical Condition|condition
Event|Event|Discharge Instructions|13668,13674|false|false|false|||called
Event|Event|Discharge Instructions|13679,13686|false|false|false|||failure
Finding|Functional Concept|Discharge Instructions|13679,13686|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|Discharge Instructions|13679,13686|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|Discharge Instructions|13679,13686|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|Discharge Instructions|13713,13717|true|false|false|||pump
Event|Event|Discharge Instructions|13723,13729|true|false|false|||enough
Drug|Substance|Discharge Instructions|13734,13739|true|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|Discharge Instructions|13734,13739|true|false|false|||fluid
Finding|Intellectual Product|Discharge Instructions|13734,13739|true|false|false|C1546638|Fluid Specimen Code|fluid
Anatomy|Body Location or Region|Discharge Instructions|13740,13745|true|false|false|C0004600||backs
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|13760,13765|false|false|false|C0024109|Lung|lungs
Event|Activity|Discharge Instructions|13775,13783|false|false|false|C1709305|Occur (action)|HAPPENED
Event|Event|Discharge Instructions|13792,13795|false|false|false|||WAS
Finding|Idea or Concept|Discharge Instructions|13803,13811|false|false|false|C1547192|Organization unit type - Hospital|HOSPITAL
Attribute|Clinical Attribute|Discharge Instructions|13830,13841|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|13830,13841|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|13830,13841|false|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|13830,13841|false|false|false|C4284232|Medications|medications
Event|Event|Discharge Instructions|13845,13849|false|false|false|||help
Event|Event|Discharge Instructions|13850,13853|false|false|false|||get
Drug|Substance|Discharge Instructions|13858,13863|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|Discharge Instructions|13858,13863|false|false|false|||fluid
Finding|Intellectual Product|Discharge Instructions|13858,13863|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|Discharge Instructions|13875,13884|false|false|false|||breathing
Event|Event|Discharge Instructions|13889,13895|false|false|false|||better
Finding|Idea or Concept|Discharge Instructions|13889,13895|false|false|false|C1550462|Observation Interpretation - better|better
Event|Event|Discharge Instructions|13905,13910|false|false|false|||ready
Event|Event|Discharge Instructions|13914,13919|false|false|false|||leave
Event|Event|Discharge Instructions|13924,13932|false|false|false|||hospital
Finding|Idea or Concept|Discharge Instructions|13924,13932|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|Discharge Instructions|13945,13948|false|false|false|||YOU
Event|Event|Discharge Instructions|13949,13953|false|false|false|||NEED
Finding|Functional Concept|Discharge Instructions|13949,13953|false|false|false|C0686904|Patient need for (contextual qualifier)|NEED
Event|Event|Discharge Instructions|13957,13959|false|false|false|||DO
Event|Event|Discharge Instructions|13969,13974|false|false|false|||LEAVE
Event|Event|Discharge Instructions|13979,13987|false|false|false|||HOSPITAL
Finding|Idea or Concept|Discharge Instructions|13979,13987|false|false|false|C1547192|Organization unit type - Hospital|HOSPITAL
Event|Event|Discharge Instructions|13993,13997|false|false|false|||Take
Attribute|Clinical Attribute|Discharge Instructions|14010,14021|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|14010,14021|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|14010,14021|false|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|14010,14021|false|false|false|C4284232|Medications|medications
Event|Event|Discharge Instructions|14025,14035|false|false|false|||prescribed
Finding|Functional Concept|Discharge Instructions|14055,14061|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|Follow
Finding|Intellectual Product|Discharge Instructions|14055,14061|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|Follow
Finding|Finding|Discharge Instructions|14055,14064|false|false|false|C0589120|Follow-up status|Follow up
Procedure|Health Care Activity|Discharge Instructions|14055,14064|false|false|false|C1522577|follow-up|Follow up
Event|Event|Discharge Instructions|14062,14064|false|false|false|||up
Attribute|Clinical Attribute|Discharge Instructions|14138,14144|false|false|false|C0944911||weight
Event|Event|Discharge Instructions|14138,14144|false|false|false|||weight
Finding|Finding|Discharge Instructions|14138,14144|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|Discharge Instructions|14138,14144|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|Discharge Instructions|14138,14144|false|false|false|C1305866|Weighing patient|weight
Event|Event|Discharge Instructions|14148,14157|false|false|false|||discharge
Finding|Body Substance|Discharge Instructions|14148,14157|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Discharge Instructions|14148,14157|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Discharge Instructions|14148,14157|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Discharge Instructions|14148,14157|false|false|false|C0030685|Patient Discharge|discharge
Procedure|Laboratory Procedure|Discharge Instructions|14169,14172|false|false|false|C3161851|liquid-based cytology (procedure)|lbs
Event|Event|Discharge Instructions|14174,14178|false|false|false|||Call
Event|Event|Discharge Instructions|14184,14190|false|false|false|||doctor
Finding|Intellectual Product|Discharge Instructions|14184,14190|false|false|false|C2348314|Doctor - Title|doctor
Attribute|Clinical Attribute|Discharge Instructions|14199,14205|false|false|false|C0944911||weight
Event|Event|Discharge Instructions|14199,14205|false|false|false|||weight
Finding|Finding|Discharge Instructions|14199,14205|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|Discharge Instructions|14199,14205|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|Discharge Instructions|14199,14205|false|false|false|C1305866|Weighing patient|weight
Event|Event|Discharge Instructions|14206,14210|false|false|false|||goes
Event|Event|Discharge Instructions|14227,14233|false|false|false|||pounds
Event|Event|Discharge Instructions|14237,14241|false|false|false|||Call
Finding|Functional Concept|Discharge Instructions|14237,14241|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|Call
Finding|Gene or Genome|Discharge Instructions|14237,14241|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|Call
Finding|Intellectual Product|Discharge Instructions|14237,14241|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|Call
Finding|Mental Process|Discharge Instructions|14237,14241|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|Call
Event|Event|Discharge Instructions|14246,14252|false|false|false|||doctor
Event|Event|Discharge Instructions|14260,14266|true|false|false|||notice
Finding|Gene or Genome|Discharge Instructions|14279,14285|true|false|false|C1428845|ITPRIP gene|danger
Event|Event|Discharge Instructions|14286,14291|true|false|false|||signs
Finding|Finding|Discharge Instructions|14286,14291|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Discharge Instructions|14286,14291|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Disorder|Disease or Syndrome|Discharge Instructions|14321,14325|false|false|false|C0339510|Vitelliform Macular Dystrophy|best
Event|Event|Discharge Instructions|14321,14325|false|false|false|||best
Finding|Gene or Genome|Discharge Instructions|14321,14325|false|false|false|C1826421;C5781213|BEST1 gene;BEST1 wt Allele|best
Event|Activity|Discharge Instructions|14338,14342|false|false|false|C1947933|care activity|Care
Finding|Finding|Discharge Instructions|14338,14342|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Discharge Instructions|14338,14342|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Attribute|Clinical Attribute|Discharge Instructions|14338,14347|false|false|false|C4321316||Care Team
Finding|Finding|Discharge Instructions|14338,14347|false|false|false|C4321315|Care team|Care Team
Procedure|Health Care Activity|Discharge Instructions|14353,14361|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|14362,14374|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|14362,14374|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|14362,14374|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

