 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Procedure|Health Care Activity|SIMPLE_SEGMENT|52,61|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|52,66|false|false|false|C2598112||Admission Date
Finding|Body Substance|SIMPLE_SEGMENT|86,95|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|86,95|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|86,95|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|86,95|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|86,100|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|118,123|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|118,123|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|118,123|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|142,145|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|142,145|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|142,145|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|142,145|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|142,145|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|153,160|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|153,160|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|162,170|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|Allergies|188,197|true|false|false|C1717415||Allergies
Finding|Pathologic Function|Allergies|188,197|true|false|false|C0020517|Hypersensitivity|Allergies
Finding|Functional Concept|Allergies|206,210|false|false|false|C0016094;C1522646;C1555017|File (record);Filed;URL Scheme - File|File
Finding|Intellectual Product|Allergies|206,210|false|false|false|C0016094;C1522646;C1555017|File (record);Filed;URL Scheme - File|File
Finding|Functional Concept|Allergies|213,222|false|false|false|C1999232|Attending (action)|Attending
Anatomy|Body Location or Region|Chief Complaint|248,253|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Chief Complaint|248,253|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Chief Complaint|248,258|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Chief Complaint|248,258|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Chief Complaint|254,258|false|true|false|C2598155||pain
Finding|Functional Concept|Chief Complaint|254,258|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Chief Complaint|254,258|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Classification|Chief Complaint|261,266|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|267,275|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|267,275|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|279,297|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|288,297|false|false|false|C0945766||Procedure
Event|Occupational Activity|Chief Complaint|288,297|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|288,297|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|288,297|false|false|false|C0184661|Interventional procedure|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|313,331|false|false|false|C0191234|Pericardiocentesis|pericardiocentesis
Finding|Conceptual Entity|History of Present Illness|371,378|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|HISTORY
Finding|Finding|History of Present Illness|371,378|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|HISTORY
Finding|Functional Concept|History of Present Illness|371,378|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|HISTORY
Finding|Finding|History of Present Illness|371,381|false|false|false|C0262926|Medical History|HISTORY OF
Finding|Idea or Concept|History of Present Illness|382,392|true|false|false|C0449450|Presentation|PRESENTING
Finding|Sign or Symptom|History of Present Illness|393,400|false|false|false|C0221423|Illness (finding)|ILLNESS
Finding|Finding|History of Present Illness|419,423|false|false|false|C1706180|Male Gender|male
Disorder|Disease or Syndrome|History of Present Illness|429,449|false|false|false|C0003873|Rheumatoid Arthritis|rheumatoid arthritis
Disorder|Disease or Syndrome|History of Present Illness|440,449|false|false|false|C0003864|Arthritis|arthritis
Drug|Pharmacologic Substance|History of Present Illness|451,456|false|false|false|C0242708|Antirheumatic Drugs, Disease-Modifying|DMARD
Event|Event|History of Present Illness|457,464|false|false|false|C0019843|Holidays|holiday
Finding|Intellectual Product|History of Present Illness|478,483|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|brief
Procedure|Health Care Activity|History of Present Illness|484,499|false|false|false|C0019993|Hospitalization|hospitalization
Disorder|Disease or Syndrome|History of Present Illness|516,528|false|false|false|C0031046|Pericarditis|pericarditis
Finding|Idea or Concept|History of Present Illness|551,559|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Finding|History of Present Illness|565,573|false|false|false|C0332148|Probable diagnosis|probable
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|574,581|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|History of Present Illness|574,581|false|true|false|C1314974|Cardiac attachment|cardiac
Disorder|Disease or Syndrome|History of Present Illness|574,591|false|true|false|C0007177|Cardiac Tamponade|cardiac tamponade
Finding|Functional Concept|History of Present Illness|582,591|false|true|false|C0332459|Compressed structure|tamponade
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|582,591|false|true|false|C0579016||tamponade
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|609,627|false|false|false|C0191234|Pericardiocentesis|pericardiocentesis
Drug|Substance|History of Present Illness|633,638|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|History of Present Illness|633,638|false|false|false|C1546604|Drain Specimen Code|drain
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|633,648|false|false|false|C3495845|Drain placement|drain placement
Procedure|Health Care Activity|History of Present Illness|639,648|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|639,648|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Finding|Functional Concept|History of Present Illness|658,666|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|History of Present Illness|658,666|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|History of Present Illness|658,666|false|false|false|C4706767|Transfer (immobility management)|transfer
Finding|Body Substance|History of Present Illness|681,688|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|681,688|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|681,688|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|725,730|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Sign or Symptom|History of Present Illness|731,751|false|false|false|C0008033|Pleuritic pain|pleuritic chest pain
Anatomy|Body Location or Region|History of Present Illness|741,746|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|741,746|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|741,751|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|741,751|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|747,751|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|747,751|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|747,751|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Idea or Concept|History of Present Illness|759,762|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|History of Present Illness|759,762|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Pharmacologic Substance|History of Present Illness|763,771|false|false|false|C0720099|Duration brand of oxymetazoline|duration
Finding|Idea or Concept|History of Present Illness|779,786|false|false|false|C0449255;C0542559;C4281677|Application Context;Context;contextual factors|context
Finding|Intellectual Product|History of Present Illness|779,786|false|false|false|C0449255;C0542559;C4281677|Application Context;Context;contextual factors|context
Finding|Mental Process|History of Present Illness|779,786|false|false|false|C0449255;C0542559;C4281677|Application Context;Context;contextual factors|context
Finding|Sign or Symptom|History of Present Illness|807,814|false|false|false|C0015672|Fatigue|fatigue
Finding|Sign or Symptom|History of Present Illness|816,823|false|false|false|C0231218|Malaise|malaise
Attribute|Clinical Attribute|History of Present Illness|831,842|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|History of Present Illness|831,842|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|History of Present Illness|831,842|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|History of Present Illness|831,842|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|History of Present Illness|843,851|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|History of Present Illness|843,851|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Drug|Organic Chemical|History of Present Illness|872,877|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|872,877|false|false|false|C3815497|Cough (guaifenesin)|cough
Finding|Sign or Symptom|History of Present Illness|872,877|false|false|false|C0010200|Coughing|cough
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|885,888|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Finding|Gene or Genome|History of Present Illness|885,888|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|History of Present Illness|885,888|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|900,909|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|History of Present Illness|900,909|false|false|false|C2707265||pulmonary
Finding|Finding|History of Present Illness|900,909|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|History of Present Illness|900,918|false|false|false|C0034065|Pulmonary Embolism|pulmonary embolism
Finding|Finding|History of Present Illness|910,918|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Finding|Pathologic Function|History of Present Illness|910,918|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|930,941|false|false|false|C0031050|Pericardial sac structure|pericardium
Finding|Body Substance|History of Present Illness|952,960|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|History of Present Illness|952,960|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|History of Present Illness|952,960|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Disorder|Disease or Syndrome|History of Present Illness|985,997|false|false|false|C0031046|Pericarditis|pericarditis
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|999,1002|false|false|false|C0018064|Equine Gonadotropins|ECG
Drug|Hormone|History of Present Illness|999,1002|false|false|false|C0018064|Equine Gonadotropins|ECG
Drug|Pharmacologic Substance|History of Present Illness|999,1002|false|false|false|C0018064|Equine Gonadotropins|ECG
Finding|Intellectual Product|History of Present Illness|999,1002|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|ECG
Procedure|Diagnostic Procedure|History of Present Illness|999,1002|false|false|false|C1623258|Electrocardiography|ECG
Disorder|Disease or Syndrome|History of Present Illness|1057,1069|false|false|false|C0031046|Pericarditis|pericarditis
Procedure|Diagnostic Procedure|History of Present Illness|1071,1085|false|false|false|C0013516|Echocardiography|Echocardiogram
Finding|Body Substance|History of Present Illness|1102,1110|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|History of Present Illness|1102,1110|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|History of Present Illness|1102,1110|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Functional Concept|History of Present Illness|1134,1143|false|false|false|C0332459|Compressed structure|tamponade
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1134,1143|false|false|false|C0579016||tamponade
Finding|Idea or Concept|History of Present Illness|1189,1192|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|History of Present Illness|1189,1192|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|History of Present Illness|1198,1207|false|false|false|C0020740|ibuprofen|ibuprofen
Drug|Pharmacologic Substance|History of Present Illness|1198,1207|false|false|false|C0020740|ibuprofen|ibuprofen
Drug|Organic Chemical|History of Present Illness|1223,1233|false|false|false|C0009262|colchicine|colchicine
Drug|Pharmacologic Substance|History of Present Illness|1223,1233|false|false|false|C0009262|colchicine|colchicine
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|1241,1244|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1241,1244|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|History of Present Illness|1241,1244|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|History of Present Illness|1241,1244|false|false|false|C1332410|BID gene|BID
Finding|Mental Process|History of Present Illness|1253,1264|false|false|false|C0546816|Persistence|persistence
Disorder|Disease or Syndrome|History of Present Illness|1268,1273|false|false|false|C1446899|minor (disease)|minor
Finding|Gene or Genome|History of Present Illness|1268,1273|false|false|false|C1417837;C3272493|NR4A3 gene;NR4A3 wt Allele|minor
Anatomy|Body Location or Region|History of Present Illness|1284,1289|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|1284,1289|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|1290,1294|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|1290,1294|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1290,1294|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|History of Present Illness|1395,1401|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|History of Present Illness|1395,1401|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Attribute|Clinical Attribute|History of Present Illness|1415,1419|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|1415,1419|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1415,1419|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Location or Region|History of Present Illness|1431,1441|false|false|false|C0230134|Structure of precordium|precordium
Anatomy|Body Location or Region|History of Present Illness|1462,1470|false|false|false|C0037004;C4299050|Shoulder;Upper extremity>Shoulder|shoulder
Procedure|Diagnostic Procedure|History of Present Illness|1462,1470|false|false|false|C0221590;C0869975|Examination of shoulder(s);Procedures on Shoulder|shoulder
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1462,1470|false|false|false|C0221590;C0869975|Examination of shoulder(s);Procedures on Shoulder|shoulder
Finding|Finding|History of Present Illness|1509,1512|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|History of Present Illness|1509,1512|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Anatomy|Body Location or Region|History of Present Illness|1535,1540|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|1535,1540|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|1541,1545|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|1541,1545|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1541,1545|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Social Behavior|History of Present Illness|1557,1565|false|false|false|C0019421|Heterosexuality|straight
Finding|Intellectual Product|History of Present Illness|1583,1587|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Finding|History of Present Illness|1595,1603|false|false|false|C0277854|dyspneic|dyspneic
Event|Activity|History of Present Illness|1627,1631|false|false|false|C1947933|care activity|care
Finding|Finding|History of Present Illness|1627,1631|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|History of Present Illness|1627,1631|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Pathologic Function|History of Present Illness|1651,1662|false|false|false|C0857353|Hypotensive|hypotensive
Attribute|Clinical Attribute|History of Present Illness|1668,1671|false|false|false|C0871470|Systolic Pressure|SBP
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1668,1671|false|false|false|C0085805|Androgen Binding Protein|SBP
Drug|Biologically Active Substance|History of Present Illness|1668,1671|false|false|false|C0085805|Androgen Binding Protein|SBP
Finding|Gene or Genome|History of Present Illness|1668,1671|false|false|false|C1705296;C3274833|CCHCR1 wt Allele;SHBG wt Allele|SBP
Procedure|Diagnostic Procedure|History of Present Illness|1668,1671|false|false|false|C1306620|Systolic blood pressure measurement|SBP
Finding|Intellectual Product|History of Present Illness|1682,1687|false|false|false|C3542016|Concept model range (foundation metadata concept)|range
Finding|Intellectual Product|History of Present Illness|1726,1730|false|false|false|C1547225|Mild Severity of Illness Code|mild
Attribute|Clinical Attribute|History of Present Illness|1731,1742|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|History of Present Illness|1731,1742|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|History of Present Illness|1731,1742|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|History of Present Illness|1731,1742|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Sign or Symptom|History of Present Illness|1731,1751|false|false|false|C0476273|Respiratory distress|respiratory distress
Finding|Finding|History of Present Illness|1743,1751|false|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|History of Present Illness|1743,1751|false|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Cell Function|History of Present Illness|1757,1768|false|false|false|C0231940;C0282636|Alveolar ventilation function;Cell Respiration|oxygenation
Finding|Organ or Tissue Function|History of Present Illness|1757,1768|false|false|false|C0231940;C0282636|Alveolar ventilation function;Cell Respiration|oxygenation
Drug|Substance|History of Present Illness|1821,1826|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|History of Present Illness|1821,1826|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Functional Concept|History of Present Illness|1843,1852|false|false|false|C0332459|Compressed structure|tamponade
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1843,1852|false|false|false|C0579016||tamponade
Finding|Intellectual Product|History of Present Illness|1876,1880|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Procedure|Diagnostic Procedure|History of Present Illness|1900,1914|false|false|false|C0013516|Echocardiography|echocardiogram
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1916,1934|false|false|false|C0191234|Pericardiocentesis|Pericardiocentesis
Finding|Body Substance|History of Present Illness|1961,1973|false|false|false|C0682554|Serous fluid|serous fluid
Drug|Substance|History of Present Illness|1968,1973|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|History of Present Illness|1968,1973|false|false|false|C1546638|Fluid Specimen Code|fluid
Anatomy|Body Location or Region|History of Present Illness|1980,1991|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1980,1991|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Drug|Substance|History of Present Illness|1992,1997|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|History of Present Illness|1992,1997|false|false|false|C1546604|Drain Specimen Code|drain
Finding|Organ or Tissue Function|History of Present Illness|2010,2022|false|false|false|C0019010|Hemodynamics|Hemodynamics
Procedure|Laboratory Procedure|History of Present Illness|2010,2022|false|false|false|C4281788|hemodynamics (procedure)|Hemodynamics
Event|Activity|History of Present Illness|2044,2051|false|false|false|C1706079||arrival
Finding|Functional Concept|History of Present Illness|2044,2051|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Finding|Body Substance|History of Present Illness|2063,2070|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|2063,2070|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|2063,2070|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|History of Present Illness|2082,2104|false|false|false|C0578150|Hemodynamically stable|hemodynamically stable
Finding|Intellectual Product|History of Present Illness|2098,2104|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Intellectual Product|History of Present Illness|2113,2117|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Finding|History of Present Illness|2121,2129|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|History of Present Illness|2121,2129|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Attribute|Clinical Attribute|History of Present Illness|2130,2141|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|History of Present Illness|2130,2141|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|History of Present Illness|2130,2141|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|History of Present Illness|2130,2141|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Sign or Symptom|History of Present Illness|2130,2150|false|false|false|C0476273|Respiratory distress|respiratory distress
Finding|Finding|History of Present Illness|2142,2150|false|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|History of Present Illness|2142,2150|false|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Drug|Organic Chemical|History of Present Illness|2191,2196|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|History of Present Illness|2191,2196|false|false|false|C0699992|Lasix|Lasix
Procedure|Diagnostic Procedure|History of Present Illness|2215,2229|false|false|false|C0013516|Echocardiography|echocardiogram
Finding|Functional Concept|History of Present Illness|2261,2271|false|false|false|C0332299|Suggestive of|suggestive
Finding|Functional Concept|History of Present Illness|2261,2274|false|false|false|C0332299|Suggestive of|suggestive of
Finding|Body Substance|History of Present Illness|2291,2299|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|History of Present Illness|2291,2299|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|History of Present Illness|2291,2299|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Body Substance|History of Present Illness|2313,2320|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|2313,2320|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|2313,2320|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Disorder|Disease or Syndrome|History of Present Illness|2341,2345|false|false|false|C0080151|Simian Acquired Immunodeficiency Syndrome|said
Anatomy|Body Location or Region|History of Present Illness|2346,2351|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|2346,2351|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|2346,2356|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|2346,2356|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|2352,2356|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|2352,2356|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|2352,2356|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|History of Present Illness|2362,2369|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|History of Present Illness|2362,2369|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Functional Concept|History of Present Illness|2387,2397|false|false|false|C1524062|Additional|additional
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2468,2475|false|false|false|C0018787|Heart|Cardiac
Finding|Intellectual Product|Past Medical History|2468,2475|false|false|false|C1314974|Cardiac attachment|Cardiac
Disorder|Disease or Syndrome|Patient History|2488,2500|false|false|false|C0031046|Pericarditis|Pericarditis
Finding|Idea or Concept|Patient History|2505,2510|false|false|false|C1552828|Table Frame - above|above
Disorder|Disease or Syndrome|Patient History|2513,2525|false|false|false|C0020538|Hypertensive disease|Hypertension
Disorder|Disease or Syndrome|Patient History|2528,2540|false|false|false|C0242339|Dyslipidemias|Dyslipidemia
Finding|Finding|Patient History|2552,2555|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|PMH
Disorder|Disease or Syndrome|Patient History|2560,2580|false|false|false|C0003873|Rheumatoid Arthritis|Rheumatoid arthritis
Disorder|Disease or Syndrome|Patient History|2571,2580|false|false|false|C0003864|Arthritis|arthritis
Finding|Functional Concept|Patient History|2591,2600|false|false|false|C0332663|Traumatic|traumatic
Anatomy|Body Location or Region|Patient History|2601,2604|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Patient History|2601,2604|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Patient History|2601,2604|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Procedure|Therapeutic or Preventive Procedure|Patient History|2607,2622|false|false|false|C0008320|Cholecystectomy procedure|Cholecystectomy
Procedure|Therapeutic or Preventive Procedure|Patient History|2625,2637|false|false|false|C0003611;C0003612|Appendectomy;Appendectomy; for ruptured appendix with abscess or generalized peritonitis|Appendectomy
Procedure|Therapeutic or Preventive Procedure|Patient History|2640,2653|false|false|false|C0040423|Tonsillectomy|Tonsillectomy
Finding|Functional Concept|Patient History|2656,2660|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|Patient History|2656,2666|false|false|false|C0230366|Structure of left wrist|Left wrist
Anatomy|Body Location or Region|Patient History|2661,2666|false|false|false|C0043262;C1322271;C4298907|Upper extremity>Wrist;Wrist;Wrist joint|wrist
Anatomy|Body Space or Junction|Patient History|2661,2666|false|false|false|C0043262;C1322271;C4298907|Upper extremity>Wrist;Wrist;Wrist joint|wrist
Procedure|Therapeutic or Preventive Procedure|Patient History|2661,2681|false|false|false|C0845620|Wrist reconstruction|wrist reconstruction
Procedure|Machine Activity|Patient History|2667,2681|false|false|false|C0020912;C0524865|Optical Image Reconstruction;Reconstructive Surgical Procedures|reconstruction
Procedure|Therapeutic or Preventive Procedure|Patient History|2667,2681|false|false|false|C0020912;C0524865|Optical Image Reconstruction;Reconstructive Surgical Procedures|reconstruction
Finding|Functional Concept|Patient History|2684,2689|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Location or Region|Patient History|2684,2702|false|false|false|C0828608|Right tendinous cuff|Right rotator cuff
Anatomy|Body Part, Organ, or Organ Component|Patient History|2690,2702|false|false|false|C0085515|Rotator Cuff|rotator cuff
Anatomy|Body Part, Organ, or Organ Component|Patient History|2698,2702|false|false|false|C1550244|Cuff - body part|cuff
Finding|Pathologic Function|Patient History|2698,2702|false|false|false|C3668885|Cuffing (morphologic abnormality)|cuff
Procedure|Machine Activity|Patient History|2703,2717|false|false|false|C0020912;C0524865|Optical Image Reconstruction;Reconstructive Surgical Procedures|reconstruction
Procedure|Therapeutic or Preventive Procedure|Patient History|2703,2717|false|false|false|C0020912;C0524865|Optical Image Reconstruction;Reconstructive Surgical Procedures|reconstruction
Finding|Finding|Family Medical History|2758,2774|false|false|false|C0424909|Family history with explicit context pertaining to father|paternal history
Finding|Conceptual Entity|Family Medical History|2767,2774|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|2767,2774|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Family Medical History|2767,2774|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|2767,2777|false|false|false|C0262926|Medical History|history of
Disorder|Neoplastic Process|Family Medical History|2790,2799|false|false|false|C0007097|Carcinoma|carcinoma
Finding|Finding|Family Medical History|2801,2809|false|false|false|C1858460|Maternal|Maternal
Finding|Finding|Family Medical History|2801,2817|false|false|false|C0559473|maternal history|Maternal history
Finding|Conceptual Entity|Family Medical History|2810,2817|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|2810,2817|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Family Medical History|2810,2817|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|2810,2820|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|Family Medical History|2821,2829|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|diabetes
Procedure|Health Care Activity|General Exam|2850,2859|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Finding|Finding|General Exam|2860,2868|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|General Exam|2860,2868|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|General Exam|2860,2868|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|General Exam|2860,2880|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAMINATION
Procedure|Health Care Activity|General Exam|2860,2880|false|false|false|C0031809|Physical Examination|PHYSICAL EXAMINATION
Event|Activity|General Exam|2869,2880|false|false|false|C4321457|Examination|EXAMINATION
Procedure|Health Care Activity|General Exam|2869,2880|false|false|false|C0031809;C0582103|Medical Examination;Physical Examination|EXAMINATION
Finding|Classification|General Exam|2961,2968|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|General Exam|2961,2968|false|false|false|C3812897|General medical service|GENERAL
Disorder|Disease or Syndrome|General Exam|2970,2975|false|false|false|C0028754|Obesity|obese
Finding|Finding|General Exam|2976,2980|false|false|false|C1706180|Male Gender|male
Finding|Intellectual Product|General Exam|2984,2988|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Finding|General Exam|2992,3000|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|General Exam|2992,3000|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Attribute|Clinical Attribute|General Exam|3001,3012|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|General Exam|3001,3012|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|General Exam|3001,3012|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|General Exam|3001,3012|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Sign or Symptom|General Exam|3001,3021|false|false|false|C0476273|Respiratory distress|respiratory distress
Finding|Finding|General Exam|3013,3021|false|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|General Exam|3013,3021|false|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|General Exam|3026,3031|false|false|false|C1512338|HEENT|HEENT
Finding|Finding|General Exam|3033,3042|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Location or Region|General Exam|3052,3062|false|false|false|C0521367|Oropharyngeal|Oropharynx
Finding|Idea or Concept|General Exam|3063,3068|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Location or Region|General Exam|3073,3077|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|General Exam|3073,3077|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|General Exam|3073,3077|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Finding|Finding|General Exam|3079,3082|false|false|false|C0428897|Jugular venous pressure|JVP
Anatomy|Body Part, Organ, or Organ Component|General Exam|3086,3096|false|false|false|C0024687|Mandible|mandibular
Anatomy|Body Part, Organ, or Organ Component|General Exam|3106,3113|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|General Exam|3106,3113|false|false|false|C1314974|Cardiac attachment|CARDIAC
Finding|Gene or Genome|General Exam|3141,3145|false|false|false|C1514917|Retinoic Acid Response Element|rare
Anatomy|Anatomical Structure|General Exam|3184,3188|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Anatomy|Body Part, Organ, or Organ Component|General Exam|3184,3188|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Finding|Intellectual Product|General Exam|3184,3188|false|false|false|C1551342|Document Body|body
Procedure|Diagnostic Procedure|General Exam|3184,3196|false|false|false|C1318474|Assessment of body build|body habitus
Anatomy|Body Location or Region|General Exam|3205,3216|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|General Exam|3205,3216|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Finding|Finding|General Exam|3205,3220|false|false|false|C0232267|Pericardial friction rub|pericardial rub
Anatomy|Body Location or Region|General Exam|3222,3233|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|Pericardial
Anatomy|Body Part, Organ, or Organ Component|General Exam|3222,3233|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|Pericardial
Drug|Substance|General Exam|3234,3239|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|General Exam|3234,3239|false|false|false|C1546604|Drain Specimen Code|drain
Finding|Body Substance|General Exam|3245,3265|false|false|false|C4518404|Serosanguinous fluid|serosanguinous fluid
Drug|Substance|General Exam|3260,3265|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|General Exam|3260,3265|false|false|false|C1546638|Fluid Specimen Code|fluid
Anatomy|Body Part, Organ, or Organ Component|General Exam|3267,3274|false|false|false|C0038293|Sternum|Sternal
Finding|Finding|General Exam|3267,3285|false|false|false|C0241246|tender sternum on palpation|Sternal tenderness
Finding|Mental Process|General Exam|3275,3285|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|General Exam|3275,3285|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Anatomy|Body Part, Organ, or Organ Component|General Exam|3289,3294|false|false|false|C0024109|Lung|LUNGS
Finding|Finding|General Exam|3311,3318|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|General Exam|3311,3318|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Finding|General Exam|3323,3332|false|false|false|C0231835|Tachypnea|tachypnea
Finding|Sign or Symptom|General Exam|3353,3361|false|false|false|C0043144|Wheezing|wheezing
Finding|Finding|General Exam|3366,3374|false|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Anatomy|Body Location or Region|General Exam|3388,3392|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|General Exam|3388,3392|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|General Exam|3388,3392|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|General Exam|3388,3392|false|false|false|C0740941|Lung Problem|lung
Anatomy|Body Location or Region|General Exam|3404,3411|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|General Exam|3404,3411|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Finding|Finding|General Exam|3404,3411|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|General Exam|3413,3418|false|false|false|C0028754|Obesity|obese
Disorder|Disease or Syndrome|General Exam|3420,3424|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Anatomy|Body Part, Organ, or Organ Component|General Exam|3439,3450|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Finding|Finding|General Exam|3452,3456|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|3452,3456|false|false|false|C0687712|warming process|Warm
Finding|Finding|General Exam|3458,3462|false|false|false|C5575035|Well (answer to question)|well
Finding|Finding|General Exam|3473,3489|false|false|false|C1720371|2+ pitting edema|2+ pitting edema
Finding|Functional Concept|General Exam|3476,3483|false|false|false|C0205323|Pitting|pitting
Finding|Finding|General Exam|3476,3489|false|false|false|C0333243|Pitting edema|pitting edema
Attribute|Clinical Attribute|General Exam|3484,3489|false|false|false|C1717255||edema
Finding|Pathologic Function|General Exam|3484,3489|false|false|false|C0013604|Edema|edema
Anatomy|Body Part, Organ, or Organ Component|General Exam|3493,3498|false|false|false|C0022742|Knee|knees
Anatomy|Body System|General Exam|3503,3507|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|General Exam|3503,3507|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|General Exam|3503,3507|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Finding|Body Substance|General Exam|3503,3507|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|General Exam|3503,3507|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|General Exam|3509,3516|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|General Exam|3509,3516|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Anatomy|Body Part, Organ, or Organ Component|General Exam|3527,3533|false|false|false|C0042449|Veins|venous
Disorder|Disease or Syndrome|General Exam|3527,3540|false|false|false|C0042344|Varicose Ulcer|venous stasis
Finding|Pathologic Function|General Exam|3527,3540|false|false|false|C4551518|Venous stasis|venous stasis
Finding|Pathologic Function|General Exam|3534,3540|false|false|false|C0333138|Stasis|stasis
Disorder|Disease or Syndrome|General Exam|3534,3551|false|false|false|C0011620|Stasis dermatitis|stasis dermatitis
Disorder|Disease or Syndrome|General Exam|3541,3551|false|false|false|C0011603|Dermatitis|dermatitis
Drug|Food|General Exam|3556,3562|false|false|false|C5890763||PULSES
Finding|Physiologic Function|General Exam|3556,3562|false|false|false|C0391850|Physiologic pulse|PULSES
Procedure|Health Care Activity|General Exam|3556,3562|false|false|false|C0034107|Pulse taking|PULSES
Attribute|Clinical Attribute|General Exam|3564,3570|false|false|false|C4522154|Distal Resection Margin|Distal
Drug|Food|General Exam|3571,3577|false|false|false|C5890763||pulses
Finding|Physiologic Function|General Exam|3571,3577|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|3571,3577|false|false|false|C0034107|Pulse taking|pulses
Finding|Conceptual Entity|General Exam|3591,3600|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|General Exam|3591,3600|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Body Substance|General Exam|3624,3633|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|3624,3633|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|3624,3633|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|3624,3633|false|false|false|C0030685|Patient Discharge|DISCHARGE
Finding|Finding|General Exam|3634,3642|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|General Exam|3634,3642|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|General Exam|3634,3642|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|General Exam|3634,3654|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAMINATION
Procedure|Health Care Activity|General Exam|3634,3654|false|false|false|C0031809|Physical Examination|PHYSICAL EXAMINATION
Event|Activity|General Exam|3643,3654|false|false|false|C4321457|Examination|EXAMINATION
Procedure|Health Care Activity|General Exam|3643,3654|false|false|false|C0031809;C0582103|Medical Examination;Physical Examination|EXAMINATION
Finding|Classification|General Exam|3692,3699|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|General Exam|3692,3699|false|false|false|C3812897|General medical service|GENERAL
Disorder|Disease or Syndrome|General Exam|3701,3706|false|false|false|C0028754|Obesity|obese
Finding|Finding|General Exam|3707,3711|false|false|false|C1706180|Male Gender|male
Finding|Intellectual Product|General Exam|3715,3719|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Finding|General Exam|3723,3731|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|General Exam|3723,3731|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Attribute|Clinical Attribute|General Exam|3732,3743|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|General Exam|3732,3743|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|General Exam|3732,3743|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|General Exam|3732,3743|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Sign or Symptom|General Exam|3732,3752|false|false|false|C0476273|Respiratory distress|respiratory distress
Finding|Finding|General Exam|3744,3752|false|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|General Exam|3744,3752|false|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|General Exam|3757,3762|false|false|false|C1512338|HEENT|HEENT
Finding|Finding|General Exam|3764,3773|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Location or Region|General Exam|3783,3793|false|false|false|C0521367|Oropharyngeal|Oropharynx
Finding|Idea or Concept|General Exam|3794,3799|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Location or Region|General Exam|3804,3808|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|General Exam|3804,3808|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|General Exam|3804,3808|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Finding|Finding|General Exam|3810,3813|true|false|false|C0428897|Jugular venous pressure|JVP
Anatomy|Body Part, Organ, or Organ Component|General Exam|3833,3840|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|General Exam|3833,3840|false|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Activity|General Exam|3849,3853|false|false|false|C0871208|Rating (action)|rate
Finding|Idea or Concept|General Exam|3849,3853|false|false|false|C1549480|Amount type - Rate|rate
Finding|Finding|General Exam|3858,3864|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|General Exam|3858,3864|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Anatomy|Anatomical Structure|General Exam|3895,3899|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Anatomy|Body Part, Organ, or Organ Component|General Exam|3895,3899|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Finding|Intellectual Product|General Exam|3895,3899|false|false|false|C1551342|Document Body|body
Procedure|Diagnostic Procedure|General Exam|3895,3907|false|false|false|C1318474|Assessment of body build|body habitus
Anatomy|Body Location or Region|General Exam|3912,3923|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|General Exam|3912,3923|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Finding|Finding|General Exam|3912,3927|true|false|false|C0232267|Pericardial friction rub|pericardial rub
Anatomy|Body Part, Organ, or Organ Component|General Exam|3943,3948|false|false|false|C0024109|Lung|LUNGS
Finding|Finding|General Exam|3950,3959|false|false|false|C0392756;C0442797|Decreasing;Reduced|Decreased
Attribute|Clinical Attribute|General Exam|3960,3971|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|General Exam|3960,3971|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|General Exam|3960,3971|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|General Exam|3960,3971|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Attribute|Clinical Attribute|General Exam|3960,3978|false|false|false|C4050166||respiratory effort
Finding|Finding|General Exam|3960,3978|false|false|false|C0425466|Respiratory effort|respiratory effort
Finding|Organism Function|General Exam|3972,3978|false|false|false|C0015264|Exertion|effort
Finding|Organism Function|General Exam|4002,4012|false|false|false|C0231800|Expiration, Respiratory|Expiratory
Finding|Sign or Symptom|General Exam|4002,4021|false|false|false|C0231875|Expiratory wheezing|Expiratory wheezing
Finding|Sign or Symptom|General Exam|4013,4021|false|false|false|C0043144|Wheezing|wheezing
Finding|Finding|General Exam|4036,4044|false|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Anatomy|Body Location or Region|General Exam|4047,4054|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|General Exam|4047,4054|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Finding|Finding|General Exam|4047,4054|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|General Exam|4056,4061|false|false|false|C0028754|Obesity|obese
Disorder|Disease or Syndrome|General Exam|4063,4067|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Anatomy|Body Part, Organ, or Organ Component|General Exam|4097,4108|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Finding|Finding|General Exam|4110,4114|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|4110,4114|false|false|false|C0687712|warming process|Warm
Finding|Finding|General Exam|4116,4120|false|false|false|C5575035|Well (answer to question)|well
Finding|Finding|General Exam|4136,4152|false|false|false|C1720371|2+ pitting edema|2+ pitting edema
Finding|Functional Concept|General Exam|4139,4146|false|false|false|C0205323|Pitting|pitting
Finding|Finding|General Exam|4139,4152|false|false|false|C0333243|Pitting edema|pitting edema
Attribute|Clinical Attribute|General Exam|4147,4152|false|false|false|C1717255||edema
Finding|Pathologic Function|General Exam|4147,4152|false|false|false|C0013604|Edema|edema
Anatomy|Body Part, Organ, or Organ Component|General Exam|4156,4161|false|false|false|C0022742|Knee|knees
Anatomy|Body System|General Exam|4166,4170|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|General Exam|4166,4170|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|General Exam|4166,4170|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Finding|Body Substance|General Exam|4166,4170|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|General Exam|4166,4170|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|General Exam|4172,4179|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|General Exam|4172,4179|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Anatomy|Body Part, Organ, or Organ Component|General Exam|4180,4186|false|false|false|C0042449|Veins|venous
Disorder|Disease or Syndrome|General Exam|4180,4193|false|false|false|C0042344|Varicose Ulcer|venous stasis
Finding|Pathologic Function|General Exam|4180,4193|false|false|false|C4551518|Venous stasis|venous stasis
Finding|Pathologic Function|General Exam|4187,4193|false|false|false|C0333138|Stasis|stasis
Disorder|Disease or Syndrome|General Exam|4187,4204|false|false|false|C0011620|Stasis dermatitis|stasis dermatitis
Disorder|Disease or Syndrome|General Exam|4194,4204|false|false|false|C0011603|Dermatitis|dermatitis
Drug|Food|General Exam|4209,4215|false|false|false|C5890763||PULSES
Finding|Physiologic Function|General Exam|4209,4215|false|false|false|C0391850|Physiologic pulse|PULSES
Procedure|Health Care Activity|General Exam|4209,4215|false|false|false|C0034107|Pulse taking|PULSES
Attribute|Clinical Attribute|General Exam|4217,4223|false|false|false|C4522154|Distal Resection Margin|Distal
Drug|Food|General Exam|4224,4230|false|false|false|C5890763||pulses
Finding|Physiologic Function|General Exam|4224,4230|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|4224,4230|false|false|false|C0034107|Pulse taking|pulses
Finding|Conceptual Entity|General Exam|4244,4253|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|General Exam|4244,4253|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Procedure|Health Care Activity|General Exam|4297,4306|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Lab|Laboratory or Test Result|General Exam|4307,4311|false|false|false|C0587081|Laboratory test finding|LABS
Anatomy|Cell|General Exam|4343,4346|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|4353,4356|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|4353,4356|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|4353,4356|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|4362,4365|false|false|false|C0019046|Hemoglobin|HGB
Drug|Biologically Active Substance|General Exam|4362,4365|false|false|false|C0019046|Hemoglobin|HGB
Finding|Gene or Genome|General Exam|4362,4365|false|false|false|C1424337|CYGB gene|HGB
Lab|Laboratory or Test Result|General Exam|4362,4365|false|false|false|C0019029|Hemoglobin concentration|HGB
Procedure|Laboratory Procedure|General Exam|4371,4374|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|General Exam|4371,4374|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Disorder|Virus|General Exam|4380,4383|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|General Exam|4380,4383|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|4380,4383|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|4380,4383|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|4388,4391|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|4388,4391|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|General Exam|4388,4391|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|4388,4391|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|4388,4391|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|4397,4401|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Finding|Body Substance|General Exam|4453,4459|false|false|false|C0024202|Lymph|LYMPHS
Drug|Antibiotic|General Exam|4465,4470|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Biomedical or Dental Material|General Exam|4465,4470|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Organic Chemical|General Exam|4465,4470|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Disorder|Disease or Syndrome|General Exam|4475,4478|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|EOS
Finding|Gene or Genome|General Exam|4475,4478|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|EOS
Disorder|Neoplastic Process|General Exam|4590,4593|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Procedure|Laboratory Procedure|General Exam|4590,4593|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Drug|Biologically Active Substance|General Exam|4617,4624|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|General Exam|4617,4624|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|General Exam|4617,4624|false|false|false|C0017725|glucose|GLUCOSE
Lab|Laboratory or Test Result|General Exam|4617,4624|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|General Exam|4617,4624|false|false|false|C0337438|Glucose measurement|GLUCOSE
Drug|Biologically Active Substance|General Exam|4630,4634|false|false|false|C0041942|urea|UREA
Drug|Organic Chemical|General Exam|4630,4634|false|false|false|C0041942|urea|UREA
Drug|Pharmacologic Substance|General Exam|4630,4634|false|false|false|C0041942|urea|UREA
Procedure|Laboratory Procedure|General Exam|4630,4634|false|false|false|C0523961|Urea measurement|UREA
Drug|Biologically Active Substance|General Exam|4650,4656|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Element, Ion, or Isotope|General Exam|4650,4656|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Pharmacologic Substance|General Exam|4650,4656|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Finding|Physiologic Function|General Exam|4650,4656|false|false|false|C4553025|Sodium metabolic function|SODIUM
Procedure|Laboratory Procedure|General Exam|4650,4656|false|false|false|C0337443|Sodium measurement|SODIUM
Drug|Biologically Active Substance|General Exam|4662,4671|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Element, Ion, or Isotope|General Exam|4662,4671|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Food|General Exam|4662,4671|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Inorganic Chemical|General Exam|4662,4671|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Pharmacologic Substance|General Exam|4662,4671|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Finding|Physiologic Function|General Exam|4662,4671|false|false|false|C4553027|Potassium metabolic function|POTASSIUM
Procedure|Laboratory Procedure|General Exam|4662,4671|false|false|false|C0202194|Potassium measurement|POTASSIUM
Drug|Element, Ion, or Isotope|General Exam|4676,4684|false|false|false|C0008203;C0596019|Chlorides;chloride ion|CHLORIDE
Finding|Physiologic Function|General Exam|4676,4684|false|false|false|C4553021|Chloride metabolic function|CHLORIDE
Procedure|Laboratory Procedure|General Exam|4676,4684|false|false|false|C0201952|Chloride measurement|CHLORIDE
Drug|Biologically Active Substance|General Exam|4695,4698|false|false|false|C0007012|carbon dioxide|CO2
Drug|Inorganic Chemical|General Exam|4695,4698|false|false|false|C0007012|carbon dioxide|CO2
Finding|Finding|General Exam|4695,4698|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Finding|Gene or Genome|General Exam|4695,4698|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Drug|Element, Ion, or Isotope|General Exam|4703,4708|false|false|false|C0003075|Anions|ANION
Attribute|Clinical Attribute|General Exam|4703,4712|false|false|false|C0003074|Anion Gap|ANION GAP
Lab|Laboratory or Test Result|General Exam|4703,4712|false|false|false|C1509129|Anion gap result|ANION GAP
Procedure|Laboratory Procedure|General Exam|4703,4712|false|false|false|C0201889;C2189246|Anion gap measurement;blood anion gap (lab test)|ANION GAP
Drug|Amino Acid, Peptide, or Protein|General Exam|4709,4712|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Drug|Biologically Active Substance|General Exam|4709,4712|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Finding|Gene or Genome|General Exam|4709,4712|false|false|false|C1419277;C2984552|RASA1 gene;RASA1 wt Allele|GAP
Drug|Biologically Active Substance|General Exam|4730,4737|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Element, Ion, or Isotope|General Exam|4730,4737|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Inorganic Chemical|General Exam|4730,4737|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Pharmacologic Substance|General Exam|4730,4737|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Vitamin|General Exam|4730,4737|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Finding|Physiologic Function|General Exam|4730,4737|false|false|false|C4553026|Calcium metabolic function|CALCIUM
Procedure|Laboratory Procedure|General Exam|4730,4737|false|false|false|C0201925|Calcium measurement|CALCIUM
Drug|Element, Ion, or Isotope|General Exam|4743,4752|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Drug|Inorganic Chemical|General Exam|4743,4752|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Drug|Pharmacologic Substance|General Exam|4743,4752|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Procedure|Laboratory Procedure|General Exam|4743,4752|false|false|false|C0523826|Phosphate measurement|PHOSPHATE
Drug|Biologically Active Substance|General Exam|4757,4766|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Element, Ion, or Isotope|General Exam|4757,4766|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Inorganic Chemical|General Exam|4757,4766|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Pharmacologic Substance|General Exam|4757,4766|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Procedure|Laboratory Procedure|General Exam|4757,4766|false|false|false|C0373675|Magnesium measurement|MAGNESIUM
Drug|Organic Chemical|General Exam|4813,4820|false|false|false|C0022924;C0376261|Lactates;lactate|LACTATE
Drug|Pharmacologic Substance|General Exam|4813,4820|false|false|false|C0022924;C0376261|Lactates;lactate|LACTATE
Procedure|Laboratory Procedure|General Exam|4813,4820|false|false|false|C0202115|Lactic acid measurement|LACTATE
Anatomy|Tissue|General Exam|4837,4844|false|false|false|C0032225|Pleura|PLEURAL
Disorder|Disease or Syndrome|General Exam|4837,4844|false|false|false|C0032226|Pleural Diseases|PLEURAL
Finding|Body Substance|General Exam|4837,4850|false|false|false|C0225778|Pleural fluid|PLEURAL FLUID
Procedure|Laboratory Procedure|General Exam|4837,4850|false|false|false|C2242629|Pleural fluid analysis|PLEURAL FLUID
Drug|Substance|General Exam|4845,4850|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|FLUID
Finding|Intellectual Product|General Exam|4845,4850|false|false|false|C1546638|Fluid Specimen Code|FLUID
Procedure|Research Activity|General Exam|4851,4858|false|false|false|C0947630|Scientific Study|STUDIES
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|4864,4869|false|false|false|C0032400;C0071360|5'-Inosinic acid, 2'-deoxy-2'-fluoro-, homopolymer;Poly A|Polys
Finding|Body Substance|General Exam|4874,4880|false|false|false|C0024202|Lymph|Lymphs
Drug|Antibiotic|General Exam|4884,4889|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|General Exam|4884,4889|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|General Exam|4884,4889|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Finding|Finding|General Exam|4894,4901|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|General Exam|4894,4901|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Procedure|Diagnostic Procedure|General Exam|4916,4919|false|false|false|C0430462|Transthoracic echocardiography|TTE
Finding|Functional Concept|General Exam|4924,4928|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|General Exam|4924,4935|false|false|false|C0225860|Left atrial structure|left atrium
Anatomy|Body Part, Organ, or Organ Component|General Exam|4929,4935|false|false|false|C0018792|Heart Atrium|atrium
Finding|Social Behavior|General Exam|4959,4967|false|false|false|C0678975|inferiority|inferior
Anatomy|Body Part, Organ, or Organ Component|General Exam|4959,4977|false|false|false|C0042458;C4266635|Abdomen>Vena cava.inferior;Inferior vena cava structure|inferior vena cava
Anatomy|Body Part, Organ, or Organ Component|General Exam|4968,4972|false|false|false|C0447122|Structure of vein of trunk|vena
Anatomy|Body Part, Organ, or Organ Component|General Exam|4968,4977|false|false|false|C0042460;C4266402|Chest+Abdomen>Vena cava.superior &or Vena cava.inferior;Vena caval structure|vena cava
Finding|Gene or Genome|General Exam|4973,4977|false|false|false|C1413046|CA5A gene|cava
Finding|Finding|General Exam|4982,4989|false|false|false|C0700124|Dilated|dilated
Finding|Functional Concept|General Exam|5017,5021|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|General Exam|5022,5033|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Space or Junction|General Exam|5063,5069|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|General Exam|5063,5069|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|General Exam|5063,5069|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|General Exam|5097,5102|false|false|false|C1846009|Intrauterine growth restriction, metaphyseal dysplasia, adrenal hypoplasia congenita, and genital anomaly syndrome|image
Finding|Intellectual Product|General Exam|5097,5102|false|false|false|C1696103;C1704254;C1704922;C3542466|Image;Image (foundation metadata concept);Medical Image;image - dosage form|image
Finding|Functional Concept|General Exam|5130,5134|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|General Exam|5135,5146|false|false|false|C0018827|Heart Ventricle|ventricular
Finding|Finding|General Exam|5147,5155|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|General Exam|5147,5155|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|General Exam|5147,5155|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|General Exam|5147,5155|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|General Exam|5157,5164|false|false|false|C0282416|Overall Publication Type|Overall
Finding|Functional Concept|General Exam|5165,5169|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|General Exam|5170,5181|false|false|false|C0018827|Heart Ventricle|ventricular
Finding|Organ or Tissue Function|General Exam|5182,5190|false|false|false|C0039155|Systole|systolic
Finding|Finding|General Exam|5191,5199|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|General Exam|5191,5199|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|General Exam|5191,5199|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|General Exam|5191,5199|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|General Exam|5233,5237|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Physiologic Function|General Exam|5233,5258|false|false|false|C2733342|Left ventricular ejection|left ventricular ejection
Anatomy|Body Part, Organ, or Organ Component|General Exam|5238,5249|false|false|false|C0018827|Heart Ventricle|ventricular
Finding|Physiologic Function|General Exam|5238,5258|false|false|false|C2733340|Ventricular ejection|ventricular ejection
Attribute|Clinical Attribute|General Exam|5250,5258|false|false|false|C0812388|Ejection time|ejection
Finding|Daily or Recreational Activity|General Exam|5250,5258|false|false|false|C0336969|Ejection as a Sports activity|ejection
Phenomenon|Phenomenon or Process|General Exam|5250,5258|false|false|false|C0302131|Ejection as a Circumstance of Injury|ejection
Finding|Intellectual Product|General Exam|5259,5267|false|false|false|C1554103|MDFAttributeType - Fraction|fraction
Finding|Functional Concept|General Exam|5277,5281|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Attribute|Clinical Attribute|General Exam|5277,5307|false|false|false|C4050538||Left ventricular cardiac index
Anatomy|Body Part, Organ, or Organ Component|General Exam|5282,5293|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Part, Organ, or Organ Component|General Exam|5294,5301|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|General Exam|5294,5301|false|false|false|C1314974|Cardiac attachment|cardiac
Finding|Finding|General Exam|5294,5307|false|false|false|C0428776|Cardiac index|cardiac index
Finding|Idea or Concept|General Exam|5302,5307|false|false|false|C0600653;C0918012;C1552854|Html Link Type - index;Index;Indexes|index
Finding|Intellectual Product|General Exam|5302,5307|false|false|false|C0600653;C0918012;C1552854|Html Link Type - index;Index;Indexes|index
Anatomy|Body Part, Organ, or Organ Component|General Exam|5339,5350|false|false|false|C0018827|Heart Ventricle|ventricular
Disorder|Congenital Abnormality|General Exam|5339,5364|true|false|false|C0018818|Ventricular Septal Defects|ventricular septal defect
Disorder|Anatomical Abnormality|General Exam|5351,5364|true|false|false|C0018816;C5779791|Congenital septal defect of heart;Heart Septal Defects|septal defect
Disorder|Congenital Abnormality|General Exam|5351,5364|true|false|false|C0018816;C5779791|Congenital septal defect of heart;Heart Septal Defects|septal defect
Disorder|Disease or Syndrome|General Exam|5358,5364|true|false|false|C1861101|THYROID HORMONE PLASMA MEMBRANE TRANSPORT DEFECT|defect
Finding|Functional Concept|General Exam|5358,5364|true|false|false|C1457869|Defect|defect
Finding|Functional Concept|General Exam|5381,5386|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Space or Junction|General Exam|5381,5405|false|false|false|C0503854|Cavity of right ventricle|right ventricular cavity
Lab|Laboratory or Test Result|General Exam|5381,5410|false|false|false|C0455865|Right ventricular cavity size|right ventricular cavity size
Anatomy|Body Part, Organ, or Organ Component|General Exam|5387,5398|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Space or Junction|General Exam|5387,5405|false|false|false|C0507083|Cavity of ventricle|ventricular cavity
Anatomy|Body Space or Junction|General Exam|5399,5405|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|General Exam|5399,5405|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|General Exam|5399,5405|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Finding|Functional Concept|General Exam|5423,5427|false|false|false|C0332296|Free of (attribute)|free
Phenomenon|Natural Phenomenon or Process|General Exam|5434,5440|false|false|false|C0026597|Motion|motion
Finding|Finding|General Exam|5451,5459|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Finding|Idea or Concept|General Exam|5451,5459|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Phenomenon|Natural Phenomenon or Process|General Exam|5484,5490|false|false|false|C0026597|Motion|motion
Anatomy|Body Part, Organ, or Organ Component|General Exam|5496,5502|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|General Exam|5496,5508|false|false|false|C0037197|Structure of sinus of Valsalva|aortic sinus
Anatomy|Body Space or Junction|General Exam|5503,5508|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|General Exam|5503,5508|false|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|General Exam|5503,5508|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|General Exam|5503,5508|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Finding|Functional Concept|General Exam|5552,5561|false|false|false|C1547175;C1962987|Ascend (action);Sequencing - Ascending|ascending
Anatomy|Body Part, Organ, or Organ Component|General Exam|5552,5567|false|false|false|C0003956|Ascending aorta structure|ascending aorta
Anatomy|Body Part, Organ, or Organ Component|General Exam|5562,5567|false|false|false|C0003483;C4037978|Aorta;Chest+Abdomen>Aorta|aorta
Procedure|Health Care Activity|General Exam|5562,5567|false|false|false|C0869784|Procedure on aorta|aorta
Finding|Finding|General Exam|5562,5576|false|false|false|C0579133|Aortic diameter|aorta diameter
Anatomy|Body Part, Organ, or Organ Component|General Exam|5593,5599|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|General Exam|5593,5604|false|false|false|C0003489;C4037976|Aortic arch structure;Chest>Aortic arch|aortic arch
Disorder|Anatomical Abnormality|General Exam|5593,5604|false|false|false|C4759703|Aortic arch malformation|aortic arch
Anatomy|Body Location or Region|General Exam|5600,5604|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Anatomy|Body Part, Organ, or Organ Component|General Exam|5600,5604|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Anatomy|Body Space or Junction|General Exam|5600,5604|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Finding|Finding|General Exam|5600,5604|false|false|false|C1538146;C4722404|Age-Related Clonal Hematopoiesis;ZBTB8OS gene|arch
Finding|Gene or Genome|General Exam|5600,5604|false|false|false|C1538146;C4722404|Age-Related Clonal Hematopoiesis;ZBTB8OS gene|arch
Finding|Idea or Concept|General Exam|5637,5645|true|false|false|C3887511|Evidence|evidence
Anatomy|Body Part, Organ, or Organ Component|General Exam|5654,5660|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|General Exam|5654,5665|false|false|false|C0003489;C4037976|Aortic arch structure;Chest>Aortic arch|aortic arch
Disorder|Anatomical Abnormality|General Exam|5654,5665|false|false|false|C4759703|Aortic arch malformation|aortic arch
Anatomy|Body Location or Region|General Exam|5661,5665|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Anatomy|Body Part, Organ, or Organ Component|General Exam|5661,5665|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Anatomy|Body Space or Junction|General Exam|5661,5665|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Finding|Finding|General Exam|5661,5665|false|false|false|C1538146;C4722404|Age-Related Clonal Hematopoiesis;ZBTB8OS gene|arch
Finding|Gene or Genome|General Exam|5661,5665|false|false|false|C1538146;C4722404|Age-Related Clonal Hematopoiesis;ZBTB8OS gene|arch
Disorder|Anatomical Abnormality|General Exam|5666,5677|false|false|false|C0003492;C0332886|Aortic coarctation;Coarctation|coarctation
Disorder|Congenital Abnormality|General Exam|5666,5677|false|false|false|C0003492;C0332886|Aortic coarctation;Coarctation|coarctation
Anatomy|Body Part, Organ, or Organ Component|General Exam|5683,5689|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|General Exam|5690,5695|false|false|false|C1186983|Anatomical valve|valve
Anatomy|Body Part, Organ, or Organ Component|General Exam|5751,5757|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|General Exam|5751,5763|false|false|false|C0003501;C4533215|Aortic valve structure;Chest>Aortic valve|aortic valve
Disorder|Congenital Abnormality|General Exam|5751,5772|false|false|false|C5193127;C5700069|AORTIC VALVE DISEASE 3;Stenosis of aorta|aortic valve stenosis
Disorder|Disease or Syndrome|General Exam|5751,5772|false|false|false|C5193127;C5700069|AORTIC VALVE DISEASE 3;Stenosis of aorta|aortic valve stenosis
Finding|Pathologic Function|General Exam|5751,5772|false|false|false|C0003507|Aortic Valve Stenosis|aortic valve stenosis
Anatomy|Body Part, Organ, or Organ Component|General Exam|5758,5763|false|false|false|C1186983|Anatomical valve|valve
Finding|Pathologic Function|General Exam|5764,5772|false|false|false|C1261287|Stenosis|stenosis
Anatomy|Body Part, Organ, or Organ Component|General Exam|5786,5792|false|false|false|C0003483|Aorta|aortic
Finding|Finding|General Exam|5793,5806|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|General Exam|5793,5806|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|General Exam|5793,5806|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Anatomy|Body Part, Organ, or Organ Component|General Exam|5812,5824|false|false|false|C0026264|Mitral Valve|mitral valve
Anatomy|Body Part, Organ, or Organ Component|General Exam|5819,5824|false|false|false|C1186983|Anatomical valve|valve
Finding|Finding|General Exam|5832,5836|true|false|false|C5575035|Well (answer to question)|well
Anatomy|Body Part, Organ, or Organ Component|General Exam|5854,5869|true|false|false|C0040960|Tricuspid valve structure|tricuspid valve
Anatomy|Body Part, Organ, or Organ Component|General Exam|5864,5869|false|false|false|C1186983|Anatomical valve|valve
Finding|Finding|General Exam|5877,5881|true|false|false|C5575035|Well (answer to question)|well
Anatomy|Body Part, Organ, or Organ Component|General Exam|5892,5901|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|General Exam|5892,5901|false|false|false|C2707265||pulmonary
Finding|Finding|General Exam|5892,5901|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Anatomy|Body Part, Organ, or Organ Component|General Exam|5902,5908|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|General Exam|5902,5908|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Finding|Organ or Tissue Function|General Exam|5909,5917|false|false|false|C0039155|Systole|systolic
Attribute|Clinical Attribute|General Exam|5909,5926|false|false|false|C0871470|Systolic Pressure|systolic pressure
Finding|Finding|General Exam|5918,5926|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|General Exam|5918,5926|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|General Exam|5918,5926|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|General Exam|5918,5926|false|false|false|C0033095||pressure
Anatomy|Body Location or Region|General Exam|5964,5975|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|General Exam|5964,5975|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Disorder|Disease or Syndrome|General Exam|5964,5984|false|false|false|C0031039|Pericardial effusion|pericardial effusion
Finding|Body Substance|General Exam|5964,5984|false|false|false|C1253937|Pericardial effusion body substance|pericardial effusion
Finding|Body Substance|General Exam|5976,5984|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|General Exam|5976,5984|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|General Exam|5976,5984|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Conceptual Entity|General Exam|5987,5992|false|false|false|C3811161;C4049106|Micro (prefix);Microbiology - Laboratory Class|MICRO
Finding|Intellectual Product|General Exam|5987,5992|false|false|false|C3811161;C4049106|Micro (prefix);Microbiology - Laboratory Class|MICRO
Procedure|Laboratory Procedure|General Exam|5987,5992|false|false|false|C0085672|Microbiology procedure|MICRO
Drug|Substance|General Exam|6013,6018|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|FLUID
Finding|Intellectual Product|General Exam|6013,6018|false|false|false|C1546638|Fluid Specimen Code|FLUID
Finding|Intellectual Product|General Exam|6013,6024|false|false|false|C1546636|Fluid, Other|FLUID,OTHER
Anatomy|Body Location or Region|General Exam|6030,6041|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|PERICARDIAL
Anatomy|Body Part, Organ, or Organ Component|General Exam|6030,6041|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|PERICARDIAL
Disorder|Disease or Syndrome|General Exam|6030,6047|false|false|false|C0031039|Pericardial effusion|PERICARDIAL FLUID
Finding|Body Substance|General Exam|6030,6047|false|false|false|C0225973|Pericardial fluid (substance)|PERICARDIAL FLUID
Procedure|Laboratory Procedure|General Exam|6030,6047|false|false|false|C3854061|pericardial fluid analysis|PERICARDIAL FLUID
Drug|Substance|General Exam|6042,6047|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|FLUID
Finding|Intellectual Product|General Exam|6042,6047|false|false|false|C1546638|Fluid Specimen Code|FLUID
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|6054,6064|false|false|false|C0061856|Gram's stain|GRAM STAIN
Drug|Organic Chemical|General Exam|6054,6064|false|false|false|C0061856|Gram's stain|GRAM STAIN
Procedure|Laboratory Procedure|General Exam|6054,6064|false|false|false|C0200966|Bacterial stain, routine|GRAM STAIN
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|6059,6064|false|false|false|C0038128|Stains|STAIN
Procedure|Laboratory Procedure|General Exam|6059,6064|false|false|false|C0487602|Staining method|STAIN
Finding|Idea or Concept|General Exam|6066,6071|false|false|false|C1546485|Diagnosis Type - Final|Final
Finding|Conceptual Entity|General Exam|6104,6109|false|false|false|C1521738;C2346620;C2349184|Field;Force Field;Knowledge Field|FIELD
Procedure|Health Care Activity|General Exam|6104,6109|false|false|false|C1553496|field - patient encounter|FIELD
Anatomy|Cell|General Exam|6133,6143|false|false|false|C0023516|Leukocytes|LEUKOCYTES
Finding|Body Substance|General Exam|6133,6143|false|false|false|C1547962;C1550647|Specimen Type - Leukocytes|LEUKOCYTES
Finding|Intellectual Product|General Exam|6133,6143|false|false|false|C1547962;C1550647|Specimen Type - Leukocytes|LEUKOCYTES
Finding|Finding|General Exam|6155,6174|false|false|false|C2924473|Microorganisms seen|MICROORGANISMS SEEN
Event|Activity|General Exam|6206,6211|false|false|false|C1947932|Smear - instruction imperative|smear
Finding|Functional Concept|General Exam|6206,6211|false|false|false|C3872789|Smearing technique|smear
Procedure|Diagnostic Procedure|General Exam|6206,6211|false|false|false|C0444186|Smear test|smear
Finding|Functional Concept|General Exam|6229,6235|false|false|false|C0025663;C0449851;C2828387|Method, LOINC Axis 6;Methods;Techniques|method
Finding|Intellectual Product|General Exam|6229,6235|false|false|false|C0025663;C0449851;C2828387|Method, LOINC Axis 6;Methods;Techniques|method
Finding|Intellectual Product|General Exam|6260,6270|false|false|false|C1547985|Diagnostic Service Section ID - Hematology|hematology
Procedure|Laboratory Procedure|General Exam|6260,6270|false|false|false|C0018941;C0200627;C2183233|Hematologic Tests;Hematology procedure;diagnostic service sources hematology (procedure)|hematology
Anatomy|Cell|General Exam|6290,6306|false|false|false|C0023516|Leukocytes|white blood cell
Lab|Laboratory or Test Result|General Exam|6290,6312|false|false|false|C0427512||white blood cell count
Procedure|Laboratory Procedure|General Exam|6290,6312|false|false|false|C0023508|White Blood Cell Count procedure|white blood cell count
Disorder|Disease or Syndrome|General Exam|6296,6301|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|General Exam|6296,6301|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Anatomy|Cell|General Exam|6296,6306|false|false|false|C0005773|Blood Cells|blood cell
Procedure|Laboratory Procedure|General Exam|6296,6312|false|false|false|C0005771;C0009555|Blood Cell Count;Complete Blood Count|blood cell count
Anatomy|Cell|General Exam|6302,6306|false|false|false|C0007634|Cells|cell
Finding|Gene or Genome|General Exam|6302,6306|false|false|false|C1413336;C1413337|CEL gene;CELP gene|cell
Procedure|Laboratory Procedure|General Exam|6302,6312|false|false|false|C0007584|Cell Count|cell count
Drug|Substance|General Exam|6320,6325|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|FLUID
Finding|Intellectual Product|General Exam|6320,6325|false|false|false|C1546638|Fluid Specimen Code|FLUID
Drug|Biomedical or Dental Material|General Exam|6326,6333|false|false|false|C1706355|Culture Dose Form|CULTURE
Finding|Functional Concept|General Exam|6326,6333|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|General Exam|6326,6333|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|General Exam|6326,6333|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Disorder|Disease or Syndrome|General Exam|6409,6423|false|false|false|C0374989|Unspecified Staphylococcus infection in conditions classified elsewhere and of unspecified site|STAPHYLOCOCCUS
Drug|Amino Acid, Peptide, or Protein|General Exam|6425,6434|false|false|false|C0009118|Coagulase|COAGULASE
Drug|Enzyme|General Exam|6425,6434|false|false|false|C0009118|Coagulase|COAGULASE
Anatomy|Cell|General Exam|6450,6456|false|false|false|C1947989|Colony (cells or organisms)|COLONY
Procedure|Laboratory Procedure|General Exam|6475,6492|false|false|false|C1273935|Anaerobic microbial culture|ANAEROBIC CULTURE
Drug|Biomedical or Dental Material|General Exam|6485,6492|false|false|false|C1706355|Culture Dose Form|CULTURE
Finding|Functional Concept|General Exam|6485,6492|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|General Exam|6485,6492|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|General Exam|6485,6492|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Finding|Functional Concept|General Exam|6539,6545|false|false|false|C0521033|Fungal|FUNGAL
Procedure|Laboratory Procedure|General Exam|6539,6553|false|false|false|C0200954|Mycology culture|FUNGAL CULTURE
Drug|Biomedical or Dental Material|General Exam|6546,6553|false|false|false|C1706355|Culture Dose Form|CULTURE
Finding|Functional Concept|General Exam|6546,6553|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|General Exam|6546,6553|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|General Exam|6546,6553|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|6574,6583|false|false|false|C1318720|Acid fast stain|ACID FAST
Finding|Finding|General Exam|6579,6583|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Finding|Gene or Genome|General Exam|6579,6583|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Finding|Molecular Function|General Exam|6579,6583|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Event|Activity|General Exam|6584,6589|false|false|false|C1947932|Smear - instruction imperative|SMEAR
Finding|Functional Concept|General Exam|6584,6589|false|false|false|C3872789|Smearing technique|SMEAR
Procedure|Diagnostic Procedure|General Exam|6584,6589|false|false|false|C0444186|Smear test|SMEAR
Finding|Idea or Concept|General Exam|6591,6596|false|false|false|C1546485|Diagnosis Type - Final|Final
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|6612,6621|true|false|false|C1318720|Acid fast stain|ACID FAST
Finding|Finding|General Exam|6617,6621|true|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Finding|Gene or Genome|General Exam|6617,6621|true|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Finding|Molecular Function|General Exam|6617,6621|true|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Finding|Intellectual Product|General Exam|6638,6644|false|false|false|C1552596;C3244286|Direct - PostalAddressUse;direct address|DIRECT
Event|Activity|General Exam|6645,6650|false|false|false|C1947932|Smear - instruction imperative|SMEAR
Finding|Functional Concept|General Exam|6645,6650|false|false|false|C3872789|Smearing technique|SMEAR
Procedure|Diagnostic Procedure|General Exam|6645,6650|false|false|false|C0444186|Smear test|SMEAR
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|6657,6666|false|false|false|C1318720|Acid fast stain|ACID FAST
Finding|Finding|General Exam|6662,6666|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Finding|Gene or Genome|General Exam|6662,6666|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Finding|Molecular Function|General Exam|6662,6666|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|FAST
Drug|Biomedical or Dental Material|General Exam|6667,6674|false|false|false|C1706355|Culture Dose Form|CULTURE
Finding|Functional Concept|General Exam|6667,6674|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|General Exam|6667,6674|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|General Exam|6667,6674|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Finding|Body Substance|General Exam|6692,6701|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|6692,6701|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|6692,6701|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|6692,6701|false|false|false|C0030685|Patient Discharge|DISCHARGE
Lab|Laboratory or Test Result|General Exam|6702,6706|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|General Exam|6736,6741|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|6736,6741|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|6742,6745|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|6752,6755|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|6752,6755|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|6752,6755|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|6762,6765|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|6762,6765|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|6762,6765|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|6762,6765|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|6772,6775|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|6772,6775|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|6783,6786|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|General Exam|6783,6786|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|6783,6786|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|6783,6786|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|6790,6793|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|6790,6793|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|General Exam|6790,6793|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|6790,6793|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|6790,6793|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|6799,6803|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|6829,6832|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|6849,6854|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|6849,6854|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|6849,6862|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|6849,6862|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|6849,6862|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|6855,6862|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|6855,6862|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|6855,6862|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|General Exam|6855,6862|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|6855,6862|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|6909,6913|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|6909,6913|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|6909,6913|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|6938,6943|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|6938,6943|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|6944,6947|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|6944,6947|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|General Exam|6944,6947|false|false|false|C0001899|Alanine Transaminase|ALT
Finding|Gene or Genome|General Exam|6944,6947|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|General Exam|6944,6947|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|General Exam|6944,6947|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|General Exam|6944,6947|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|General Exam|6952,6955|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|General Exam|6952,6955|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|6952,6955|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|General Exam|6952,6955|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|General Exam|6952,6955|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Finding|Gene or Genome|General Exam|6952,6955|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|6959,6966|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|General Exam|6959,6966|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|General Exam|6994,6999|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|6994,6999|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|6994,7007|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|General Exam|7000,7007|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|7000,7007|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|7000,7007|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|7000,7007|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|7000,7007|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Finding|Physiologic Function|General Exam|7000,7007|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|7000,7007|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|General Exam|7041,7046|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|7041,7046|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|7047,7053|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Drug|Hormone|General Exam|7047,7053|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Disorder|Disease or Syndrome|General Exam|7070,7075|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|7070,7075|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Attribute|Clinical Attribute|General Exam|7076,7079|false|false|false|C2708739||TSH
Drug|Amino Acid, Peptide, or Protein|General Exam|7076,7079|false|false|false|C0040160|thyrotropin|TSH
Drug|Hormone|General Exam|7076,7079|false|false|false|C0040160|thyrotropin|TSH
Drug|Pharmacologic Substance|General Exam|7076,7079|false|false|false|C0040160|thyrotropin|TSH
Procedure|Laboratory Procedure|General Exam|7076,7079|false|false|false|C0202230|Thyroid stimulating hormone measurement|TSH
Disorder|Disease or Syndrome|General Exam|7097,7102|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|7097,7102|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Classification|General Exam|7107,7110|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|pO2
Finding|Molecular Function|General Exam|7107,7110|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|pO2
Procedure|Laboratory Procedure|General Exam|7107,7110|false|false|false|C1283004|PO2 measurement|pO2
Lab|Laboratory or Test Result|General Exam|7115,7119|false|false|false|C0391839|Carbon dioxide, partial pressure|pCO2
Procedure|Laboratory Procedure|General Exam|7115,7119|false|false|false|C0201931|Carbon dioxide measurement, partial pressure|pCO2
Anatomy|Body Location or Region|General Exam|7144,7148|false|false|false|C2987514|Anatomical base|Base
Drug|Biomedical or Dental Material|General Exam|7144,7148|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Drug|Chemical Viewed Functionally|General Exam|7144,7148|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|7144,7148|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Finding|Gene or Genome|General Exam|7144,7148|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|Base
Finding|Idea or Concept|General Exam|7144,7148|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|Base
Finding|Intellectual Product|Hospital Course|7180,7187|false|false|false|C1552616;C1706244|Summary (document);summary - ActRelationshipSubset|SUMMARY
Finding|Finding|Hospital Course|7217,7221|false|false|false|C1706180|Male Gender|male
Disorder|Disease or Syndrome|Hospital Course|7227,7247|false|false|false|C0003873|Rheumatoid Arthritis|rheumatoid arthritis
Disorder|Disease or Syndrome|Hospital Course|7238,7247|false|false|false|C0003864|Arthritis|arthritis
Drug|Pharmacologic Substance|Hospital Course|7249,7254|false|false|false|C0242708|Antirheumatic Drugs, Disease-Modifying|DMARD
Event|Event|Hospital Course|7255,7262|false|false|false|C0019843|Holidays|holiday
Finding|Intellectual Product|Hospital Course|7276,7281|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|brief
Procedure|Health Care Activity|Hospital Course|7282,7297|false|false|false|C0019993|Hospitalization|hospitalization
Disorder|Disease or Syndrome|Hospital Course|7314,7326|false|false|false|C0031046|Pericarditis|pericarditis
Finding|Idea or Concept|Hospital Course|7348,7356|false|false|false|C1547192|Organization unit type - Hospital|hospital
Anatomy|Body Location or Region|Hospital Course|7362,7373|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7362,7373|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Disorder|Disease or Syndrome|Hospital Course|7362,7382|false|false|false|C0031039|Pericardial effusion|pericardial effusion
Finding|Body Substance|Hospital Course|7362,7382|false|false|false|C1253937|Pericardial effusion body substance|pericardial effusion
Finding|Body Substance|Hospital Course|7374,7382|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|Hospital Course|7374,7382|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|Hospital Course|7374,7382|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Finding|Hospital Course|7389,7397|false|false|false|C0332149|Possible|possible
Finding|Functional Concept|Hospital Course|7398,7407|false|true|false|C0332459|Compressed structure|tamponade
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7398,7407|false|true|false|C0579016||tamponade
Finding|Physiologic Function|Hospital Course|7408,7418|false|true|false|C0031843|physiological aspects|physiology
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7437,7455|false|false|false|C0191234|Pericardiocentesis|pericardiocentesis
Finding|Functional Concept|Hospital Course|7465,7473|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|Hospital Course|7465,7473|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|Hospital Course|7465,7473|false|false|false|C4706767|Transfer (immobility management)|transfer
Anatomy|Body Location or Region|Hospital Course|7492,7503|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7492,7503|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Disorder|Disease or Syndrome|Hospital Course|7492,7512|false|false|false|C0031039|Pericardial effusion|pericardial effusion
Finding|Body Substance|Hospital Course|7492,7512|false|false|false|C1253937|Pericardial effusion body substance|pericardial effusion
Finding|Body Substance|Hospital Course|7504,7512|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|Hospital Course|7504,7512|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|Hospital Course|7504,7512|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Drug|Substance|Hospital Course|7521,7526|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|Hospital Course|7521,7526|false|false|false|C1546604|Drain Specimen Code|drain
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7521,7536|false|false|false|C3495845|Drain placement|drain placement
Procedure|Health Care Activity|Hospital Course|7527,7536|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7527,7536|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Finding|Intellectual Product|Hospital Course|7565,7570|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Attribute|Clinical Attribute|Hospital Course|7584,7595|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|Hospital Course|7584,7595|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|Hospital Course|7584,7595|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|Hospital Course|7584,7595|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Sign or Symptom|Hospital Course|7584,7604|false|false|false|C0476273|Respiratory distress|respiratory distress
Finding|Finding|Hospital Course|7596,7604|false|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|Hospital Course|7596,7604|false|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7621,7628|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Immunologic Factor|Hospital Course|7621,7628|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Pharmacologic Substance|Hospital Course|7621,7628|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Finding|Finding|Hospital Course|7621,7628|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Functional Concept|Hospital Course|7621,7628|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Idea or Concept|Hospital Course|7621,7628|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Intellectual Product|Hospital Course|7621,7628|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Molecular Function|Hospital Course|7631,7635|false|false|false|C1150186|matrix metalloproteinase 7 activity|PUMP
Finding|Finding|Hospital Course|7672,7680|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|Hospital Course|7672,7680|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|Hospital Course|7672,7680|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|Hospital Course|7672,7680|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Finding|Hospital Course|7684,7690|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|RHYTHM
Finding|Physiologic Function|Hospital Course|7684,7690|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|RHYTHM
Finding|Molecular Function|Hospital Course|7692,7695|false|false|false|C1704493;C2700623|Neutral Sidebent Rotated|NSR
Finding|Pathologic Function|Hospital Course|7692,7695|false|false|false|C1704493;C2700623|Neutral Sidebent Rotated|NSR
Disorder|Disease or Syndrome|Hospital Course|7697,7700|false|false|false|C0235480;C0393911|Paroxysmal atrial fibrillation;Pure Autonomic Failure|pAF
Drug|Immunologic Factor|Hospital Course|7697,7700|false|false|false|C0032172|Platelet Activating Factor|pAF
Drug|Organic Chemical|Hospital Course|7697,7700|false|false|false|C0032172|Platelet Activating Factor|pAF
Finding|Gene or Genome|Hospital Course|7697,7700|false|false|false|C1537443|PCLAF gene|pAF
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7697,7700|false|false|false|C0279389|doxorubicin/fluorouracil/melphalan protocol|pAF
Finding|Idea or Concept|Hospital Course|7706,7718|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Drug|Organic Chemical|Hospital Course|7772,7781|false|false|false|C0020740|ibuprofen|ibuprofen
Drug|Pharmacologic Substance|Hospital Course|7772,7781|false|false|false|C0020740|ibuprofen|ibuprofen
Drug|Organic Chemical|Hospital Course|7796,7806|false|false|false|C0009262|colchicine|colchicine
Drug|Pharmacologic Substance|Hospital Course|7796,7806|false|false|false|C0009262|colchicine|colchicine
Disorder|Mental or Behavioral Dysfunction|Hospital Course|7814,7817|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7814,7817|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|7814,7817|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|7814,7817|false|false|false|C1332410|BID gene|BID
Finding|Functional Concept|Hospital Course|7826,7838|false|false|false|C0333348|Inflammatory|inflammatory
Disorder|Disease or Syndrome|Hospital Course|7839,7851|false|false|false|C0031046|Pericarditis|pericarditis
Drug|Organic Chemical|Hospital Course|7873,7883|false|false|false|C0009262|colchicine|colchicine
Drug|Pharmacologic Substance|Hospital Course|7873,7883|false|false|false|C0009262|colchicine|colchicine
Drug|Organic Chemical|Hospital Course|7917,7926|false|false|false|C0020740|ibuprofen|ibuprofen
Drug|Pharmacologic Substance|Hospital Course|7917,7926|false|false|false|C0020740|ibuprofen|ibuprofen
Finding|Conceptual Entity|Hospital Course|7953,7963|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolution
Finding|Pathologic Function|Hospital Course|7953,7963|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolution
Finding|Functional Concept|Hospital Course|7971,7979|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Hospital Course|7971,7979|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Idea or Concept|Hospital Course|8008,8012|false|false|false|C0035647|Risk|risk
Finding|Idea or Concept|Hospital Course|8008,8015|false|false|false|C0035647|Risk|risk of
Disorder|Neoplastic Process|Hospital Course|8016,8026|false|false|false|C1458156|Recurrent Malignant Neoplasm|recurrence
Finding|Pathologic Function|Hospital Course|8016,8026|false|false|false|C2825055|Recurrence (disease attribute)|recurrence
Phenomenon|Phenomenon or Process|Hospital Course|8016,8026|false|false|false|C0034897|Recurrence|recurrence
Drug|Pharmacologic Substance|Hospital Course|8055,8058|false|false|false|C0358591|Proton Pump Inhibitors|PPI
Finding|Physiologic Function|Hospital Course|8055,8058|false|false|false|C0871125|Prepulse Inhibition|PPI
Drug|Organic Chemical|Hospital Course|8094,8103|false|false|false|C0020740|ibuprofen|ibuprofen
Drug|Pharmacologic Substance|Hospital Course|8094,8103|false|false|false|C0020740|ibuprofen|ibuprofen
Finding|Body Substance|Hospital Course|8133,8140|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|8133,8140|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|8133,8140|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Classification|Hospital Course|8149,8159|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|8149,8159|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Finding|Hospital Course|8172,8176|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|Hospital Course|8172,8176|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|Hospital Course|8172,8176|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Mental Process|Hospital Course|8177,8186|false|false|false|C0242114|Suspicion|suspicion
Drug|Biomedical or Dental Material|Hospital Course|8191,8199|false|false|false|C0168634|BaseLine dental cement|baseline
Finding|Idea or Concept|Hospital Course|8191,8199|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Functional Concept|Hospital Course|8200,8211|false|false|false|C0549186|Obstructed|obstructive
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8224,8233|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Hospital Course|8224,8233|false|false|false|C2707265||pulmonary
Finding|Finding|Hospital Course|8224,8233|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Disorder|Disease or Syndrome|Hospital Course|8235,8242|false|false|false|C0012634|Disease|disease
Finding|Body Substance|Hospital Course|8247,8254|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|8247,8254|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|8247,8254|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Disorder|Disease or Syndrome|Hospital Course|8276,8280|false|false|false|C0004238|Atrial Fibrillation|afib
Lab|Laboratory or Test Result|Hospital Course|8276,8280|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|afib
Finding|Finding|Hospital Course|8286,8289|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Finding|Gene or Genome|Hospital Course|8286,8289|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Procedure|Health Care Activity|Hospital Course|8303,8312|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Finding|Hospital Course|8324,8327|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Hospital Course|8324,8327|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Finding|Hospital Course|8324,8337|false|false|false|C2585997|New diagnosis (finding)|new diagnosis
Procedure|Diagnostic Procedure|Hospital Course|8324,8337|false|false|false|C1882082|New Diagnosis Procedure|new diagnosis
Attribute|Clinical Attribute|Hospital Course|8328,8337|false|false|false|C0945731||diagnosis
Finding|Classification|Hospital Course|8328,8337|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|Hospital Course|8328,8337|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|Hospital Course|8328,8337|false|false|false|C0011900|Diagnosis|diagnosis
Disorder|Disease or Syndrome|Hospital Course|8355,8367|false|false|false|C0020538|Hypertensive disease|hypertension
Disorder|Disease or Syndrome|Hospital Course|8373,8381|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|diabetes
Finding|Finding|Hospital Course|8383,8398|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|Anticoagulation
Finding|Physiologic Function|Hospital Course|8383,8398|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|Anticoagulation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8383,8398|false|false|false|C0003281|Anticoagulation Therapy|Anticoagulation
Procedure|Health Care Activity|Hospital Course|8428,8437|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Finding|Hospital Course|8480,8483|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Hospital Course|8480,8483|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Finding|Hospital Course|8480,8488|false|false|false|C5201228;C5202762|International Prognostic Index Low Risk Group;Low risk|low risk
Finding|Idea or Concept|Hospital Course|8484,8488|false|false|false|C0035647|Risk|risk
Disorder|Disease or Syndrome|Hospital Course|8494,8497|false|false|false|C0001365;C0038454|Acute ill-defined cerebrovascular disease;Cerebrovascular accident|CVA
Drug|Pharmacologic Substance|Hospital Course|8494,8497|false|false|false|C5779650|Cyclophosphamide/Doxorubicin/Vincristine|CVA
Finding|Finding|Hospital Course|8534,8537|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Hospital Course|8534,8537|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Finding|Hospital Course|8534,8547|false|false|false|C2585997|New diagnosis (finding)|new diagnosis
Procedure|Diagnostic Procedure|Hospital Course|8534,8547|false|false|false|C1882082|New Diagnosis Procedure|new diagnosis
Attribute|Clinical Attribute|Hospital Course|8538,8547|false|false|false|C0945731||diagnosis
Finding|Classification|Hospital Course|8538,8547|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|Hospital Course|8538,8547|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|Hospital Course|8538,8547|false|false|false|C0011900|Diagnosis|diagnosis
Finding|Functional Concept|Hospital Course|8562,8566|false|false|false|C0686904|Patient need for (contextual qualifier)|need
Finding|Functional Concept|Hospital Course|8562,8570|false|false|false|C0686904|Patient need for (contextual qualifier)|need for
Finding|Finding|Hospital Course|8571,8586|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|Hospital Course|8571,8586|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8571,8586|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Finding|Idea or Concept|Hospital Course|8624,8629|false|false|false|C0750546|newly|newly
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8649,8654|false|false|false|C0019018|Glycosylated hemoglobin A|HbA1c
Drug|Biologically Active Substance|Hospital Course|8649,8654|false|false|false|C0019018|Glycosylated hemoglobin A|HbA1c
Procedure|Laboratory Procedure|Hospital Course|8649,8654|false|false|false|C0202054|Glucohemoglobin measurement|HbA1c
Drug|Organic Chemical|Hospital Course|8693,8702|false|false|false|C0025598|metformin|metformin
Drug|Pharmacologic Substance|Hospital Course|8693,8702|false|false|false|C0025598|metformin|metformin
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8707,8710|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8707,8710|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8707,8710|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|8707,8710|false|false|false|C1332410|BID gene|BID
Finding|Classification|Hospital Course|8726,8736|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|8726,8736|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Functional Concept|Hospital Course|8737,8743|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|Hospital Course|8737,8743|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|Hospital Course|8737,8746|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|Hospital Course|8737,8746|false|false|false|C1522577|follow-up|follow-up
Finding|Classification|Hospital Course|8793,8803|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|8793,8803|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Mental Process|Hospital Course|8804,8811|false|false|false|C0542559|contextual factors|setting
Drug|Pharmacologic Substance|Hospital Course|8842,8850|false|false|false|C0012798;C5399719|Diuretic [APC];Diuretics|diuretic
Finding|Classification|Hospital Course|8858,8868|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|8858,8868|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Mental Process|Hospital Course|8869,8876|false|false|false|C0542559|contextual factors|setting
Finding|Idea or Concept|Hospital Course|8907,8915|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Hospital Course|8907,8918|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8919,8924|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Hospital Course|8919,8924|true|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Hospital Course|8919,8924|true|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|Hospital Course|8919,8932|true|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Finding|Functional Concept|Hospital Course|8925,8932|true|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|Hospital Course|8925,8932|true|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|Hospital Course|8925,8932|true|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Procedure|Health Care Activity|Hospital Course|8946,8955|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Drug|Pharmacologic Substance|Hospital Course|8981,8990|false|false|false|C0012798|Diuretics|diuretics
Finding|Finding|Hospital Course|8994,8997|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Finding|Idea or Concept|Hospital Course|8994,8997|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Drug|Pharmacologic Substance|Hospital Course|8994,9009|false|false|false|C1718097|New medications|New medications
Attribute|Clinical Attribute|Hospital Course|8998,9009|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Hospital Course|8998,9009|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|Hospital Course|8998,9009|false|false|false|C4284232|Medications|medications
Drug|Organic Chemical|Hospital Course|9011,9020|false|false|false|C0025598|metformin|Metformin
Drug|Pharmacologic Substance|Hospital Course|9011,9020|false|false|false|C0025598|metformin|Metformin
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9027,9030|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9027,9030|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9027,9030|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|9027,9030|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|9031,9041|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|Hospital Course|9031,9041|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|Hospital Course|9054,9064|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Pharmacologic Substance|Hospital Course|9054,9064|false|false|false|C0028978|omeprazole|Omeprazole
Attribute|Clinical Attribute|Hospital Course|9085,9096|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Hospital Course|9085,9096|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|Hospital Course|9085,9096|false|false|false|C4284232|Medications|medications
Drug|Organic Chemical|Hospital Course|9098,9110|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|9098,9110|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|Hospital Course|9120,9130|false|false|false|C0009262|colchicine|Colchicine
Drug|Pharmacologic Substance|Hospital Course|9120,9130|false|false|false|C0009262|colchicine|Colchicine
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9137,9140|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9137,9140|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9137,9140|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|9137,9140|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|9141,9150|false|false|false|C0020740|ibuprofen|Ibuprofen
Drug|Pharmacologic Substance|Hospital Course|9141,9150|false|false|false|C0020740|ibuprofen|Ibuprofen
Drug|Organic Chemical|Hospital Course|9161,9171|false|false|false|C0016410|folic acid|Folic acid
Drug|Pharmacologic Substance|Hospital Course|9161,9171|false|false|false|C0016410|folic acid|Folic acid
Drug|Vitamin|Hospital Course|9161,9171|false|false|false|C0016410|folic acid|Folic acid
Procedure|Laboratory Procedure|Hospital Course|9161,9171|false|false|false|C0523631|Folic acid measurement|Folic acid
Drug|Organic Chemical|Hospital Course|9182,9192|false|false|false|C0074393|sertraline|Sertraline
Drug|Pharmacologic Substance|Hospital Course|9182,9192|false|false|false|C0074393|sertraline|Sertraline
Attribute|Clinical Attribute|Hospital Course|9214,9225|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Hospital Course|9214,9225|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|Hospital Course|9214,9225|false|false|false|C4284232|Medications|medications
Drug|Organic Chemical|Hospital Course|9228,9240|false|false|false|C0025677|methotrexate|Methotrexate
Drug|Pharmacologic Substance|Hospital Course|9228,9240|false|false|false|C0025677|methotrexate|Methotrexate
Procedure|Laboratory Procedure|Hospital Course|9228,9240|false|false|false|C5399953|Drug assay methotrexate|Methotrexate
Drug|Organic Chemical|Hospital Course|9249,9259|false|false|false|C0015620|famotidine|Famotidine
Drug|Pharmacologic Substance|Hospital Course|9249,9259|false|false|false|C0015620|famotidine|Famotidine
Finding|Intellectual Product|Hospital Course|9269,9274|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|ACUTE
Finding|Intellectual Product|Hospital Course|9301,9306|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Disorder|Disease or Syndrome|Hospital Course|9301,9319|false|false|false|C0155679|Acute pericarditis|Acute pericarditis
Disorder|Disease or Syndrome|Hospital Course|9307,9319|false|false|false|C0031046|Pericarditis|pericarditis
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9323,9330|false|false|false|C0018787|Heart|Cardiac
Finding|Intellectual Product|Hospital Course|9323,9330|false|false|false|C1314974|Cardiac attachment|Cardiac
Disorder|Disease or Syndrome|Hospital Course|9323,9340|false|false|false|C0007177|Cardiac Tamponade|Cardiac tamponade
Finding|Functional Concept|Hospital Course|9331,9340|false|false|false|C0332459|Compressed structure|tamponade
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9331,9340|false|false|false|C0579016||tamponade
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9350,9368|false|false|false|C0191234|Pericardiocentesis|pericardiocentesis
Drug|Substance|Hospital Course|9373,9378|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|Hospital Course|9373,9378|false|false|false|C1546604|Drain Specimen Code|drain
Procedure|Health Care Activity|Hospital Course|9379,9388|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9379,9388|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Finding|Functional Concept|Hospital Course|9408,9420|false|false|false|C0333348|Inflammatory|inflammatory
Disorder|Disease or Syndrome|Hospital Course|9421,9433|false|false|false|C0031046|Pericarditis|pericarditis
Finding|Finding|Hospital Course|9437,9445|false|false|false|C0332148|Probable diagnosis|probable
Finding|Functional Concept|Hospital Course|9446,9451|false|true|false|C0521026|Viral|viral
Finding|Functional Concept|Hospital Course|9453,9459|false|false|false|C0349590;C1262865|Nature;Natures|nature
Finding|Idea or Concept|Hospital Course|9453,9459|false|false|false|C0349590;C1262865|Nature;Natures|nature
Finding|Idea or Concept|Hospital Course|9467,9474|false|false|false|C0449255;C0542559;C4281677|Application Context;Context;contextual factors|context
Finding|Intellectual Product|Hospital Course|9467,9474|false|false|false|C0449255;C0542559;C4281677|Application Context;Context;contextual factors|context
Finding|Mental Process|Hospital Course|9467,9474|false|false|false|C0449255;C0542559;C4281677|Application Context;Context;contextual factors|context
Finding|Functional Concept|Hospital Course|9478,9483|false|false|false|C0521026|Viral|viral
Finding|Sign or Symptom|Hospital Course|9489,9497|false|false|false|C0240805|Prodrome|prodrome
Disorder|Disease or Syndrome|Hospital Course|9505,9514|false|false|false|C0035435|Rheumatism|rheumatic
Disorder|Disease or Syndrome|Hospital Course|9516,9528|false|false|false|C0031046|Pericarditis|pericarditis
Finding|Functional Concept|Hospital Course|9536,9545|false|false|false|C0205473|Serologic|serologic
Disorder|Cell or Molecular Dysfunction|Hospital Course|9546,9554|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Finding|Classification|Hospital Course|9546,9554|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|Hospital Course|9546,9554|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Disorder|Disease or Syndrome|Hospital Course|9562,9569|false|false|false|C0012634|Disease|disease
Disorder|Anatomical Abnormality|Hospital Course|9578,9585|false|false|false|C1689985|Absence (morphologic abnormality)|absence
Finding|Functional Concept|Hospital Course|9578,9585|false|false|false|C0332197|Absent|absence
Finding|Functional Concept|Hospital Course|9578,9588|false|false|false|C0332197|Absent|absence of
Drug|Pharmacologic Substance|Hospital Course|9589,9594|false|false|false|C0242708|Antirheumatic Drugs, Disease-Modifying|DMARD
Anatomy|Body Location or Region|Hospital Course|9596,9607|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|Pericardial
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9596,9607|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|Pericardial
Disorder|Disease or Syndrome|Hospital Course|9596,9613|false|false|false|C0031039|Pericardial effusion|Pericardial fluid
Finding|Body Substance|Hospital Course|9596,9613|false|false|false|C0225973|Pericardial fluid (substance)|Pericardial fluid
Procedure|Laboratory Procedure|Hospital Course|9596,9613|false|false|false|C3854061|pericardial fluid analysis|Pericardial fluid
Drug|Substance|Hospital Course|9608,9613|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|9608,9613|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Idea or Concept|Hospital Course|9614,9622|false|true|false|C0010453|Culture (Anthropological)|cultures
Finding|Classification|Hospital Course|9633,9641|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|9633,9641|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|9633,9641|false|false|false|C5237010|Expression Negative|negative
Finding|Idea or Concept|Hospital Course|9643,9651|false|false|false|C0010453|Culture (Anthropological)|cultures
Anatomy|Cell|Hospital Course|9664,9670|false|false|false|C1947989|Colony (cells or organisms)|colony
Procedure|Laboratory Procedure|Hospital Course|9685,9689|false|false|false|C0005790|Blood coagulation tests|coag
Finding|Classification|Hospital Course|9691,9699|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|9691,9699|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|9691,9699|false|false|false|C5237010|Expression Negative|negative
Disorder|Disease or Syndrome|Hospital Course|9700,9705|false|false|false|C0038160|Staphylococcal Infections|staph
Drug|Substance|Hospital Course|9717,9728|true|false|false|C2827365|Contaminant|contaminant
Finding|Classification|Hospital Course|9730,9738|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|9730,9738|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|9730,9738|false|false|false|C5237010|Expression Negative|negative
Drug|Indicator, Reagent, or Diagnostic Aid|Hospital Course|9739,9748|false|false|false|C1318720|Acid fast stain|acid fast
Finding|Finding|Hospital Course|9744,9748|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|fast
Finding|Gene or Genome|Hospital Course|9744,9748|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|fast
Finding|Molecular Function|Hospital Course|9744,9748|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|fast
Event|Activity|Hospital Course|9749,9754|false|false|false|C1947932|Smear - instruction imperative|smear
Finding|Functional Concept|Hospital Course|9749,9754|false|false|false|C3872789|Smearing technique|smear
Procedure|Diagnostic Procedure|Hospital Course|9749,9754|false|false|false|C0444186|Smear test|smear
Finding|Functional Concept|Hospital Course|9760,9771|false|false|false|C0205474|Biochemical|biochemical
Finding|Idea or Concept|Hospital Course|9772,9780|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Hospital Course|9772,9783|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Anatomy|Tissue|Hospital Course|9784,9794|false|false|false|C0027061|Myocardium|myocardial
Disorder|Injury or Poisoning|Hospital Course|9784,9801|true|false|false|C0746730|Myocardial injury|myocardial injury
Disorder|Injury or Poisoning|Hospital Course|9795,9801|true|false|false|C3263722;C3263723|Traumatic AND/OR non-traumatic injury;Traumatic injury|injury
Procedure|Health Care Activity|Hospital Course|9805,9814|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Finding|Hospital Course|9817,9825|false|false|false|C0750558|Unlikely|unlikely
Disorder|Disease or Syndrome|Hospital Course|9845,9856|false|false|false|C0027059|Myocarditis|myocarditis
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9860,9867|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|Hospital Course|9860,9867|false|false|false|C1314974|Cardiac attachment|cardiac
Disorder|Disease or Syndrome|Hospital Course|9860,9873|false|true|false|C0741923|Cardiac Events|cardiac event
Event|Event|Hospital Course|9868,9873|false|false|false|C0441471|Event|event
Finding|Pathologic Function|Hospital Course|9875,9883|false|false|false|C0243088;C0543419|Sequela of disorder;sequelae aspects|sequelae
Anatomy|Body Space or Junction|Hospital Course|9920,9924|false|false|false|C0228216|Structure of subparietal sulcus|SBPs
Drug|Substance|Hospital Course|9950,9955|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|9950,9955|false|false|false|C1546638|Fluid Specimen Code|fluid
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9950,9969|false|false|false|C0150238|Fluid resuscitation|fluid resuscitation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9956,9969|false|false|false|C0035273|Resuscitation (procedure)|resuscitation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9974,9992|false|false|false|C0191234|Pericardiocentesis|pericardiocentesis
Finding|Idea or Concept|Hospital Course|10000,10007|false|false|false|C2699424|Concern|concern
Finding|Functional Concept|Hospital Course|10012,10021|false|false|false|C0332459|Compressed structure|tamponade
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10012,10021|false|false|false|C0579016||tamponade
Finding|Physiologic Function|Hospital Course|10022,10032|false|false|false|C0031843|physiological aspects|physiology
Finding|Organ or Tissue Function|Hospital Course|10034,10046|false|false|false|C0019010|Hemodynamics|Hemodynamics
Procedure|Laboratory Procedure|Hospital Course|10034,10046|false|false|false|C4281788|hemodynamics (procedure)|Hemodynamics
Drug|Pharmacologic Substance|Hospital Course|10103,10111|false|false|false|C0720099|Duration brand of oxymetazoline|duration
Procedure|Health Care Activity|Hospital Course|10120,10129|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Procedure|Diagnostic Procedure|Hospital Course|10136,10139|false|false|false|C0430462|Transthoracic echocardiography|TTE
Anatomy|Body Location or Region|Hospital Course|10157,10168|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10157,10168|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Finding|Body Substance|Hospital Course|10170,10178|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|Hospital Course|10170,10178|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|Hospital Course|10170,10178|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Anatomy|Body Location or Region|Hospital Course|10180,10191|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|Pericardial
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10180,10191|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|Pericardial
Drug|Substance|Hospital Course|10192,10197|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|Hospital Course|10192,10197|false|false|false|C1546604|Drain Specimen Code|drain
Finding|Functional Concept|Hospital Course|10212,10216|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Phenomenon|Natural Phenomenon or Process|Hospital Course|10220,10227|false|false|false|C0282189|Gravity (physical force)|gravity
Finding|Conceptual Entity|Hospital Course|10246,10252|false|false|false|C1709366|system output|output
Procedure|Health Care Activity|Hospital Course|10246,10252|false|false|false|C3251815|Measurement of fluid output|output
Drug|Organic Chemical|Hospital Course|10296,10306|false|false|false|C0009262|colchicine|colchicine
Drug|Pharmacologic Substance|Hospital Course|10296,10306|false|false|false|C0009262|colchicine|colchicine
Disorder|Mental or Behavioral Dysfunction|Hospital Course|10313,10316|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10313,10316|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|10313,10316|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|10313,10316|false|false|false|C1332410|BID gene|BID
Finding|Body Substance|Hospital Course|10360,10369|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|10360,10369|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|10360,10369|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|10360,10369|false|false|false|C0030685|Patient Discharge|discharge
Drug|Organic Chemical|Hospital Course|10388,10397|false|false|false|C0020740|ibuprofen|ibuprofen
Drug|Pharmacologic Substance|Hospital Course|10388,10397|false|false|false|C0020740|ibuprofen|ibuprofen
Procedure|Health Care Activity|Hospital Course|10445,10450|false|false|false|C0441640||taper
Drug|Pharmacologic Substance|Hospital Course|10464,10467|false|false|false|C0358591|Proton Pump Inhibitors|PPI
Finding|Physiologic Function|Hospital Course|10464,10467|false|false|false|C0871125|Prepulse Inhibition|PPI
Drug|Pharmacologic Substance|Hospital Course|10485,10491|false|false|false|C0003211;C0358845|Analgesics and non-steroidal anti-inflammatory drugs;Anti-Inflammatory Agents, Non-Steroidal|NSAIDs
Finding|Intellectual Product|Hospital Course|10498,10503|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Disorder|Disease or Syndrome|Hospital Course|10498,10535|false|false|false|C4040419|Acute Hypercapnic Respiratory Failure|Acute hypercapnic respiratory failure
Finding|Finding|Hospital Course|10504,10515|false|false|false|C0020440|Hypercapnia|hypercapnic
Finding|Pathologic Function|Hospital Course|10504,10535|false|false|false|C0398353|Hypercapnic respiratory failure|hypercapnic respiratory failure
Attribute|Clinical Attribute|Hospital Course|10516,10527|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|Hospital Course|10516,10527|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|Hospital Course|10516,10527|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|Hospital Course|10516,10527|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Disorder|Disease or Syndrome|Hospital Course|10516,10535|false|false|false|C1145670|Respiratory Failure|respiratory failure
Finding|Functional Concept|Hospital Course|10528,10535|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|Hospital Course|10528,10535|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|Hospital Course|10528,10535|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Finding|Hospital Course|10548,10556|false|false|false|C0332148|Probable diagnosis|Probable
Finding|Gene or Genome|Hospital Course|10557,10562|false|true|false|C1413133;C4284306|CASP8AP2 gene;CASP8AP2 wt Allele|flash
Procedure|Diagnostic Procedure|Hospital Course|10557,10562|false|true|false|C0262485|Flash|flash
Disorder|Disease or Syndrome|Hospital Course|10557,10578|false|true|false|C1168329|Flash pulmonary oedema|flash pulmonary edema
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10563,10572|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Hospital Course|10563,10572|false|true|false|C2707265||pulmonary
Finding|Finding|Hospital Course|10563,10572|false|true|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|Hospital Course|10563,10578|false|true|false|C0034063|Pulmonary Edema|pulmonary edema
Attribute|Clinical Attribute|Hospital Course|10573,10578|false|true|false|C1717255||edema
Finding|Pathologic Function|Hospital Course|10573,10578|false|true|false|C0013604|Edema|edema
Finding|Gene or Genome|Hospital Course|10590,10595|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Finding|Intellectual Product|Hospital Course|10596,10602|false|false|false|C1705102|Volume (publication)|volume
Drug|Substance|Hospital Course|10603,10608|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|10603,10608|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Occupational Activity|Hospital Course|10610,10624|false|false|false|C0001554|Administration occupational activities|administration
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10610,10624|false|false|false|C1533734|Administration (procedure)|administration
Finding|Functional Concept|Hospital Course|10628,10637|false|false|false|C0332459|Compressed structure|tamponade
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10628,10637|false|false|false|C0579016||tamponade
Phenomenon|Natural Phenomenon or Process|Hospital Course|10655,10667|false|false|false|C0444708|Radiographic|radiographic
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10669,10678|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Hospital Course|10669,10678|false|false|false|C2707265||pulmonary
Finding|Finding|Hospital Course|10669,10678|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|Hospital Course|10669,10684|false|false|false|C0034063|Pulmonary Edema|pulmonary edema
Attribute|Clinical Attribute|Hospital Course|10679,10684|false|false|false|C1717255||edema
Finding|Pathologic Function|Hospital Course|10679,10684|false|false|false|C0013604|Edema|edema
Procedure|Diagnostic Procedure|Hospital Course|10694,10708|false|false|false|C0013516|Echocardiography|echocardiogram
Finding|Functional Concept|Hospital Course|10723,10733|true|false|false|C0332299|Suggestive of|suggestive
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10738,10749|false|false|false|C0018827|Heart Ventricle|ventricular
Finding|Pathologic Function|Hospital Course|10738,10761|false|false|false|C0242973|Ventricular Dysfunction|ventricular dysfunction
Disorder|Disease or Syndrome|Hospital Course|10750,10761|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Finding|Conceptual Entity|Hospital Course|10750,10761|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|Hospital Course|10750,10761|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|Hospital Course|10750,10761|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10766,10769|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Hormone|Hospital Course|10766,10769|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Pharmacologic Substance|Hospital Course|10766,10769|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Finding|Gene or Genome|Hospital Course|10766,10769|false|false|false|C1417808;C2982014|NPPB gene;NPPB wt Allele|BNP
Procedure|Laboratory Procedure|Hospital Course|10766,10769|false|false|false|C1095989|Brain natriuretic peptide measurement|BNP
Procedure|Diagnostic Procedure|Hospital Course|10795,10798|false|false|false|C0430462|Transthoracic echocardiography|TTE
Finding|Idea or Concept|Hospital Course|10819,10827|false|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Hospital Course|10819,10830|false|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10831,10838|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|Hospital Course|10831,10838|true|false|false|C1314974|Cardiac attachment|cardiac
Disorder|Disease or Syndrome|Hospital Course|10831,10847|true|false|false|C0741922|CARDIAC ETIOLOGY|cardiac etiology
Finding|Conceptual Entity|Hospital Course|10839,10847|true|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|etiology
Finding|Functional Concept|Hospital Course|10839,10847|true|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|etiology
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10857,10866|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Hospital Course|10857,10866|false|false|false|C2707265||pulmonary
Finding|Finding|Hospital Course|10857,10866|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|Hospital Course|10857,10872|false|false|false|C0034063|Pulmonary Edema|pulmonary edema
Attribute|Clinical Attribute|Hospital Course|10867,10872|false|false|false|C1717255||edema
Finding|Pathologic Function|Hospital Course|10867,10872|false|false|false|C0013604|Edema|edema
Attribute|Clinical Attribute|Hospital Course|10873,10884|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|Hospital Course|10873,10884|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|Hospital Course|10873,10884|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|Hospital Course|10873,10884|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Disorder|Disease or Syndrome|Hospital Course|10873,10892|false|false|false|C1145670|Respiratory Failure|respiratory failure
Finding|Functional Concept|Hospital Course|10885,10892|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|Hospital Course|10885,10892|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|Hospital Course|10885,10892|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Body Substance|Hospital Course|10894,10901|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|10894,10901|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|10894,10901|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Finding|Hospital Course|10902,10908|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|10902,10908|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10939,10948|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Hospital Course|10939,10948|false|false|false|C2707265||pulmonary
Finding|Finding|Hospital Course|10939,10948|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Physiologic Function|Hospital Course|10950,10960|false|false|false|C0031843|physiological aspects|physiology
Finding|Functional Concept|Hospital Course|10979,10992|true|false|false|C0333159|Emphysematous|emphysematous
Finding|Functional Concept|Hospital Course|10993,11000|true|false|false|C0392747|Changing|changes
Finding|Intellectual Product|Hospital Course|11018,11022|false|false|false|C1561540|Transaction counts and value totals - week|week
Finding|Gene or Genome|Hospital Course|11023,11026|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Finding|Conceptual Entity|Hospital Course|11032,11042|false|false|false|C1706907|Background|background
Finding|Functional Concept|Hospital Course|11043,11054|false|false|false|C0549186|Obstructed|obstructive
Disorder|Disease or Syndrome|Hospital Course|11055,11061|false|false|false|C1861101|THYROID HORMONE PLASMA MEMBRANE TRANSPORT DEFECT|defect
Finding|Functional Concept|Hospital Course|11055,11061|false|false|false|C1457869|Defect|defect
Finding|Conceptual Entity|Hospital Course|11103,11110|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|11103,11110|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|11103,11110|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Classification|Hospital Course|11121,11129|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|11121,11129|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|11121,11129|false|false|false|C5237010|Expression Negative|negative
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11130,11133|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Finding|Gene or Genome|Hospital Course|11130,11133|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|Hospital Course|11130,11133|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Finding|Intellectual Product|Hospital Course|11138,11142|false|false|false|C1561540|Transaction counts and value totals - week|week
Procedure|Health Care Activity|Hospital Course|11153,11162|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Body Substance|Hospital Course|11164,11171|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|11164,11171|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|11164,11171|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Disorder|Disease or Syndrome|Hospital Course|11176,11188|false|false|false|C0023518|Leukocytosis|leukocytosis
Finding|Finding|Hospital Course|11176,11188|false|false|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Procedure|Health Care Activity|Hospital Course|11192,11201|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Idea or Concept|Hospital Course|11210,11215|false|false|false|C1550016|Remote control command - Clear|clear
Phenomenon|Natural Phenomenon or Process|Hospital Course|11217,11229|false|false|false|C0444708|Radiographic|radiographic
Disorder|Disease or Syndrome|Hospital Course|11230,11243|false|false|false|C0521530|Lung consolidation|consolidation
Finding|Functional Concept|Hospital Course|11244,11254|false|false|false|C0332299|Suggestive of|suggestive
Finding|Functional Concept|Hospital Course|11244,11257|false|false|false|C0332299|Suggestive of|suggestive of
Disorder|Disease or Syndrome|Hospital Course|11258,11267|false|false|false|C0032285|Pneumonia|pneumonia
Drug|Antibiotic|Hospital Course|11291,11303|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|Hospital Course|11291,11303|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|Hospital Course|11291,11303|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Finding|Organ or Tissue Function|Hospital Course|11365,11373|false|false|false|C0012797|Diuresis|diuresis
Finding|Idea or Concept|Hospital Course|11379,11390|false|false|false|C0750502|Significant|significant
Finding|Conceptual Entity|Hospital Course|11391,11402|false|false|false|C2986411|Improvement|improvement
Attribute|Clinical Attribute|Hospital Course|11411,11422|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|Hospital Course|11411,11422|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|Hospital Course|11411,11422|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|Hospital Course|11411,11422|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Attribute|Clinical Attribute|Hospital Course|11411,11429|false|false|false|C2598168||respiratory status
Finding|Finding|Hospital Course|11411,11429|false|false|false|C1998827|Respiratory Status|respiratory status
Attribute|Clinical Attribute|Hospital Course|11423,11429|false|false|false|C5889824||status
Finding|Idea or Concept|Hospital Course|11423,11429|false|false|false|C1546481|What subject filter - Status|status
Finding|Finding|Hospital Course|11497,11501|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Hospital Course|11497,11501|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Hospital Course|11497,11501|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Body Substance|Hospital Course|11505,11514|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|11505,11514|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|11505,11514|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|11505,11514|false|false|false|C0030685|Patient Discharge|discharge
Finding|Functional Concept|Hospital Course|11520,11530|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|ambulatory
Finding|Idea or Concept|Hospital Course|11520,11530|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|ambulatory
Finding|Intellectual Product|Hospital Course|11520,11530|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|ambulatory
Procedure|Health Care Activity|Hospital Course|11520,11530|false|false|false|C1561560|ambulatory encounter|ambulatory
Phenomenon|Natural Phenomenon or Process|Hospital Course|11532,11543|false|false|false|C0522534|Saturated|saturations
Disorder|Disease or Syndrome|Hospital Course|11566,11570|false|false|false|C0004238|Atrial Fibrillation|AFib
Lab|Laboratory or Test Result|Hospital Course|11566,11570|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|AFib
Finding|Finding|Hospital Course|11572,11575|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Hospital Course|11572,11575|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Finding|Hospital Course|11572,11585|false|false|false|C2585997|New diagnosis (finding)|new diagnosis
Procedure|Diagnostic Procedure|Hospital Course|11572,11585|false|false|false|C1882082|New Diagnosis Procedure|new diagnosis
Attribute|Clinical Attribute|Hospital Course|11576,11585|false|false|false|C0945731||diagnosis
Finding|Classification|Hospital Course|11576,11585|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|Hospital Course|11576,11585|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|Hospital Course|11576,11585|false|false|false|C0011900|Diagnosis|diagnosis
Finding|Body Substance|Hospital Course|11587,11594|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|11587,11594|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|11587,11594|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Disorder|Disease or Syndrome|Hospital Course|11605,11609|false|false|false|C0004238|Atrial Fibrillation|Afib
Lab|Laboratory or Test Result|Hospital Course|11605,11609|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Afib
Finding|Finding|Hospital Course|11615,11618|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Finding|Gene or Genome|Hospital Course|11615,11618|false|false|false|C1417822;C3540498;C4050414|NR1D2 gene;NR1D2 wt Allele;Rapid Virologic Response|RVR
Drug|Organic Chemical|Hospital Course|11654,11664|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|Hospital Course|11654,11664|false|false|false|C0025859|metoprolol|metoprolol
Finding|Molecular Function|Hospital Course|11700,11703|false|false|false|C1704493;C2700623|Neutral Sidebent Rotated|NSR
Finding|Pathologic Function|Hospital Course|11700,11703|false|false|false|C1704493;C2700623|Neutral Sidebent Rotated|NSR
Disorder|Disease or Syndrome|Hospital Course|11729,11732|false|false|false|C0020538|Hypertensive disease|HTN
Finding|Finding|Hospital Course|11735,11750|false|false|true|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|Anticoagulation
Finding|Physiologic Function|Hospital Course|11735,11750|false|false|true|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|Anticoagulation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11735,11750|false|false|true|C0003281|Anticoagulation Therapy|Anticoagulation
Finding|Finding|Hospital Course|11797,11801|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Hospital Course|11797,11801|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Hospital Course|11797,11801|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Body Substance|Hospital Course|11805,11814|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|11805,11814|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|11805,11814|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|11805,11814|false|false|false|C0030685|Patient Discharge|discharge
Finding|Body Substance|Hospital Course|11825,11832|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|11825,11832|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|11825,11832|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Anatomy|Body Location or Region|Hospital Course|11836,11841|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|Hospital Course|11836,11841|false|false|false|C2003888|Lower (action)|lower
Finding|Intellectual Product|Hospital Course|11842,11849|false|false|false|C0282416|Overall Publication Type|overall
Finding|Idea or Concept|Hospital Course|11850,11854|false|false|false|C0035647|Risk|risk
Disorder|Disease or Syndrome|Hospital Course|11859,11862|false|false|false|C0001365;C0038454|Acute ill-defined cerebrovascular disease;Cerebrovascular accident|CVA
Drug|Pharmacologic Substance|Hospital Course|11859,11862|false|false|false|C5779650|Cyclophosphamide/Doxorubicin/Vincristine|CVA
Drug|Pharmacologic Substance|Hospital Course|11886,11896|false|false|false|C0013227|Pharmaceutical Preparations|medication
Finding|Intellectual Product|Hospital Course|11886,11896|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Finding|Functional Concept|Hospital Course|11898,11907|false|false|false|C1510802|Adherence (attribute)|adherence
Finding|Functional Concept|Hospital Course|11908,11912|false|false|false|C0220812;C4050363|Comprehensive Score for Financial Toxicity;Cost aspects|cost
Finding|Intellectual Product|Hospital Course|11908,11912|false|false|false|C0220812;C4050363|Comprehensive Score for Financial Toxicity;Cost aspects|cost
Drug|Organic Chemical|Hospital Course|11935,11945|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|Hospital Course|11935,11945|false|false|false|C0025859|metoprolol|metoprolol
Finding|Functional Concept|Hospital Course|11967,11971|false|false|false|C0686904|Patient need for (contextual qualifier)|need
Finding|Functional Concept|Hospital Course|11967,11975|false|false|false|C0686904|Patient need for (contextual qualifier)|need for
Finding|Finding|Hospital Course|11976,11991|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|Hospital Course|11976,11991|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11976,11991|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Finding|Classification|Hospital Course|12009,12019|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|12009,12019|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Gene or Genome|Hospital Course|12052,12056|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|Type
Finding|Intellectual Product|Hospital Course|12052,12056|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|Type
Disorder|Disease or Syndrome|Hospital Course|12052,12068|false|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|Type II diabetes
Disorder|Disease or Syndrome|Hospital Course|12060,12068|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|diabetes
Finding|Idea or Concept|Hospital Course|12078,12083|false|false|false|C0750546|newly|newly
Finding|Classification|Hospital Course|12109,12112|false|false|false|C4521595|United States Military enlisted E3 (qualifier value)|A1C
Procedure|Laboratory Procedure|Hospital Course|12109,12112|false|false|false|C0474680|Hemoglobin A1c measurement|A1C
Procedure|Health Care Activity|Hospital Course|12134,12143|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12169,12176|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|Hospital Course|12169,12176|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|Hospital Course|12169,12176|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Finding|Gene or Genome|Hospital Course|12169,12176|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|Hospital Course|12169,12176|false|false|false|C0202098|Insulin measurement|insulin
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12185,12190|false|false|false|C0222045|Integumentary scale|scale
Event|Activity|Hospital Course|12185,12190|false|false|false|C1947916|Scaling|scale
Finding|Conceptual Entity|Hospital Course|12185,12190|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Finding|Intellectual Product|Hospital Course|12185,12190|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Procedure|Health Care Activity|Hospital Course|12204,12213|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Drug|Organic Chemical|Hospital Course|12240,12249|false|false|false|C0025598|metformin|metformin
Drug|Pharmacologic Substance|Hospital Course|12240,12249|false|false|false|C0025598|metformin|metformin
Disorder|Mental or Behavioral Dysfunction|Hospital Course|12256,12259|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12256,12259|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|12256,12259|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|12256,12259|false|false|false|C1332410|BID gene|BID
Finding|Intellectual Product|Hospital Course|12263,12270|false|false|false|C1547296|Chronic - Admission Level of Care Code|CHRONIC
Procedure|Health Care Activity|Hospital Course|12263,12270|false|false|false|C1555457|Provision of recurring care for chronic illness|CHRONIC
Finding|Intellectual Product|Hospital Course|12271,12277|false|false|false|C1547311|Patient Condition Code - Stable|STABLE
Disorder|Disease or Syndrome|Hospital Course|12310,12330|false|false|false|C0003873|Rheumatoid Arthritis|Rheumatoid arthritis
Disorder|Disease or Syndrome|Hospital Course|12321,12330|false|false|false|C0003864|Arthritis|arthritis
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12340,12348|false|false|false|C4318437|Anti-Cyclic Citrullinated Protein Antibodies|anti-CCP
Drug|Immunologic Factor|Hospital Course|12340,12348|false|false|false|C4318437|Anti-Cyclic Citrullinated Protein Antibodies|anti-CCP
Disorder|Cell or Molecular Dysfunction|Hospital Course|12349,12357|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Finding|Classification|Hospital Course|12349,12357|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|Hospital Course|12349,12357|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Classification|Hospital Course|12362,12372|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|12362,12372|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Functional Concept|Hospital Course|12414,12424|false|false|false|C0332299|Suggestive of|suggestive
Finding|Functional Concept|Hospital Course|12414,12427|false|false|false|C0332299|Suggestive of|suggestive of
Finding|Finding|Hospital Course|12431,12436|false|false|false|C1517205;C3540542|Exacerbation of cGVHD;Flare|flare
Finding|Sign or Symptom|Hospital Course|12431,12436|false|false|false|C1517205;C3540542|Exacerbation of cGVHD;Flare|flare
Finding|Social Behavior|Hospital Course|12442,12452|false|false|false|C2584313|Discussion (communication)|discussion
Procedure|Therapeutic or Preventive Procedure|Hospital Course|12442,12452|false|false|false|C0557061|Discussion (procedure)|discussion
Drug|Organic Chemical|Hospital Course|12497,12500|false|false|false|C0025677|methotrexate|MTX
Drug|Pharmacologic Substance|Hospital Course|12497,12500|false|false|false|C0025677|methotrexate|MTX
Finding|Gene or Genome|Hospital Course|12497,12500|false|false|false|C1417487;C5891182|MTX1 gene;Matrix Market File Format|MTX
Finding|Intellectual Product|Hospital Course|12497,12500|false|false|false|C1417487;C5891182|MTX1 gene;Matrix Market File Format|MTX
Drug|Pharmacologic Substance|Hospital Course|12514,12519|false|false|false|C0242708|Antirheumatic Drugs, Disease-Modifying|DMARD
Finding|Classification|Hospital Course|12526,12536|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|12526,12536|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Disorder|Disease or Syndrome|Hospital Course|12542,12545|false|false|false|C0020538|Hypertensive disease|HTN
Finding|Idea or Concept|Hospital Course|12550,12554|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|12550,12554|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|12550,12554|false|false|false|C1553498|home health encounter|home
Disorder|Disease or Syndrome|Hospital Course|12558,12562|false|false|false|C3280240|MICROCEPHALY, EPILEPSY, AND DIABETES SYNDROME 1|meds
Finding|Intellectual Product|Hospital Course|12558,12562|false|false|false|C4284232|Medications|meds
Disorder|Disease or Syndrome|Hospital Course|12590,12594|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Disorder|Disease or Syndrome|Hospital Course|12595,12598|false|false|false|C1849718|POPLITEAL PTERYGIUM SYNDROME, LETHAL TYPE|BPs
Drug|Organic Chemical|Hospital Course|12595,12598|false|false|false|C2740858|BPS|BPs
Drug|Pharmacologic Substance|Hospital Course|12595,12598|false|false|false|C2740858|BPS|BPs
Finding|Finding|Hospital Course|12624,12628|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Hospital Course|12624,12628|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Hospital Course|12624,12628|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Body Substance|Hospital Course|12632,12641|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|12632,12641|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|12632,12641|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|12632,12641|false|false|false|C0030685|Patient Discharge|discharge
Anatomy|Cell Component|Hospital Course|12673,12677|false|false|false|C1167518|viral nucleocapsid location|CORE
Finding|Body Substance|Hospital Course|12673,12677|false|false|false|C3274653|Core Specimen|CORE
Finding|Functional Concept|Hospital Course|12678,12686|false|false|false|C1879489|Measures (attribute)|MEASURES
Event|Occupational Activity|Hospital Course|12706,12710|false|false|false|C0009219|Coding|CODE
Finding|Intellectual Product|Hospital Course|12706,12710|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|CODE
Attribute|Clinical Attribute|Hospital Course|12712,12715|false|false|false|C4285234||DNR
Drug|Antibiotic|Hospital Course|12712,12715|false|false|false|C0011015|daunorubicin|DNR
Drug|Organic Chemical|Hospital Course|12712,12715|false|false|false|C0011015|daunorubicin|DNR
Finding|Finding|Hospital Course|12712,12715|false|false|false|C0079252;C0582114|Do not resuscitate status;Do-Not-Resuscitate Orders|DNR
Finding|Intellectual Product|Hospital Course|12712,12715|false|false|false|C0079252;C0582114|Do not resuscitate status;Do-Not-Resuscitate Orders|DNR
Event|Activity|Hospital Course|12722,12729|false|false|false|C3812666|Personal Contact|CONTACT
Finding|Functional Concept|Hospital Course|12722,12729|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Idea or Concept|Hospital Course|12722,12729|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Intellectual Product|Hospital Course|12722,12729|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Phenomenon|Phenomenon or Process|Hospital Course|12722,12729|false|false|false|C0392367|Physical contact|CONTACT
Disorder|Disease or Syndrome|Hospital Course|12730,12733|false|false|false|C0162531|Hereditary Coproporphyria|HCP
Finding|Gene or Genome|Hospital Course|12730,12733|false|false|false|C1335283;C1412376;C1413681;C1705637;C5780748|AMBP gene;AMBP wt Allele;CPOX gene;PTPN6 gene;PTPN6 wt Allele|HCP
Attribute|Clinical Attribute|Hospital Course|12757,12768|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|12757,12768|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Hospital Course|12757,12768|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|12757,12781|false|false|false|C1627937|Medications on admission|Medications on Admission
Procedure|Health Care Activity|Hospital Course|12772,12781|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|Hospital Course|12800,12810|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Hospital Course|12800,12810|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|Hospital Course|12800,12815|false|false|false|C0746470|MEDICATION LIST|Medication list
Finding|Intellectual Product|Hospital Course|12811,12815|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Drug|Organic Chemical|Hospital Course|12832,12840|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Hospital Course|12832,12840|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Hospital Course|12832,12840|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Finding|Functional Concept|Hospital Course|12832,12840|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|12832,12840|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|Hospital Course|12845,12857|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|12845,12857|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|Hospital Course|12875,12885|false|false|false|C0009262|colchicine|Colchicine
Drug|Pharmacologic Substance|Hospital Course|12875,12885|false|false|false|C0009262|colchicine|Colchicine
Disorder|Mental or Behavioral Dysfunction|Hospital Course|12896,12899|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12896,12899|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|12896,12899|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|12896,12899|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|12904,12913|false|false|false|C0020740|ibuprofen|Ibuprofen
Drug|Pharmacologic Substance|Hospital Course|12904,12913|false|false|false|C0020740|ibuprofen|Ibuprofen
Drug|Organic Chemical|Hospital Course|12932,12942|false|false|false|C0015620|famotidine|Famotidine
Drug|Pharmacologic Substance|Hospital Course|12932,12942|false|false|false|C0015620|famotidine|Famotidine
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12962,12972|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|Hospital Course|12962,12972|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|Hospital Course|12962,12992|false|false|false|C0717824|hydrochlorothiazide / lisinopril|lisinopril-hydrochlorothiazide
Drug|Organic Chemical|Hospital Course|12973,12992|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Drug|Pharmacologic Substance|Hospital Course|12973,12992|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Anatomy|Body Space or Junction|Hospital Course|13000,13004|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|13000,13004|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|13000,13004|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|13000,13004|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Organic Chemical|Hospital Course|13015,13027|false|false|false|C0025677|methotrexate|Methotrexate
Drug|Pharmacologic Substance|Hospital Course|13015,13027|false|false|false|C0025677|methotrexate|Methotrexate
Procedure|Laboratory Procedure|Hospital Course|13015,13027|false|false|false|C5399953|Drug assay methotrexate|Methotrexate
Finding|Intellectual Product|Hospital Course|13040,13044|false|false|false|C1561540|Transaction counts and value totals - week|WEEK
Drug|Organic Chemical|Hospital Course|13055,13065|false|false|false|C0074393|sertraline|Sertraline
Drug|Pharmacologic Substance|Hospital Course|13055,13065|false|false|false|C0074393|sertraline|Sertraline
Drug|Organic Chemical|Hospital Course|13086,13096|false|false|false|C0016410|folic acid|FoLIC Acid
Drug|Pharmacologic Substance|Hospital Course|13086,13096|false|false|false|C0016410|folic acid|FoLIC Acid
Drug|Vitamin|Hospital Course|13086,13096|false|false|false|C0016410|folic acid|FoLIC Acid
Procedure|Laboratory Procedure|Hospital Course|13086,13096|false|false|false|C0523631|Folic acid measurement|FoLIC Acid
Finding|Body Substance|Hospital Course|13115,13124|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|13115,13124|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|13115,13124|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|13115,13124|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|13115,13136|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|13125,13136|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|13125,13136|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Hospital Course|13125,13136|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|13142,13151|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|Hospital Course|13142,13151|false|false|false|C0001927|albuterol|Albuterol
Finding|Functional Concept|Hospital Course|13152,13159|false|false|false|C4319647|Inhaler (unit of presentation)|Inhaler
Finding|Gene or Genome|Hospital Course|13174,13177|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Body Substance|Hospital Course|13202,13208|false|false|false|C0225386|Breath|breath
Drug|Organic Chemical|Hospital Course|13214,13223|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|Hospital Course|13214,13223|false|false|false|C0001927|albuterol|albuterol
Drug|Organic Chemical|Hospital Course|13214,13231|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|Hospital Course|13214,13231|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|Hospital Course|13224,13231|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|Hospital Course|13224,13231|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|Hospital Course|13224,13231|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Organic Chemical|Hospital Course|13233,13239|false|false|false|C0162684;C1739179|Pro-Air Procaterol;ProAir|ProAir
Drug|Pharmacologic Substance|Hospital Course|13233,13239|false|false|false|C0162684;C1739179|Pro-Air Procaterol;ProAir|ProAir
Drug|Organic Chemical|Hospital Course|13233,13243|false|false|false|C1739179|ProAir|ProAir HFA
Drug|Pharmacologic Substance|Hospital Course|13233,13243|false|false|false|C1739179|ProAir|ProAir HFA
Disorder|Disease or Syndrome|Hospital Course|13240,13243|false|false|false|C0015458|Facial Hemiatrophy|HFA
Procedure|Diagnostic Procedure|Hospital Course|13240,13243|false|false|false|C0430649|High frequency audiometry|HFA
Finding|Functional Concept|Hospital Course|13297,13304|false|false|false|C4319647|Inhaler (unit of presentation)|Inhaler
Finding|Idea or Concept|Hospital Course|13305,13312|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|13321,13330|false|false|false|C0025598|metformin|MetFORMIN
Drug|Pharmacologic Substance|Hospital Course|13321,13330|false|false|false|C0025598|metformin|MetFORMIN
Drug|Organic Chemical|Hospital Course|13332,13342|false|false|false|C0591573|Glucophage|Glucophage
Drug|Pharmacologic Substance|Hospital Course|13332,13342|false|false|false|C0591573|Glucophage|Glucophage
Disorder|Mental or Behavioral Dysfunction|Hospital Course|13354,13357|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|13354,13357|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|13354,13357|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|13354,13357|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|13363,13372|false|false|false|C0025598|metformin|metformin
Drug|Pharmacologic Substance|Hospital Course|13363,13372|false|false|false|C0025598|metformin|metformin
Drug|Biomedical or Dental Material|Hospital Course|13382,13388|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|13392,13400|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|13395,13400|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|13395,13400|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|Hospital Course|13409,13412|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|13409,13412|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biomedical or Dental Material|Hospital Course|13424,13430|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|13431,13438|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|13447,13457|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|Hospital Course|13447,13457|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|Hospital Course|13447,13467|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Pharmacologic Substance|Hospital Course|13447,13467|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Organic Chemical|Hospital Course|13458,13467|false|false|false|C0038617;C0220918|Succinates;succinate|Succinate
Drug|Organic Chemical|Hospital Course|13491,13501|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|Hospital Course|13491,13501|false|false|false|C0025859|metoprolol|metoprolol
Drug|Organic Chemical|Hospital Course|13491,13511|false|false|false|C0724633|metoprolol succinate|metoprolol succinate
Drug|Pharmacologic Substance|Hospital Course|13491,13511|false|false|false|C0724633|metoprolol succinate|metoprolol succinate
Drug|Organic Chemical|Hospital Course|13502,13511|false|false|false|C0038617;C0220918|Succinates;succinate|succinate
Drug|Biomedical or Dental Material|Hospital Course|13520,13526|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|13530,13538|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|13533,13538|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|13533,13538|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Activity|Hospital Course|13545,13549|false|false|false|C1880359|Dispense (activity)|Disp
Finding|Gene or Genome|Hospital Course|13545,13549|false|false|false|C2828567|PRSS30P gene|Disp
Drug|Biomedical or Dental Material|Hospital Course|13556,13562|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|13563,13570|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|13579,13589|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Pharmacologic Substance|Hospital Course|13579,13589|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Organic Chemical|Hospital Course|13610,13620|false|false|false|C0028978|omeprazole|omeprazole
Drug|Pharmacologic Substance|Hospital Course|13610,13620|false|false|false|C0028978|omeprazole|omeprazole
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|13629,13636|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|Hospital Course|13629,13636|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|Hospital Course|13629,13636|false|false|false|C0006935|capsule (pharmacologic)|capsule
Finding|Functional Concept|Hospital Course|13640,13648|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|13643,13648|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|13643,13648|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|13666,13673|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|13666,13673|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|13666,13673|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Finding|Idea or Concept|Hospital Course|13674,13681|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|13690,13702|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|13690,13702|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|Hospital Course|13722,13732|false|false|false|C0009262|colchicine|Colchicine
Drug|Pharmacologic Substance|Hospital Course|13722,13732|false|false|false|C0009262|colchicine|Colchicine
Disorder|Mental or Behavioral Dysfunction|Hospital Course|13743,13746|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|13743,13746|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|13743,13746|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|13743,13746|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|13752,13762|false|false|false|C0009262|colchicine|colchicine
Drug|Pharmacologic Substance|Hospital Course|13752,13762|false|false|false|C0009262|colchicine|colchicine
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|13772,13779|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|Hospital Course|13772,13779|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|Hospital Course|13772,13779|false|false|false|C0006935|capsule (pharmacologic)|capsule
Finding|Functional Concept|Hospital Course|13783,13791|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|13786,13791|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|13786,13791|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|Hospital Course|13800,13803|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|13800,13803|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Activity|Hospital Course|13804,13808|false|false|false|C1880359|Dispense (activity)|Disp
Finding|Gene or Genome|Hospital Course|13804,13808|false|false|false|C2828567|PRSS30P gene|Disp
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|13815,13822|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|13815,13822|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|13815,13822|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Finding|Idea or Concept|Hospital Course|13823,13830|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|13839,13849|false|false|false|C0016410|folic acid|FoLIC Acid
Drug|Pharmacologic Substance|Hospital Course|13839,13849|false|false|false|C0016410|folic acid|FoLIC Acid
Drug|Vitamin|Hospital Course|13839,13849|false|false|false|C0016410|folic acid|FoLIC Acid
Procedure|Laboratory Procedure|Hospital Course|13839,13849|false|false|false|C0523631|Folic acid measurement|FoLIC Acid
Drug|Organic Chemical|Hospital Course|13870,13879|false|false|false|C0020740|ibuprofen|Ibuprofen
Drug|Pharmacologic Substance|Hospital Course|13870,13879|false|false|false|C0020740|ibuprofen|Ibuprofen
Drug|Organic Chemical|Hospital Course|13900,13910|false|false|false|C0074393|sertraline|Sertraline
Drug|Pharmacologic Substance|Hospital Course|13900,13910|false|false|false|C0074393|sertraline|Sertraline
Drug|Amino Acid, Peptide, or Protein|Hospital Course|13933,13937|false|false|false|C0675390|ARID1A protein, human|HELD
Drug|Biologically Active Substance|Hospital Course|13933,13937|false|false|false|C0675390|ARID1A protein, human|HELD
Finding|Gene or Genome|Hospital Course|13933,13937|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|HELD
Finding|Idea or Concept|Hospital Course|13933,13937|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|HELD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|13939,13949|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|Hospital Course|13939,13949|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|Hospital Course|13939,13969|false|false|false|C0717824|hydrochlorothiazide / lisinopril|lisinopril-hydrochlorothiazide
Drug|Organic Chemical|Hospital Course|13950,13969|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Drug|Pharmacologic Substance|Hospital Course|13950,13969|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Anatomy|Body Space or Junction|Hospital Course|13977,13981|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|13977,13981|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|13977,13981|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|13977,13981|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Pharmacologic Substance|Hospital Course|13995,14005|false|false|false|C0013227|Pharmaceutical Preparations|medication
Finding|Intellectual Product|Hospital Course|13995,14005|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Drug|Amino Acid, Peptide, or Protein|Hospital Course|14032,14042|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|Hospital Course|14032,14042|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|Hospital Course|14032,14062|false|false|false|C0717824|hydrochlorothiazide / lisinopril|lisinopril-hydrochlorothiazide
Drug|Organic Chemical|Hospital Course|14043,14062|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Drug|Pharmacologic Substance|Hospital Course|14043,14062|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Event|Activity|Hospital Course|14097,14101|false|false|false|C1947933|care activity|care
Finding|Finding|Hospital Course|14097,14101|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Hospital Course|14097,14101|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Hospital Course|14102,14108|false|false|false|C2348314|Doctor - Title|doctor
Drug|Amino Acid, Peptide, or Protein|Hospital Course|14129,14133|false|false|false|C0675390|ARID1A protein, human|HELD
Drug|Biologically Active Substance|Hospital Course|14129,14133|false|false|false|C0675390|ARID1A protein, human|HELD
Finding|Gene or Genome|Hospital Course|14129,14133|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|HELD
Finding|Idea or Concept|Hospital Course|14129,14133|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|HELD
Drug|Organic Chemical|Hospital Course|14135,14147|false|false|false|C0025677|methotrexate|Methotrexate
Drug|Pharmacologic Substance|Hospital Course|14135,14147|false|false|false|C0025677|methotrexate|Methotrexate
Procedure|Laboratory Procedure|Hospital Course|14135,14147|false|false|false|C5399953|Drug assay methotrexate|Methotrexate
Finding|Intellectual Product|Hospital Course|14160,14164|false|false|false|C1561540|Transaction counts and value totals - week|WEEK
Drug|Pharmacologic Substance|Hospital Course|14177,14187|false|false|false|C0013227|Pharmaceutical Preparations|medication
Finding|Intellectual Product|Hospital Course|14177,14187|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Drug|Organic Chemical|Hospital Course|14214,14226|false|false|false|C0025677|methotrexate|Methotrexate
Drug|Pharmacologic Substance|Hospital Course|14214,14226|false|false|false|C0025677|methotrexate|Methotrexate
Procedure|Laboratory Procedure|Hospital Course|14214,14226|false|false|false|C5399953|Drug assay methotrexate|Methotrexate
Finding|Intellectual Product|Hospital Course|14235,14241|false|false|false|C2348314|Doctor - Title|doctor
Finding|Body Substance|Hospital Course|14259,14268|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|14259,14268|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|14259,14268|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|14259,14268|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|14259,14280|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|14259,14280|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|14269,14280|false|false|false|C2926604||Disposition
Procedure|Health Care Activity|Hospital Course|14269,14280|false|false|false|C0184758|Patient disposition|Disposition
Finding|Idea or Concept|Hospital Course|14282,14286|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|14282,14286|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|14282,14286|false|false|false|C1553498|home health encounter|Home
Finding|Body Substance|Hospital Course|14289,14298|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|14289,14298|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|14289,14298|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|14289,14298|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|14289,14308|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|14299,14308|false|false|false|C0945731||Diagnosis
Finding|Classification|Hospital Course|14299,14308|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|14299,14308|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|14299,14308|false|false|false|C0011900|Diagnosis|Diagnosis
Attribute|Clinical Attribute|Hospital Course|14310,14327|false|false|false|C0801658||Primary Diagnosis
Attribute|Clinical Attribute|Hospital Course|14318,14327|false|false|false|C0945731||Diagnosis
Finding|Classification|Hospital Course|14318,14327|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|14318,14327|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|14318,14327|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Functional Concept|Hospital Course|14329,14341|false|false|false|C0333348|Inflammatory|inflammatory
Disorder|Disease or Syndrome|Hospital Course|14342,14354|false|false|false|C0031046|Pericarditis|pericarditis
Disorder|Neoplastic Process|Hospital Course|14355,14364|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Finding|Functional Concept|Hospital Course|14355,14364|false|false|false|C1522484|metastatic qualifier|Secondary
Attribute|Clinical Attribute|Hospital Course|14355,14374|false|false|false|C4255018||Secondary Diagnosis
Finding|Finding|Hospital Course|14355,14374|false|false|false|C0332138|Secondary diagnosis|Secondary Diagnosis
Attribute|Clinical Attribute|Hospital Course|14365,14374|false|false|false|C0945731||Diagnosis
Finding|Classification|Hospital Course|14365,14374|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|14365,14374|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|14365,14374|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Disease or Syndrome|Hospital Course|14376,14396|false|false|false|C0003873|Rheumatoid Arthritis|rheumatoid arthritis
Disorder|Disease or Syndrome|Hospital Course|14387,14396|false|false|false|C0003864|Arthritis|arthritis
Finding|Mental Process|Discharge Condition|14422,14428|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|14422,14435|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|14422,14435|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|14429,14435|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|14429,14435|false|false|false|C1546481|What subject filter - Status|Status
Finding|Idea or Concept|Discharge Condition|14437,14442|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Finding|Discharge Condition|14447,14455|false|false|false|C4068804|Coherent|coherent
Attribute|Clinical Attribute|Discharge Condition|14457,14479|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|14457,14479|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Finding|Finding|Discharge Condition|14466,14479|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|14466,14479|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|14481,14486|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|14481,14486|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|14481,14486|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|Discharge Condition|14481,14486|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|14481,14486|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|14481,14486|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|14491,14502|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|14504,14512|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|14504,14512|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|14504,14512|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|14513,14519|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|14513,14519|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|Discharge Condition|14521,14531|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|14521,14531|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|14521,14531|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|14521,14531|false|false|false|C1561560|ambulatory encounter|Ambulatory
Finding|Finding|Discharge Condition|14534,14545|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Condition|14534,14545|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Gene or Genome|Discharge Instructions|14574,14578|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Finding|Idea or Concept|Discharge Instructions|14621,14629|false|false|false|C1547192|Organization unit type - Hospital|HOSPITAL
Finding|Idea or Concept|Discharge Instructions|14660,14668|false|false|false|C1547192|Organization unit type - Hospital|hospital
Anatomy|Body Location or Region|Discharge Instructions|14674,14679|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Discharge Instructions|14674,14679|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Discharge Instructions|14674,14684|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Discharge Instructions|14674,14684|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Discharge Instructions|14680,14684|false|false|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|14680,14684|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|14680,14684|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Idea or Concept|Discharge Instructions|14725,14733|false|false|false|C1547192|Organization unit type - Hospital|HOSPITAL
Finding|Pathologic Function|Discharge Instructions|14763,14775|false|false|false|C0021368|Inflammation|inflammation
Finding|Conceptual Entity|Discharge Instructions|14782,14787|false|false|false|C1707059|Pre-Release Version|build
Drug|Substance|Discharge Instructions|14794,14799|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Discharge Instructions|14794,14799|false|false|false|C1546638|Fluid Specimen Code|fluid
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|14822,14827|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|14822,14827|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Discharge Instructions|14822,14827|false|false|false|C0795691|HEART PROBLEM|heart
Attribute|Clinical Attribute|Discharge Instructions|14841,14850|false|false|false|C0945766||procedure
Event|Occupational Activity|Discharge Instructions|14841,14850|false|false|false|C1546467|Act Class - procedure|procedure
Finding|Functional Concept|Discharge Instructions|14841,14850|false|false|false|C2700391|Procedure (set of actions)|procedure
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|14841,14850|false|false|false|C0184661|Interventional procedure|procedure
Drug|Substance|Discharge Instructions|14865,14870|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Discharge Instructions|14865,14870|false|false|false|C1546638|Fluid Specimen Code|fluid
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|14895,14900|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|14895,14900|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Discharge Instructions|14895,14900|false|false|false|C0795691|HEART PROBLEM|heart
Finding|Idea or Concept|Discharge Instructions|14907,14916|false|false|false|C1548539;C3245481|EntityNameUseR2 - temporary;Job Status - Temporary|temporary
Finding|Intellectual Product|Discharge Instructions|14907,14916|false|false|false|C1548539;C3245481|EntityNameUseR2 - temporary;Job Status - Temporary|temporary
Drug|Substance|Discharge Instructions|14917,14922|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|Discharge Instructions|14917,14922|false|false|false|C1546604|Drain Specimen Code|drain
Finding|Idea or Concept|Discharge Instructions|14969,14977|false|false|false|C1547192|Organization unit type - Hospital|hospital
Drug|Pharmacologic Substance|Discharge Instructions|14995,15005|false|false|false|C0013227|Pharmaceutical Preparations|medication
Finding|Intellectual Product|Discharge Instructions|14995,15005|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Finding|Pathologic Function|Discharge Instructions|15030,15042|false|false|false|C0013604;C0546817|Edema;Hypervolemia (finding)|excess fluid
Drug|Substance|Discharge Instructions|15037,15042|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Discharge Instructions|15037,15042|false|false|false|C1546638|Fluid Specimen Code|fluid
Anatomy|Anatomical Structure|Discharge Instructions|15052,15056|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|15052,15056|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Finding|Intellectual Product|Discharge Instructions|15052,15056|false|false|false|C1551342|Document Body|body
Finding|Finding|Discharge Instructions|15078,15086|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Finding|Idea or Concept|Discharge Instructions|15078,15086|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|15087,15092|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|15087,15092|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Discharge Instructions|15087,15092|false|false|false|C0795691|HEART PROBLEM|heart
Finding|Organ or Tissue Function|Discharge Instructions|15087,15099|false|false|false|C0232187|Cardiac rhythm type|heart rhythm
Finding|Finding|Discharge Instructions|15093,15099|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|Discharge Instructions|15093,15099|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Disorder|Disease or Syndrome|Discharge Instructions|15101,15105|false|false|false|C0004238|Atrial Fibrillation|afib
Lab|Laboratory or Test Result|Discharge Instructions|15101,15105|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|afib
Finding|Idea or Concept|Discharge Instructions|15121,15129|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Finding|Discharge Instructions|15153,15156|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Discharge Instructions|15153,15156|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Drug|Pharmacologic Substance|Discharge Instructions|15157,15167|false|false|false|C0013227|Pharmaceutical Preparations|medication
Finding|Intellectual Product|Discharge Instructions|15157,15167|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Drug|Organic Chemical|Discharge Instructions|15179,15189|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|Discharge Instructions|15179,15189|false|false|false|C0025859|metoprolol|metoprolol
Disorder|Disease or Syndrome|Discharge Instructions|15218,15226|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|diabetes
Procedure|Health Care Activity|Discharge Instructions|15239,15248|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Finding|Discharge Instructions|15273,15276|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Discharge Instructions|15273,15276|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Drug|Pharmacologic Substance|Discharge Instructions|15277,15287|false|false|false|C0013227|Pharmaceutical Preparations|medication
Finding|Intellectual Product|Discharge Instructions|15277,15287|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Drug|Organic Chemical|Discharge Instructions|15298,15307|false|false|false|C0025598|metformin|metformin
Drug|Pharmacologic Substance|Discharge Instructions|15298,15307|false|false|false|C0025598|metformin|metformin
Finding|Functional Concept|Discharge Instructions|15325,15329|false|false|false|C0686904|Patient need for (contextual qualifier)|NEED
Finding|Idea or Concept|Discharge Instructions|15355,15363|false|false|false|C1547192|Organization unit type - Hospital|HOSPITAL
Attribute|Clinical Attribute|Discharge Instructions|15386,15397|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|15386,15397|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|Discharge Instructions|15386,15397|false|false|false|C4284232|Medications|medications
Finding|Functional Concept|Discharge Instructions|15431,15437|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|Follow
Finding|Intellectual Product|Discharge Instructions|15431,15437|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|Follow
Finding|Finding|Discharge Instructions|15431,15440|false|false|false|C0589120|Follow-up status|Follow up
Procedure|Health Care Activity|Discharge Instructions|15431,15440|false|false|false|C1522577|follow-up|Follow up
Finding|Functional Concept|Discharge Instructions|15514,15521|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|Discharge Instructions|15514,15521|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|Discharge Instructions|15514,15521|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|Discharge Instructions|15514,15521|false|false|false|C0199168|Medical service|medical
Finding|Intellectual Product|Discharge Instructions|15522,15531|false|false|false|C0004268;C4281780|Attention;Attention - G-code|attention
Finding|Mental Process|Discharge Instructions|15522,15531|false|false|false|C0004268;C4281780|Attention;Attention - G-code|attention
Attribute|Clinical Attribute|Discharge Instructions|15541,15547|false|false|false|C0944911||weight
Finding|Finding|Discharge Instructions|15541,15547|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|Discharge Instructions|15541,15547|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|Discharge Instructions|15541,15547|false|false|false|C1305866|Weighing patient|weight
Procedure|Laboratory Procedure|Discharge Instructions|15568,15571|false|false|false|C3161851|liquid-based cytology (procedure)|lbs
Finding|Intellectual Product|Discharge Instructions|15577,15581|false|false|false|C5239649|PANEL.SURVEY.SEEK|Seek
Finding|Functional Concept|Discharge Instructions|15582,15589|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|Discharge Instructions|15582,15589|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|Discharge Instructions|15582,15589|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|Discharge Instructions|15582,15589|false|false|false|C0199168|Medical service|medical
Finding|Intellectual Product|Discharge Instructions|15590,15599|false|false|false|C0004268;C4281780|Attention;Attention - G-code|attention
Finding|Mental Process|Discharge Instructions|15590,15599|false|false|false|C0004268;C4281780|Attention;Attention - G-code|attention
Finding|Finding|Discharge Instructions|15612,15615|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Discharge Instructions|15612,15615|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Functional Concept|Discharge Instructions|15630,15638|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Discharge Instructions|15630,15638|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Finding|Discharge Instructions|15655,15663|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|Discharge Instructions|15655,15663|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|15672,15676|false|false|false|C1140621|Leg|legs
Attribute|Clinical Attribute|Discharge Instructions|15672,15676|false|false|false|C5781420||legs
Anatomy|Body Location or Region|Discharge Instructions|15678,15687|false|false|false|C0000726|Abdomen|abdominal
Finding|Finding|Discharge Instructions|15678,15698|false|false|false|C0000731|Abdomen distended|abdominal distention
Finding|Finding|Discharge Instructions|15688,15698|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Finding|Pathologic Function|Discharge Instructions|15688,15698|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Attribute|Clinical Attribute|Discharge Instructions|15704,15723|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|Discharge Instructions|15704,15723|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|Discharge Instructions|15717,15723|false|false|false|C0225386|Breath|breath
Finding|Idea or Concept|Discharge Instructions|15763,15774|false|false|false|C0870705;C1533716;C1561527;C1561528|Acknowledgement Detail Type - Information;Error severity - Information;Information;control act - information|information
Finding|Intellectual Product|Discharge Instructions|15763,15774|false|false|false|C0870705;C1533716;C1561527;C1561528|Acknowledgement Detail Type - Information;Error severity - Information;Information;control act - information|information
Procedure|Health Care Activity|Discharge Instructions|15783,15798|false|false|false|C0019993|Hospitalization|hospitalization
Finding|Intellectual Product|Discharge Instructions|15810,15818|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|Discharge Instructions|15810,15818|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Idea or Concept|Discharge Instructions|15826,15830|false|false|false|C1552020|Role Class - part|part
Event|Activity|Discharge Instructions|15839,15843|false|false|false|C1947933|care activity|care
Finding|Finding|Discharge Instructions|15839,15843|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|15839,15843|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Disorder|Disease or Syndrome|Discharge Instructions|15880,15884|false|false|false|C0339510|Vitelliform Macular Dystrophy|best
Finding|Gene or Genome|Discharge Instructions|15880,15884|false|false|false|C1826421;C5781213|BEST1 gene;BEST1 wt Allele|best
Event|Activity|Discharge Instructions|15900,15904|false|false|false|C1947933|care activity|Care
Finding|Finding|Discharge Instructions|15900,15904|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Discharge Instructions|15900,15904|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Attribute|Clinical Attribute|Discharge Instructions|15900,15909|false|false|false|C4321316||Care Team
Finding|Finding|Discharge Instructions|15900,15909|false|false|false|C4321315|Care team|Care Team
Procedure|Health Care Activity|Discharge Instructions|15914,15922|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|15923,15935|false|false|false|C3263700||Instructions
Finding|Intellectual Product|Discharge Instructions|15923,15935|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

