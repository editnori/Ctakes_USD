 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|39,48|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|39,48|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|39,53|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|73,82|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|73,82|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|73,82|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|73,82|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|73,82|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|73,87|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|105,110|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|105,110|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|105,110|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|129,132|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|140,147|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|140,147|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|149,157|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|Allergies|181,190|false|false|false|C1717415||Allergies
Event|Event|Allergies|181,190|false|false|false|||Allergies
Finding|Pathologic Function|Allergies|181,190|false|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|Allergies|193,215|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|Allergies|201,205|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|Allergies|201,205|false|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|Allergies|201,215|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Event|Event|Allergies|206,215|false|false|false|||Reactions
Event|Event|Allergies|218,227|false|false|false|||Attending
Finding|Functional Concept|Allergies|218,227|false|false|false|C1999232|Attending (action)|Attending
Event|Event|Chief Complaint|253,260|false|false|false|||Dyspnea
Finding|Finding|Chief Complaint|253,260|false|false|false|C0013404;C2024878|Dyspnea|Dyspnea
Finding|Sign or Symptom|Chief Complaint|253,260|false|false|false|C0013404;C2024878|Dyspnea|Dyspnea
Anatomy|Body Location or Region|Chief Complaint|265,270|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Chief Complaint|265,270|false|false|false|C0741025|Chest problem|chest
Finding|Sign or Symptom|Chief Complaint|265,280|false|false|false|C0232292|Chest tightness|chest tightness
Event|Event|Chief Complaint|271,280|false|false|false|||tightness
Finding|Classification|Chief Complaint|283,288|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|289,297|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|289,297|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|301,319|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|310,319|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|310,319|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|310,319|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|310,319|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|310,319|false|false|false|C0184661|Interventional procedure|Procedure
Finding|Functional Concept|Chief Complaint|325,338|false|false|false|C0205464|pharmacological|Pharmacologic
Procedure|Diagnostic Procedure|Chief Complaint|339,358|false|false|false|C2825165|Nuclear stress test|nuclear stress test
Attribute|Clinical Attribute|Chief Complaint|347,353|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|Chief Complaint|347,353|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|Chief Complaint|347,353|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Finding|Finding|Chief Complaint|347,353|false|false|false|C0038435|Stress|stress
Procedure|Diagnostic Procedure|Chief Complaint|347,358|false|false|false|C0015260;C3494508|Exercise stress test;Stress Test|stress test
Anatomy|Body Location or Region|Chief Complaint|354,358|false|false|false|C4318744|Test - temporal region|test
Event|Event|Chief Complaint|354,358|false|false|false|||test
Finding|Functional Concept|Chief Complaint|354,358|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|Chief Complaint|354,358|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|Chief Complaint|354,358|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|Chief Complaint|354,358|false|false|false|C0022885|Laboratory Procedures|test
Finding|Idea or Concept|History of Present Illness|393,397|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|History of Present Illness|393,397|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|History of Present Illness|398,401|false|false|false|||old
Event|Event|History of Present Illness|414,421|false|false|false|||history
Finding|Conceptual Entity|History of Present Illness|414,421|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|414,421|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|414,421|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|414,424|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|History of Present Illness|425,428|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|History of Present Illness|425,428|false|false|false|||HTN
Event|Event|History of Present Illness|430,433|false|false|false|||HLD
Disorder|Disease or Syndrome|History of Present Illness|441,444|false|false|false|C0001365;C0038454|Acute ill-defined cerebrovascular disease;Cerebrovascular accident|CVA
Drug|Pharmacologic Substance|History of Present Illness|441,444|false|false|false|C5779650|Cyclophosphamide/Doxorubicin/Vincristine|CVA
Event|Event|History of Present Illness|441,444|false|false|false|||CVA
Disorder|Disease or Syndrome|History of Present Illness|446,449|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|446,449|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|History of Present Illness|446,449|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|History of Present Illness|446,449|false|false|false|||CAD
Finding|Gene or Genome|History of Present Illness|446,449|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|History of Present Illness|446,449|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|History of Present Illness|446,449|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|446,449|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|History of Present Illness|455,458|false|false|false|C0006430|Burning Mouth Syndrome|BMS
Event|Event|History of Present Illness|455,458|false|false|false|||BMS
Event|Event|History of Present Illness|462,472|false|false|false|||circumflex
Event|Event|History of Present Illness|477,481|false|false|false|||POBA
Drug|Organic Chemical|History of Present Illness|492,499|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|History of Present Illness|492,499|false|false|false|C0004057|aspirin|Aspirin
Event|Event|History of Present Illness|492,499|false|false|false|||Aspirin
Drug|Organic Chemical|History of Present Illness|504,510|false|false|false|C0633084|Plavix|Plavix
Drug|Pharmacologic Substance|History of Present Illness|504,510|false|false|false|C0633084|Plavix|Plavix
Event|Event|History of Present Illness|504,510|false|false|false|||Plavix
Anatomy|Body Space or Junction|History of Present Illness|512,515|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|History of Present Illness|512,515|false|false|false|C0018802|Congestive heart failure|CHF
Event|Event|History of Present Illness|512,515|false|false|false|||CHF
Disorder|Disease or Syndrome|History of Present Illness|533,541|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|diabetes
Event|Event|History of Present Illness|533,541|false|false|false|||diabetes
Event|Event|History of Present Illness|543,553|false|false|false|||presenting
Finding|Intellectual Product|History of Present Illness|559,564|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Intellectual Product|History of Present Illness|559,570|false|false|false|C1272517|Sudden onset (contextual qualifier) (qualifier value)|acute onset
Event|Event|History of Present Illness|565,570|false|false|false|||onset
Event|Event|History of Present Illness|572,581|false|false|false|||shortness
Attribute|Clinical Attribute|History of Present Illness|572,591|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|History of Present Illness|572,591|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|History of Present Illness|585,591|false|false|false|C0225386|Breath|breath
Anatomy|Body Location or Region|History of Present Illness|607,612|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|607,612|false|false|false|C0741025|Chest problem|chest
Finding|Sign or Symptom|History of Present Illness|607,622|false|false|false|C0232292|Chest tightness|chest tightness
Event|Event|History of Present Illness|613,622|false|false|false|||tightness
Event|Event|History of Present Illness|634,641|false|false|false|||evening
Finding|Body Substance|History of Present Illness|645,652|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|645,652|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|645,652|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|History of Present Illness|653,658|false|false|false|||notes
Finding|Gene or Genome|History of Present Illness|682,687|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Drug|Food|History of Present Illness|688,695|false|false|false|C0206208|Seafood|seafood
Event|Event|History of Present Illness|696,702|false|false|false|||dinner
Finding|Daily or Recreational Activity|History of Present Illness|696,702|false|false|false|C4048877|Dinner|dinner
Event|Event|History of Present Illness|717,722|false|false|false|||usual
Finding|Intellectual Product|History of Present Illness|736,740|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|History of Present Illness|763,768|false|false|false|||acute
Finding|Intellectual Product|History of Present Illness|763,768|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|History of Present Illness|770,775|false|false|false|||onset
Finding|Sign or Symptom|History of Present Illness|779,782|false|false|false|C0013404|Dyspnea|SOB
Event|Event|History of Present Illness|783,790|false|false|false|||feeling
Finding|Mental Process|History of Present Illness|783,790|false|false|false|C1527305|Feelings|feeling
Event|Event|History of Present Illness|810,814|false|false|false|||take
Attribute|Clinical Attribute|History of Present Illness|815,819|false|true|false|C4318566|Deep Resection Margin|deep
Event|Event|History of Present Illness|820,827|false|false|false|||breaths
Finding|Body Substance|History of Present Illness|820,827|false|true|false|C0225386|Breath|breaths
Anatomy|Body Location or Region|History of Present Illness|834,839|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|834,839|false|false|false|C0741025|Chest problem|chest
Finding|Sign or Symptom|History of Present Illness|834,849|false|false|false|C0232292|Chest tightness|chest tightness
Event|Event|History of Present Illness|840,849|false|false|false|||tightness
Finding|Body Substance|History of Present Illness|851,858|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|851,858|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|851,858|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|859,864|false|false|false|||notes
Attribute|Clinical Attribute|History of Present Illness|878,884|false|false|false|C2926611||angina
Event|Event|History of Present Illness|878,884|false|false|false|||angina
Finding|Finding|History of Present Illness|878,884|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Finding|Sign or Symptom|History of Present Illness|878,884|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Event|Event|History of Present Illness|888,894|false|false|false|||Denies
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|906,915|false|false|false|C1179435|Protein Component|component
Drug|Biologically Active Substance|History of Present Illness|906,915|false|false|false|C1179435|Protein Component|component
Event|Event|History of Present Illness|906,915|false|false|false|||component
Finding|Conceptual Entity|History of Present Illness|906,915|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Idea or Concept|History of Present Illness|906,915|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Intellectual Product|History of Present Illness|906,915|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Event|Event|History of Present Illness|923,932|false|false|false|||described
Drug|Pharmacologic Substance|History of Present Illness|936,943|false|false|false|C0719205|Central brand of multivitamin with minerals|central
Drug|Vitamin|History of Present Illness|936,943|false|false|false|C0719205|Central brand of multivitamin with minerals|central
Event|Event|History of Present Illness|936,943|false|false|false|||central
Procedure|Laboratory Procedure|History of Present Illness|936,943|false|false|false|C1879652|Central Minus|central
Anatomy|Body Location or Region|History of Present Illness|955,960|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|History of Present Illness|955,960|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|962,965|false|false|false|C0035561|Bone structure of rib|rib
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|962,970|false|false|false|C0222762|Rib Cage|rib cage
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|966,970|false|false|false|C4555210|CAGE Antibody|cage
Drug|Immunologic Factor|History of Present Illness|966,970|false|false|false|C4555210|CAGE Antibody|cage
Drug|Pharmacologic Substance|History of Present Illness|966,970|false|false|false|C4555210|CAGE Antibody|cage
Event|Event|History of Present Illness|966,970|false|false|false|||cage
Finding|Gene or Genome|History of Present Illness|966,970|false|false|false|C1426669|DDX53 gene|cage
Procedure|Laboratory Procedure|History of Present Illness|966,970|false|false|false|C5552712|CAP Analysis of Gene Expression|cage
Event|Event|History of Present Illness|972,982|false|false|false|||persistent
Event|Event|History of Present Illness|989,994|false|false|false|||onset
Event|Event|History of Present Illness|999,1008|false|false|false|||radiation
Phenomenon|Natural Phenomenon or Process|History of Present Illness|999,1008|true|false|false|C0034519;C0851346|Electromagnetic Radiation;Radiation|radiation
Procedure|Research Activity|History of Present Illness|999,1008|true|false|false|C1522449;C1524020;C1524021|Radiation Ionizing Radiotherapy;Radiation therapy (procedure);Radiotherapy Research|radiation
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|999,1008|true|false|false|C1522449;C1524020;C1524021|Radiation Ionizing Radiotherapy;Radiation therapy (procedure);Radiotherapy Research|radiation
Anatomy|Body Location or Region|History of Present Illness|1017,1026|false|false|false|C0037004|Shoulder|shoulders
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1027,1030|false|false|false|C0022359|Jaw|jaw
Event|Event|History of Present Illness|1040,1051|false|false|false|||diaphoreses
Event|Event|History of Present Illness|1053,1060|false|false|false|||Worsens
Event|Activity|History of Present Illness|1066,1074|false|false|false|C0441655|Activities|activity
Event|Event|History of Present Illness|1066,1074|false|false|false|||activity
Finding|Daily or Recreational Activity|History of Present Illness|1066,1074|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Finding|Finding|History of Present Illness|1066,1074|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Event|Event|History of Present Illness|1077,1085|false|false|false|||improves
Finding|Finding|History of Present Illness|1086,1094|false|false|false|C2984079|Somewhat|somewhat
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1100,1104|false|false|false|C1742913|REST protein, human|rest
Drug|Biologically Active Substance|History of Present Illness|1100,1104|false|false|false|C1742913|REST protein, human|rest
Event|Event|History of Present Illness|1100,1104|false|false|false|||rest
Finding|Daily or Recreational Activity|History of Present Illness|1100,1104|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Gene or Genome|History of Present Illness|1100,1104|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Molecular Function|History of Present Illness|1100,1104|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Body Substance|History of Present Illness|1106,1113|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|1106,1113|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|1106,1113|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|History of Present Illness|1126,1131|false|false|false|||feels
Event|Event|History of Present Illness|1144,1152|false|false|false|||episodes
Finding|Intellectual Product|History of Present Illness|1162,1166|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|History of Present Illness|1167,1175|false|false|false|||required
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1180,1195|false|false|false|C2348535|Stenting|stent placement
Event|Event|History of Present Illness|1186,1195|false|false|false|||placement
Procedure|Health Care Activity|History of Present Illness|1186,1195|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1186,1195|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Event|Event|History of Present Illness|1218,1226|false|false|false|||improved
Event|Event|History of Present Illness|1231,1239|false|false|false|||symptoms
Finding|Functional Concept|History of Present Illness|1231,1239|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|History of Present Illness|1231,1239|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|History of Present Illness|1253,1262|false|false|false|||persisted
Event|Event|History of Present Illness|1288,1291|false|false|false|||led
Anatomy|Body Location or Region|History of Present Illness|1295,1304|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|History of Present Illness|1295,1315|false|false|false|C0232487|Abdominal discomfort|abdominal discomfort
Event|Event|History of Present Illness|1305,1315|false|false|false|||discomfort
Finding|Sign or Symptom|History of Present Illness|1305,1315|false|false|false|C2364135|Discomfort|discomfort
Event|Event|History of Present Illness|1321,1329|false|false|false|||vomiting
Finding|Sign or Symptom|History of Present Illness|1321,1329|false|false|false|C0042963|Vomiting|vomiting
Event|Event|History of Present Illness|1335,1344|false|false|false|||nonbloody
Finding|Daily or Recreational Activity|History of Present Illness|1350,1356|false|false|false|C4048877|Dinner|dinner
Event|Event|History of Present Illness|1357,1363|false|false|false|||pieces
Event|Event|History of Present Illness|1367,1368|false|false|false|||_
Finding|Idea or Concept|History of Present Illness|1372,1375|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|History of Present Illness|1372,1375|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|History of Present Illness|1385,1394|false|false|false|||admission
Procedure|Health Care Activity|History of Present Illness|1385,1394|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|History of Present Illness|1397,1404|false|false|false|||decided
Event|Event|History of Present Illness|1408,1411|false|false|false|||see
Attribute|Clinical Attribute|History of Present Illness|1419,1423|false|false|false|C2598155||pain
Event|Event|History of Present Illness|1419,1423|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|1419,1423|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1419,1423|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|1424,1432|false|false|false|||improved
Finding|Finding|History of Present Illness|1440,1443|false|false|false|C5939094|Own|own
Finding|Intellectual Product|History of Present Illness|1445,1449|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|History of Present Illness|1459,1468|false|false|false|||persisted
Event|Event|History of Present Illness|1485,1493|false|false|false|||arranged
Drug|Biologically Active Substance|History of Present Illness|1501,1505|false|false|false|C0245203|4-azido-7-phenylpyrazolo-(1,5a)-1,3,5-triazine|appt
Drug|Organic Chemical|History of Present Illness|1501,1505|false|false|false|C0245203|4-azido-7-phenylpyrazolo-(1,5a)-1,3,5-triazine|appt
Event|Event|History of Present Illness|1501,1505|false|false|false|||appt
Disorder|Disease or Syndrome|History of Present Illness|1522,1525|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|1522,1525|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|History of Present Illness|1522,1525|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1522,1525|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|History of Present Illness|1522,1525|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|History of Present Illness|1522,1525|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|History of Present Illness|1522,1525|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|History of Present Illness|1522,1525|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|History of Present Illness|1522,1525|false|false|false|||PCP
Finding|Gene or Genome|History of Present Illness|1522,1525|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|History of Present Illness|1522,1525|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Attribute|Clinical Attribute|History of Present Illness|1532,1535|false|false|false|C0871470|Systolic Pressure|SBP
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1532,1535|false|false|false|C0085805|Androgen Binding Protein|SBP
Drug|Biologically Active Substance|History of Present Illness|1532,1535|false|false|false|C0085805|Androgen Binding Protein|SBP
Event|Event|History of Present Illness|1532,1535|false|false|false|||SBP
Finding|Gene or Genome|History of Present Illness|1532,1535|false|false|false|C1705296;C3274833|CCHCR1 wt Allele;SHBG wt Allele|SBP
Procedure|Diagnostic Procedure|History of Present Illness|1532,1535|false|false|false|C1306620|Systolic blood pressure measurement|SBP
Event|Event|History of Present Illness|1548,1551|false|false|false|||EKG
Finding|Intellectual Product|History of Present Illness|1548,1551|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|History of Present Illness|1548,1551|false|false|false|C1623258|Electrocardiography|EKG
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|1561,1572|false|false|false|C0011570|Mental Depression|depressions
Event|Event|History of Present Illness|1561,1572|false|false|false|||depressions
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1643,1646|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Enzyme|History of Present Illness|1643,1646|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Organic Chemical|History of Present Illness|1643,1646|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Pharmacologic Substance|History of Present Illness|1643,1646|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Event|Event|History of Present Illness|1643,1646|false|false|false|||ASA
Finding|Gene or Genome|History of Present Illness|1643,1646|false|false|false|C1412553|ARSA gene|ASA
Event|Event|History of Present Illness|1662,1666|false|false|false|||sent
Finding|Functional Concept|History of Present Illness|1662,1666|false|false|false|C1519246|Send (transmission)|sent
Event|Event|History of Present Illness|1683,1690|false|false|false|||concern
Finding|Idea or Concept|History of Present Illness|1683,1690|false|false|false|C2699424|Concern|concern
Anatomy|Body Space or Junction|History of Present Illness|1696,1699|false|false|false|C0262187|anterior calcarine sulcus (human only)|ACS
Disorder|Disease or Syndrome|History of Present Illness|1696,1699|false|false|false|C0742343;C0796147|Acrocallosal Syndrome;Acute Chest Syndrome|ACS
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1696,1699|false|false|false|C4042561|ACSS2 protein, human|ACS
Drug|Enzyme|History of Present Illness|1696,1699|false|false|false|C4042561|ACSS2 protein, human|ACS
Event|Event|History of Present Illness|1696,1699|false|false|false|||ACS
Finding|Gene or Genome|History of Present Illness|1696,1699|false|false|false|C1150760;C1424787;C1825842;C1842089;C2266615;C4318612;C5400867;C5551036|ACCS gene;ACS - Activity Card Sort;ACSS2 gene;ACSS2 wt Allele;American Community Survey;CO-methylating acetyl-CoA synthase activity;PLA2G15 gene;acetate-CoA ligase activity|ACS
Finding|Intellectual Product|History of Present Illness|1696,1699|false|false|false|C1150760;C1424787;C1825842;C1842089;C2266615;C4318612;C5400867;C5551036|ACCS gene;ACS - Activity Card Sort;ACSS2 gene;ACSS2 wt Allele;American Community Survey;CO-methylating acetyl-CoA synthase activity;PLA2G15 gene;acetate-CoA ligase activity|ACS
Finding|Molecular Function|History of Present Illness|1696,1699|false|false|false|C1150760;C1424787;C1825842;C1842089;C2266615;C4318612;C5400867;C5551036|ACCS gene;ACS - Activity Card Sort;ACSS2 gene;ACSS2 wt Allele;American Community Survey;CO-methylating acetyl-CoA synthase activity;PLA2G15 gene;acetate-CoA ligase activity|ACS
Disorder|Disease or Syndrome|History of Present Illness|1707,1710|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|History of Present Illness|1707,1710|false|false|false|||HTN
Event|Event|History of Present Illness|1711,1720|false|false|false|||emergency
Finding|Finding|History of Present Illness|1711,1720|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Idea or Concept|History of Present Illness|1711,1720|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Intellectual Product|History of Present Illness|1711,1720|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Pathologic Function|History of Present Illness|1711,1720|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Phenomenon|Phenomenon or Process|History of Present Illness|1711,1720|false|false|false|C0013956|Emergency Situation|emergency
Procedure|Health Care Activity|History of Present Illness|1711,1720|false|false|false|C1553500|emergency encounter|emergency
Finding|Body Substance|History of Present Illness|1724,1731|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|1724,1731|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|1724,1731|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|History of Present Illness|1732,1741|false|false|false|||reporting
Drug|Biomedical or Dental Material|History of Present Illness|1742,1750|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|History of Present Illness|1742,1750|false|false|false|||baseline
Finding|Idea or Concept|History of Present Illness|1742,1750|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|History of Present Illness|1751,1757|false|false|false|||sleeps
Event|Event|History of Present Illness|1774,1783|false|false|false|||unchanged
Finding|Finding|History of Present Illness|1774,1783|false|false|false|C0442739||unchanged
Drug|Organic Chemical|History of Present Illness|1798,1803|true|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|1798,1803|true|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|History of Present Illness|1798,1803|false|false|false|||cough
Finding|Sign or Symptom|History of Present Illness|1798,1803|true|false|false|C0010200|Coughing|cough
Disorder|Disease or Syndrome|History of Present Illness|1805,1808|true|false|false|C1956415|Paroxysmal nocturnal dyspnea|PND
Event|Event|History of Present Illness|1805,1808|false|false|false|||PND
Finding|Gene or Genome|History of Present Illness|1805,1808|true|false|false|C1417807;C4552608|NPPA gene;NPPA wt Allele|PND
Event|Event|History of Present Illness|1810,1819|false|false|false|||orthopnea
Finding|Finding|History of Present Illness|1810,1819|true|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Finding|Sign or Symptom|History of Present Illness|1810,1819|true|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Event|Event|History of Present Illness|1827,1834|false|false|false|||pillows
Finding|Idea or Concept|History of Present Illness|1836,1845|false|false|false|C1546960|Patient Outcome - Worsening|Worsening
Event|Event|History of Present Illness|1846,1849|false|false|false|||DOE
Finding|Sign or Symptom|History of Present Illness|1846,1849|false|false|false|C0231807|Dyspnea on exertion|DOE
Event|Event|History of Present Illness|1866,1874|false|false|false|||symptoms
Finding|Functional Concept|History of Present Illness|1866,1874|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|History of Present Illness|1866,1874|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|History of Present Illness|1880,1886|false|false|false|||unable
Finding|Finding|History of Present Illness|1880,1886|false|false|false|C1299582|Unable|unable
Finding|Finding|History of Present Illness|1880,1898|false|false|false|C3842772|Unable to complete|unable to complete
Event|Event|History of Present Illness|1890,1898|false|false|false|||complete
Drug|Biomedical or Dental Material|History of Present Illness|1901,1906|false|false|false|C1706085|Block Dosage Form|block
Event|Event|History of Present Illness|1901,1906|false|false|false|||block
Finding|Body Substance|History of Present Illness|1901,1906|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|block
Finding|Finding|History of Present Illness|1901,1906|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|block
Finding|Functional Concept|History of Present Illness|1901,1906|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|block
Event|Event|History of Present Illness|1918,1922|false|false|false|||used
Event|Event|History of Present Illness|1929,1933|false|false|false|||able
Finding|Finding|History of Present Illness|1929,1933|false|false|false|C1299581|Able (qualifier value)|able
Event|Event|History of Present Illness|1937,1941|false|false|false|||walk
Event|Event|History of Present Illness|1948,1954|false|false|false|||blocks
Finding|Body Substance|History of Present Illness|1948,1954|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|blocks
Finding|Finding|History of Present Illness|1948,1954|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|blocks
Finding|Functional Concept|History of Present Illness|1948,1954|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|blocks
Finding|Finding|History of Present Illness|1960,1964|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|History of Present Illness|1960,1964|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|History of Present Illness|1960,1964|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|History of Present Illness|1974,1982|false|false|false|||stopping
Event|Event|History of Present Illness|1987,1990|false|false|false|||SOB
Finding|Sign or Symptom|History of Present Illness|1987,1990|false|false|false|C0013404|Dyspnea|SOB
Event|Event|History of Present Illness|1995,2001|false|false|false|||Denies
Finding|Finding|History of Present Illness|2002,2005|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|History of Present Illness|2002,2005|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Attribute|Clinical Attribute|History of Present Illness|2010,2015|false|false|false|C1717255||edema
Event|Event|History of Present Illness|2010,2015|false|false|false|||edema
Finding|Pathologic Function|History of Present Illness|2010,2015|false|false|false|C0013604|Edema|edema
Drug|Biomedical or Dental Material|History of Present Illness|2017,2025|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|History of Present Illness|2017,2025|false|false|false|||baseline
Finding|Idea or Concept|History of Present Illness|2017,2025|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|History of Present Illness|2026,2030|false|false|false|||says
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2033,2036|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Event|Event|History of Present Illness|2054,2060|false|false|false|||emesis
Finding|Body Substance|History of Present Illness|2054,2060|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Physiologic Function|History of Present Illness|2054,2060|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Sign or Symptom|History of Present Illness|2054,2060|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Event|Event|History of Present Illness|2080,2091|false|false|false|||diaphoresis
Finding|Finding|History of Present Illness|2080,2091|true|false|false|C0700590|Increased sweating|diaphoresis
Anatomy|Body Location or Region|History of Present Illness|2096,2101|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|2096,2101|true|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|2096,2106|true|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|2096,2106|true|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|2102,2106|true|false|false|C2598155||pain
Event|Event|History of Present Illness|2102,2106|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|2102,2106|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|2102,2106|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|2112,2121|false|false|false|||radiation
Phenomenon|Natural Phenomenon or Process|History of Present Illness|2112,2121|true|false|false|C0034519;C0851346|Electromagnetic Radiation;Radiation|radiation
Procedure|Research Activity|History of Present Illness|2112,2121|true|false|false|C1522449;C1524020;C1524021|Radiation Ionizing Radiotherapy;Radiation therapy (procedure);Radiotherapy Research|radiation
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|2112,2121|true|false|false|C1522449;C1524020;C1524021|Radiation Ionizing Radiotherapy;Radiation therapy (procedure);Radiotherapy Research|radiation
Event|Event|History of Present Illness|2125,2133|false|false|false|||symptoms
Finding|Functional Concept|History of Present Illness|2125,2133|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|History of Present Illness|2125,2133|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|History of Present Illness|2147,2155|false|false|false|||diarrhea
Finding|Finding|History of Present Illness|2147,2155|true|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|History of Present Illness|2147,2155|true|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Event|Event|History of Present Illness|2159,2171|false|false|false|||constipation
Finding|Sign or Symptom|History of Present Illness|2159,2171|true|false|false|C0009806|Constipation|constipation
Event|Event|History of Present Illness|2177,2184|false|false|false|||dysuria
Finding|Sign or Symptom|History of Present Illness|2177,2184|true|false|false|C0013428|Dysuria|dysuria
Event|Event|History of Present Illness|2195,2203|false|false|false|||weakness
Finding|Sign or Symptom|History of Present Illness|2195,2203|true|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Event|Event|History of Present Illness|2204,2212|false|false|false|||numbness
Finding|Finding|History of Present Illness|2204,2212|true|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|History of Present Illness|2204,2212|true|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Anatomy|Body Space or Junction|History of Present Illness|2217,2220|false|false|false|C0262327|rostral sulcus|ROS
Drug|Biologically Active Substance|History of Present Illness|2217,2220|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Element, Ion, or Isotope|History of Present Illness|2217,2220|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Organic Chemical|History of Present Illness|2217,2220|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Pharmacologic Substance|History of Present Illness|2217,2220|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Event|Event|History of Present Illness|2217,2220|false|false|false|||ROS
Finding|Gene or Genome|History of Present Illness|2217,2220|false|false|false|C0812281;C1709820|ROS1 gene;ROS1 wt Allele|ROS
Procedure|Health Care Activity|History of Present Illness|2217,2220|false|false|false|C0489633|Review of systems (procedure)|ROS
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2240,2243|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Disorder|Disease or Syndrome|History of Present Illness|2244,2252|false|false|false|C0030554|Paresthesia|tingling
Event|Event|History of Present Illness|2244,2252|false|false|false|||tingling
Finding|Sign or Symptom|History of Present Illness|2244,2252|false|false|false|C2242996|Has tingling sensation|tingling
Event|Event|History of Present Illness|2269,2275|false|false|false|||stable
Finding|Intellectual Product|History of Present Illness|2269,2275|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|History of Present Illness|2280,2287|false|false|false|||chronic
Finding|Intellectual Product|History of Present Illness|2280,2287|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|History of Present Illness|2280,2287|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Event|Event|History of Present Illness|2293,2301|false|false|false|||diarrhea
Finding|Finding|History of Present Illness|2293,2301|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|History of Present Illness|2293,2301|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Drug|Food|History of Present Illness|2327,2334|false|false|false|C0206208|Seafood|seafood
Event|Event|History of Present Illness|2335,2341|false|false|false|||dinner
Finding|Daily or Recreational Activity|History of Present Illness|2335,2341|false|false|false|C4048877|Dinner|dinner
Disorder|Disease or Syndrome|History of Present Illness|2350,2353|false|false|false|C0006430|Burning Mouth Syndrome|BMs
Finding|Intellectual Product|History of Present Illness|2361,2365|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Idea or Concept|History of Present Illness|2380,2387|false|false|false|C1555582|Initial (abbreviation)|initial
Drug|Food|History of Present Illness|2388,2393|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|vital
Attribute|Clinical Attribute|History of Present Illness|2388,2399|false|false|false|C0488614;C0518766|Vital signs|vital signs
Procedure|Health Care Activity|History of Present Illness|2388,2399|false|false|false|C0150404|Taking vital signs|vital signs
Event|Event|History of Present Illness|2394,2399|false|false|false|||signs
Finding|Finding|History of Present Illness|2394,2399|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|History of Present Illness|2394,2399|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|2430,2433|false|false|false|C2744672|SAT1 protein, human|Sat
Drug|Enzyme|History of Present Illness|2430,2433|false|false|false|C2744672|SAT1 protein, human|Sat
Event|Event|History of Present Illness|2430,2433|false|false|false|||Sat
Finding|Gene or Genome|History of Present Illness|2430,2433|false|false|false|C0871290;C1705827;C1822614|College Entrance Examination Board Scholastic Aptitude Test;SAT1 gene;SAT1 wt Allele|Sat
Finding|Intellectual Product|History of Present Illness|2430,2433|false|false|false|C0871290;C1705827;C1822614|College Entrance Examination Board Scholastic Aptitude Test;SAT1 gene;SAT1 wt Allele|Sat
Event|Event|History of Present Illness|2439,2441|false|false|false|||3L
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2442,2447|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|History of Present Illness|2442,2447|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|History of Present Illness|2442,2447|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|History of Present Illness|2442,2447|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|History of Present Illness|2442,2447|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|History of Present Illness|2442,2447|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2448,2455|false|false|false|C1550232|Body Parts - Cannula|cannula
Finding|Body Substance|History of Present Illness|2448,2455|false|false|false|C1546577;C1550622|Specimen Type - Cannula|cannula
Finding|Intellectual Product|History of Present Illness|2448,2455|false|false|false|C1546577;C1550622|Specimen Type - Cannula|cannula
Lab|Laboratory or Test Result|History of Present Illness|2457,2461|false|false|false|C0587081|Laboratory test finding|Labs
Event|Event|History of Present Illness|2462,2469|false|false|false|||notable
Drug|Biomedical or Dental Material|History of Present Illness|2482,2490|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|History of Present Illness|2482,2490|false|false|false|||baseline
Finding|Idea or Concept|History of Present Illness|2482,2490|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Drug|Biologically Active Substance|History of Present Illness|2502,2505|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Drug|Inorganic Chemical|History of Present Illness|2502,2505|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Event|Event|History of Present Illness|2502,2505|false|false|false|||BUN
Procedure|Laboratory Procedure|History of Present Illness|2502,2505|false|false|false|C0005845|Blood urea nitrogen measurement|BUN
Anatomy|Cell|History of Present Illness|2510,2513|false|false|false|C0023516|Leukocytes|wbc
Event|Event|History of Present Illness|2533,2536|false|false|false|||Plt
Procedure|Laboratory Procedure|History of Present Illness|2533,2536|false|false|false|C0201617|Primed lymphocyte test|Plt
Finding|Idea or Concept|History of Present Illness|2542,2549|false|false|false|C1555582|Initial (abbreviation)|Initial
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|2569,2572|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Hormone|History of Present Illness|2569,2572|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Pharmacologic Substance|History of Present Illness|2569,2572|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Event|Event|History of Present Illness|2569,2572|false|false|false|||BNP
Finding|Gene or Genome|History of Present Illness|2569,2572|false|false|false|C1417808;C2982014|NPPB gene;NPPB wt Allele|BNP
Procedure|Laboratory Procedure|History of Present Illness|2569,2572|false|false|false|C1095989|Brain natriuretic peptide measurement|BNP
Event|Event|History of Present Illness|2579,2582|false|false|false|||CXR
Procedure|Diagnostic Procedure|History of Present Illness|2579,2582|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|History of Present Illness|2583,2589|false|false|false|||showed
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2593,2602|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|History of Present Illness|2593,2602|false|false|false|C2707265||pulmonary
Finding|Finding|History of Present Illness|2593,2602|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|History of Present Illness|2593,2608|true|false|false|C0034063|Pulmonary Edema|pulmonary edema
Attribute|Clinical Attribute|History of Present Illness|2603,2608|true|false|false|C1717255||edema
Event|Event|History of Present Illness|2603,2608|false|false|false|||edema
Finding|Pathologic Function|History of Present Illness|2603,2608|true|false|false|C0013604|Edema|edema
Anatomy|Tissue|History of Present Illness|2610,2617|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|History of Present Illness|2610,2617|false|false|false|C0032226|Pleural Diseases|pleural
Event|Event|History of Present Illness|2619,2628|false|false|false|||effusions
Finding|Pathologic Function|History of Present Illness|2619,2628|false|false|false|C0013687|effusion|effusions
Disorder|Disease or Syndrome|History of Present Illness|2633,2646|false|false|false|C0521530|Lung consolidation|consolidation
Event|Event|History of Present Illness|2633,2646|false|false|false|||consolidation
Event|Event|History of Present Illness|2659,2671|false|false|false|||cardiomegaly
Finding|Finding|History of Present Illness|2659,2671|false|false|false|C0018800|Cardiomegaly|cardiomegaly
Finding|Body Substance|History of Present Illness|2678,2685|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|2678,2685|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|2678,2685|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Organic Chemical|History of Present Illness|2695,2705|false|false|false|C0054836|carvedilol|carvedilol
Drug|Pharmacologic Substance|History of Present Illness|2695,2705|false|false|false|C0054836|carvedilol|carvedilol
Event|Event|History of Present Illness|2695,2705|false|false|false|||carvedilol
Drug|Pharmacologic Substance|History of Present Illness|2707,2717|false|false|false|C2064916|nebulizers (medication)|nebulizers
Event|Event|History of Present Illness|2707,2717|false|false|false|||nebulizers
Drug|Organic Chemical|History of Present Illness|2726,2731|false|false|false|C0699992|Lasix|lasix
Drug|Pharmacologic Substance|History of Present Illness|2726,2731|false|false|false|C0699992|Lasix|lasix
Event|Event|History of Present Illness|2726,2731|false|false|false|||lasix
Finding|Finding|History of Present Illness|2752,2756|false|false|false|C4281574|Much|much
Event|Event|History of Present Illness|2757,2760|false|false|false|||UOP
Finding|Body Substance|History of Present Illness|2765,2772|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|2765,2772|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|2765,2772|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|History of Present Illness|2765,2776|false|false|false|C0332310|Has patient|patient has
Event|Event|History of Present Illness|2791,2801|false|false|false|||documented
Finding|Body Substance|History of Present Illness|2820,2827|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|2820,2827|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|2820,2827|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|2832,2836|false|false|false|||seen
Anatomy|Body System|History of Present Illness|2840,2850|false|false|false|C0007226|Cardiovascular system|cardiology
Event|Event|History of Present Illness|2865,2869|false|false|false|||felt
Event|Event|History of Present Illness|2883,2890|false|false|false|||setting
Finding|Mental Process|History of Present Illness|2883,2890|false|false|false|C0542559|contextual factors|setting
Finding|Organ or Tissue Function|History of Present Illness|2894,2902|false|false|false|C0039155|Systole|systolic
Disorder|Disease or Syndrome|History of Present Illness|2894,2916|false|false|false|C1135191|Heart Failure, Systolic|systolic heart failure
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2903,2908|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|History of Present Illness|2903,2908|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|History of Present Illness|2903,2908|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|History of Present Illness|2903,2916|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Event|Event|History of Present Illness|2909,2916|false|false|false|||failure
Finding|Functional Concept|History of Present Illness|2909,2916|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|History of Present Illness|2909,2916|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|History of Present Illness|2909,2916|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|History of Present Illness|2922,2929|false|false|false|||dyspnea
Finding|Finding|History of Present Illness|2922,2929|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|History of Present Illness|2922,2929|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Finding|History of Present Illness|2934,2940|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|History of Present Illness|2934,2940|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Anatomy|Body Space or Junction|History of Present Illness|2951,2954|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|History of Present Illness|2951,2954|false|false|false|C0018802|Congestive heart failure|CHF
Event|Event|History of Present Illness|2955,2967|false|false|false|||exacerbation
Finding|Finding|History of Present Illness|2955,2967|false|true|false|C4086268|Exacerbation|exacerbation
Event|Event|History of Present Illness|2975,2982|false|false|false|||setting
Finding|Mental Process|History of Present Illness|2975,2982|false|false|false|C0542559|contextual factors|setting
Drug|Food|History of Present Illness|2986,2993|false|false|false|C0012155|Diet|dietary
Event|Event|History of Present Illness|2986,2993|false|false|false|||dietary
Event|Event|History of Present Illness|2995,3007|false|false|false|||indiscretion
Event|Event|History of Present Illness|3009,3017|false|false|false|||Diuresis
Finding|Organ or Tissue Function|History of Present Illness|3009,3017|false|false|false|C0012797|Diuresis|Diuresis
Event|Event|History of Present Illness|3022,3033|false|false|false|||recommended
Finding|Functional Concept|History of Present Illness|3034,3048|false|false|false|C0332287|In addition to|in addition to
Event|Event|History of Present Illness|3037,3045|false|false|false|||addition
Finding|Functional Concept|History of Present Illness|3037,3045|false|false|false|C0332287;C1883712|Add - instruction imperative;In addition to|addition
Event|Event|History of Present Illness|3049,3059|false|false|false|||increasing
Drug|Organic Chemical|History of Present Illness|3061,3071|false|false|false|C0054836|carvedilol|carvedilol
Drug|Pharmacologic Substance|History of Present Illness|3061,3071|false|false|false|C0054836|carvedilol|carvedilol
Event|Event|History of Present Illness|3061,3071|false|false|false|||carvedilol
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|3082,3085|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|3082,3085|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|History of Present Illness|3082,3085|false|false|false|C1530795|BID protein, human|BID
Event|Event|History of Present Illness|3082,3085|false|false|false|||BID
Finding|Gene or Genome|History of Present Illness|3082,3085|false|false|false|C1332410|BID gene|BID
Finding|Finding|History of Present Illness|3090,3094|false|false|false|C5575035|Well (answer to question)|well
Procedure|Diagnostic Procedure|History of Present Illness|3100,3119|false|false|false|C2825165|Nuclear stress test|nuclear stress test
Attribute|Clinical Attribute|History of Present Illness|3108,3114|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|History of Present Illness|3108,3114|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|History of Present Illness|3108,3114|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Finding|Finding|History of Present Illness|3108,3114|false|false|false|C0038435|Stress|stress
Procedure|Diagnostic Procedure|History of Present Illness|3108,3119|false|false|false|C0015260;C3494508|Exercise stress test;Stress Test|stress test
Anatomy|Body Location or Region|History of Present Illness|3115,3119|false|false|false|C4318744|Test - temporal region|test
Finding|Functional Concept|History of Present Illness|3115,3119|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|History of Present Illness|3115,3119|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|History of Present Illness|3115,3119|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|History of Present Illness|3115,3119|false|false|false|C0022885|Laboratory Procedures|test
Anatomy|Anatomical Structure|History of Present Illness|3143,3148|false|false|false|C3714591|Floor (anatomic)|floor
Finding|Body Substance|History of Present Illness|3154,3161|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|3154,3161|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|3154,3161|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|3163,3164|false|false|false|||/
Finding|Finding|History of Present Illness|3174,3182|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Finding|Intellectual Product|History of Present Illness|3174,3182|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Event|Event|History of Present Illness|3183,3190|false|false|false|||dyspnea
Finding|Finding|History of Present Illness|3183,3190|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|History of Present Illness|3183,3190|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Anatomy|Body Location or Region|History of Present Illness|3191,3196|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|3191,3196|false|false|false|C0741025|Chest problem|chest
Event|Event|History of Present Illness|3198,3207|false|false|false|||tightness
Finding|Finding|History of Present Illness|3211,3215|false|false|false|C5575035|Well (answer to question)|well
Event|Event|History of Present Illness|3219,3227|false|false|false|||wheezing
Finding|Sign or Symptom|History of Present Illness|3219,3227|false|false|false|C0043144|Wheezing|wheezing
Disorder|Disease or Syndrome|History of Present Illness|3232,3236|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|History of Present Illness|3232,3236|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|History of Present Illness|3232,3236|false|false|false|||COPD
Finding|Gene or Genome|History of Present Illness|3232,3236|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|History of Present Illness|3237,3243|false|false|false|C0004096|Asthma|asthma
Event|Event|History of Present Illness|3244,3251|false|false|false|||history
Finding|Conceptual Entity|History of Present Illness|3244,3251|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|3244,3251|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|3244,3251|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Event|Event|History of Present Illness|3253,3255|false|false|false|||no
Finding|Idea or Concept|History of Present Illness|3257,3268|false|false|false|C0750502|Significant|significant
Event|Event|History of Present Illness|3269,3276|false|false|false|||smoking
Finding|Individual Behavior|History of Present Illness|3269,3276|false|false|false|C0037369;C0453996;C1548578|Location characteristic ID - Smoking;Smoking;Tobacco smoking behavior|smoking
Finding|Intellectual Product|History of Present Illness|3269,3276|false|false|false|C0037369;C0453996;C1548578|Location characteristic ID - Smoking;Smoking;Tobacco smoking behavior|smoking
Finding|Finding|History of Present Illness|3269,3284|false|false|false|C4721824|Smoking History|smoking history
Event|Event|History of Present Illness|3277,3284|false|false|false|||history
Finding|Conceptual Entity|History of Present Illness|3277,3284|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|3277,3284|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|3277,3284|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Event|Event|History of Present Illness|3308,3313|false|false|false|||acute
Finding|Intellectual Product|History of Present Illness|3308,3313|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|History of Present Illness|3315,3325|false|false|false|||complaints
Finding|Finding|History of Present Illness|3315,3325|false|false|false|C5441521|Complaint (finding)|complaints
Finding|Idea or Concept|History of Present Illness|3337,3346|false|false|false|C0549178|Continuous|continued
Event|Event|History of Present Illness|3347,3350|false|false|false|||SOB
Finding|Sign or Symptom|History of Present Illness|3347,3350|false|false|false|C0013404|Dyspnea|SOB
Event|Event|History of Present Illness|3355,3363|false|false|false|||wheezing
Finding|Sign or Symptom|History of Present Illness|3355,3363|false|false|false|C0043144|Wheezing|wheezing
Event|Event|History of Present Illness|3374,3381|false|false|false|||written
Drug|Pharmacologic Substance|History of Present Illness|3386,3396|false|false|false|C2064916|nebulizers (medication)|nebulizers
Event|Event|History of Present Illness|3386,3396|false|false|false|||nebulizers
Drug|Organic Chemical|History of Present Illness|3401,3409|false|false|false|C0038317|Steroids|steroids
Drug|Pharmacologic Substance|History of Present Illness|3401,3409|false|false|false|C0038317|Steroids|steroids
Event|Event|History of Present Illness|3401,3409|false|false|false|||steroids
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|3414,3422|false|false|false|C4722408|Reactive Therapy|reactive
Disorder|Disease or Syndrome|History of Present Illness|3414,3437|false|false|false|C3714496;C3714497|Chronic obstructive pulmonary disease of horses;Reactive airway disease|reactive airway disease
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|3423,3429|false|false|false|C0458827;C4071894|Airway structure;Chest>Airway|airway
Disorder|Disease or Syndrome|History of Present Illness|3423,3437|false|false|false|C0699949|airway disease|airway disease
Disorder|Disease or Syndrome|History of Present Illness|3430,3437|false|false|false|C0012634|Disease|disease
Event|Event|History of Present Illness|3430,3437|false|false|false|||disease
Event|Event|History of Present Illness|3439,3448|false|false|false|||overnight
Disorder|Disease or Syndrome|Past Medical History|3476,3488|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|Past Medical History|3476,3488|false|false|false|||hypertension
Disorder|Disease or Syndrome|Past Medical History|3493,3501|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|diabetes
Event|Event|Past Medical History|3493,3501|false|false|false|||diabetes
Disorder|Disease or Syndrome|Past Medical History|3509,3512|false|false|false|C0001365;C0038454|Acute ill-defined cerebrovascular disease;Cerebrovascular accident|CVA
Drug|Pharmacologic Substance|Past Medical History|3509,3512|false|false|false|C5779650|Cyclophosphamide/Doxorubicin/Vincristine|CVA
Event|Event|Past Medical History|3509,3512|false|false|false|||CVA
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|3514,3524|false|false|false|C0007765|Cerebellum|cerebellar
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|3525,3534|false|false|false|C0001629;C0025148;C1550278|Adrenal Medulla;Medulla Oblongata;Medullary - body parts|medullary
Disorder|Disease or Syndrome|Past Medical History|3535,3541|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|Past Medical History|3535,3541|false|false|false|||stroke
Finding|Finding|Past Medical History|3535,3541|false|false|false|C5977286|Stroke (heart beat)|stroke
Disorder|Disease or Syndrome|Past Medical History|3553,3556|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Past Medical History|3553,3556|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Past Medical History|3553,3556|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Past Medical History|3553,3556|false|false|false|||CAD
Finding|Gene or Genome|Past Medical History|3553,3556|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Past Medical History|3553,3556|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Past Medical History|3553,3556|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Past Medical History|3553,3556|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|Past Medical History|3574,3577|false|false|false|C0006430|Burning Mouth Syndrome|BMS
Event|Event|Past Medical History|3574,3577|false|false|false|||BMS
Disorder|Disease or Syndrome|Past Medical History|3609,3636|false|false|false|C0085096;C1704436|Peripheral Arterial Diseases;Peripheral Vascular Diseases|peripheral arterial disease
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|3620,3628|false|false|false|C0003842|Arteries|arterial
Disorder|Disease or Syndrome|Past Medical History|3620,3636|false|false|false|C0852949|Arteriopathic disease|arterial disease
Disorder|Disease or Syndrome|Past Medical History|3629,3636|false|false|false|C0012634|Disease|disease
Event|Event|Past Medical History|3629,3636|false|false|false|||disease
Disorder|Disease or Syndrome|Past Medical History|3638,3650|false|true|false|C0021775|Intermittent Claudication|claudication
Event|Event|Past Medical History|3638,3650|false|false|false|||claudication
Finding|Finding|Past Medical History|3638,3650|false|true|false|C0311395;C1456822|Claudication (finding);Lameness|claudication
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|3665,3673|false|false|false|C0005847|Blood Vessel|vascular
Event|Event|Past Medical History|3675,3682|false|false|false|||managed
Attribute|Clinical Attribute|Past Medical History|3700,3705|false|false|false|C1300072|Tumor stage|stage
Finding|Intellectual Product|Past Medical History|3700,3708|false|false|false|C0441772|Stage level 4|stage IV
Disorder|Disease or Syndrome|Past Medical History|3709,3712|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Event|Event|Past Medical History|3709,3712|false|false|false|||CKD
Drug|Biomedical or Dental Material|Past Medical History|3714,3722|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|Past Medical History|3714,3722|false|false|false|||baseline
Finding|Idea or Concept|Past Medical History|3714,3722|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Disorder|Disease or Syndrome|Past Medical History|3736,3740|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|Past Medical History|3736,3740|false|false|false|||GERD
Disorder|Disease or Syndrome|Past Medical History|3741,3751|false|false|false|C0014852|Esophageal Diseases|esophageal
Disorder|Disease or Syndrome|Past Medical History|3741,3757|false|false|false|C0267081|Terminal esophageal web|esophageal rings
Event|Event|Past Medical History|3752,3757|false|false|false|||rings
Event|Activity|Family Medical History|3811,3815|false|false|false|C1947906|Sorting|sort
Event|Event|Family Medical History|3811,3815|false|false|false|||sort
Finding|Cell Function|Family Medical History|3811,3815|false|false|false|C0237886;C0700314|Sorting (Cognition);Sorting - Cell Movement|sort
Finding|Mental Process|Family Medical History|3811,3815|false|false|false|C0237886;C0700314|Sorting (Cognition);Sorting - Cell Movement|sort
Disorder|Neoplastic Process|Family Medical History|3819,3825|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Family Medical History|3819,3825|false|false|false|||cancer
Finding|Conceptual Entity|Family Medical History|3827,3833|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|Family Medical History|3827,3833|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Event|Event|Family Medical History|3834,3838|false|false|false|||died
Anatomy|Body Location or Region|Family Medical History|3858,3862|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3858,3862|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Family Medical History|3858,3862|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Family Medical History|3858,3862|false|false|false|C0740941|Lung Problem|lung
Disorder|Disease or Syndrome|Family Medical History|3858,3870|false|false|false|C0024115|Lung diseases|lung disease
Disorder|Disease or Syndrome|Family Medical History|3863,3870|false|false|false|C0012634|Disease|disease
Event|Event|Family Medical History|3863,3870|false|false|false|||disease
Finding|Idea or Concept|Family Medical History|3873,3879|false|false|false|C1546508|Relationship - Mother|Mother
Event|Event|Family Medical History|3880,3884|false|false|false|||died
Drug|Amino Acid, Peptide, or Protein|Family Medical History|3906,3913|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Immunologic Factor|Family Medical History|3906,3913|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Pharmacologic Substance|Family Medical History|3906,3913|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Event|Event|Family Medical History|3906,3913|false|false|false|||unknown
Finding|Finding|Family Medical History|3906,3913|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Functional Concept|Family Medical History|3906,3913|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Idea or Concept|Family Medical History|3906,3913|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Intellectual Product|Family Medical History|3906,3913|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Event|Event|Family Medical History|3914,3919|false|false|false|||cause
Finding|Conceptual Entity|Family Medical History|3914,3919|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Finding|Functional Concept|Family Medical History|3914,3919|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Disorder|Disease or Syndrome|Family Medical History|3932,3935|true|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Family Medical History|3932,3935|true|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Family Medical History|3932,3935|true|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Family Medical History|3932,3935|false|false|false|||CAD
Finding|Gene or Genome|Family Medical History|3932,3935|true|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Family Medical History|3932,3935|true|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Family Medical History|3932,3935|true|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Family Medical History|3932,3935|true|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Finding|Pathologic Function|Family Medical History|3939,3959|true|false|false|C0085298|Sudden Cardiac Death|sudden cardiac death
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3946,3953|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|Family Medical History|3946,3953|false|false|false|C1314974|Cardiac attachment|cardiac
Finding|Pathologic Function|Family Medical History|3946,3959|true|false|false|C0376297|Cardiac Death|cardiac death
Event|Event|Family Medical History|3954,3959|false|false|false|||death
Finding|Finding|Family Medical History|3954,3959|false|false|false|C0011065;C1306577;C1546949|Cessation of life;Death (finding);Event Consequence - Death|death
Finding|Idea or Concept|Family Medical History|3954,3959|false|false|false|C0011065;C1306577;C1546949|Cessation of life;Death (finding);Event Consequence - Death|death
Finding|Organism Function|Family Medical History|3954,3959|false|false|false|C0011065;C1306577;C1546949|Cessation of life;Death (finding);Event Consequence - Death|death
Event|Event|Family Medical History|3976,3983|false|false|false|||history
Finding|Conceptual Entity|Family Medical History|3976,3983|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|3976,3983|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Family Medical History|3976,3983|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|3976,3986|true|false|false|C0262926|Medical History|history of
Disorder|Neoplastic Process|Family Medical History|3988,3994|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Family Medical History|3988,3994|false|false|false|||cancer
Procedure|Health Care Activity|General Exam|4013,4022|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|General Exam|4023,4031|false|false|false|||PHYSICAL
Finding|Finding|General Exam|4023,4031|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|General Exam|4023,4031|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|General Exam|4023,4031|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|General Exam|4023,4036|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|General Exam|4023,4036|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Event|Event|General Exam|4032,4036|false|false|false|||EXAM
Finding|Functional Concept|General Exam|4032,4036|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|4032,4036|false|false|false|C0582103|Medical Examination|EXAM
Event|Activity|General Exam|4149,4154|false|false|false|C1283174||check
Event|Event|General Exam|4149,4154|false|false|false|||check
Finding|Functional Concept|General Exam|4149,4154|false|false|false|C4321547|Check|check
Drug|Amino Acid, Peptide, or Protein|General Exam|4160,4163|false|false|false|C2744672|SAT1 protein, human|Sat
Drug|Enzyme|General Exam|4160,4163|false|false|false|C2744672|SAT1 protein, human|Sat
Finding|Gene or Genome|General Exam|4160,4163|false|false|false|C0871290;C1705827;C1822614|College Entrance Examination Board Scholastic Aptitude Test;SAT1 gene;SAT1 wt Allele|Sat
Finding|Intellectual Product|General Exam|4160,4163|false|false|false|C0871290;C1705827;C1822614|College Entrance Examination Board Scholastic Aptitude Test;SAT1 gene;SAT1 wt Allele|Sat
Event|Event|General Exam|4184,4191|false|false|false|||General
Finding|Classification|General Exam|4184,4191|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|General Exam|4184,4191|false|false|false|C3812897|General medical service|General
Disorder|Disease or Syndrome|General Exam|4193,4198|false|false|false|C0028754|Obesity|Obese
Event|Event|General Exam|4205,4210|false|false|false|||lying
Disorder|Disease or Syndrome|General Exam|4214,4217|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Event|Event|General Exam|4214,4217|false|false|false|||bed
Finding|Intellectual Product|General Exam|4214,4217|false|false|false|C2346952|Bachelor of Education|bed
Disorder|Disease or Syndrome|General Exam|4221,4224|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|4221,4224|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|4221,4224|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|4221,4224|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|4221,4224|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|General Exam|4221,4224|false|false|false|||NAD
Finding|Finding|General Exam|4221,4224|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Event|Event|General Exam|4234,4242|false|false|false|||wheezing
Finding|Sign or Symptom|General Exam|4234,4242|false|false|false|C0043144|Wheezing|wheezing
Event|Event|General Exam|4254,4263|false|false|false|||tachypnea
Finding|Finding|General Exam|4254,4263|false|false|false|C0231835|Tachypnea|tachypnea
Event|Event|General Exam|4265,4273|false|false|false|||Speaking
Finding|Individual Behavior|General Exam|4265,4273|false|false|false|C0234856|Speaking (function)|Speaking
Finding|Idea or Concept|General Exam|4281,4285|false|false|false|C1705313|Term (lexical)|word
Event|Event|General Exam|4286,4295|false|false|false|||sentences
Finding|Intellectual Product|General Exam|4286,4295|false|false|true|C0876929|Sentence|sentences
Finding|Finding|General Exam|4301,4312|false|false|true|C0278085|Bradylalia|slow speech
Event|Event|General Exam|4306,4312|false|false|false|||speech
Finding|Organism Function|General Exam|4306,4312|false|false|false|C0037817|Speech|speech
Procedure|Diagnostic Procedure|General Exam|4306,4312|false|false|false|C0846595|Speech assessment|speech
Anatomy|Body Location or Region|General Exam|4314,4319|false|false|false|C1512338|HEENT|HEENT
Event|Event|General Exam|4321,4326|false|false|false|||PERRL
Finding|Finding|General Exam|4321,4326|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Event|Event|General Exam|4328,4332|false|false|false|||EOMI
Disorder|Disease or Syndrome|General Exam|4351,4360|false|false|false|C0028738|Nystagmus|nystagmus
Event|Event|General Exam|4351,4360|false|false|false|||nystagmus
Event|Event|General Exam|4374,4378|false|false|false|||gaze
Finding|Finding|General Exam|4374,4378|false|false|false|C0553544|Gaze|gaze
Anatomy|Body Part, Organ, or Organ Component|General Exam|4383,4392|false|false|false|C0229118|Structure of both eyes|both eyes
Anatomy|Body Part, Organ, or Organ Component|General Exam|4388,4392|false|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|General Exam|4388,4392|false|false|false|C5848506||eyes
Disorder|Disease or Syndrome|General Exam|4403,4412|true|false|false|C0028738|Nystagmus|nystagmus
Event|Event|General Exam|4403,4412|false|false|false|||nystagmus
Anatomy|Body Part, Organ, or Organ Component|General Exam|4414,4420|false|false|false|C0036410|Sclera|sclera
Disorder|Disease or Syndrome|General Exam|4414,4420|false|false|false|C0036412|Scleral Diseases|sclera
Event|Event|General Exam|4414,4420|false|false|false|||sclera
Procedure|Health Care Activity|General Exam|4414,4420|false|false|false|C2228481|examination of sclera|sclera
Event|Event|General Exam|4421,4430|false|false|false|||anicteris
Event|Event|General Exam|4432,4436|false|false|false|||some
Event|Event|General Exam|4451,4457|false|false|false|||pallor
Finding|Finding|General Exam|4451,4457|false|false|false|C0241137|Pallor of skin|pallor
Anatomy|Body Part, Organ, or Organ Component|General Exam|4459,4462|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|General Exam|4459,4462|false|false|false|C0026987|Myelofibrosis|MMM
Finding|Idea or Concept|General Exam|4464,4469|false|false|false|C1550016|Remote control command - Clear|clear
Disorder|Disease or Syndrome|General Exam|4470,4479|false|false|false|C0751438|Posterior pituitary disease|posterior
Event|Event|General Exam|4487,4494|false|false|false|||lesions
Finding|Finding|General Exam|4487,4494|true|false|false|C0221198|Lesion|lesions
Finding|Conceptual Entity|General Exam|4497,4506|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|General Exam|4497,4506|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Anatomy|Body Part, Organ, or Organ Component|General Exam|4507,4513|false|false|false|C0700374|Palate|palate
Event|Event|General Exam|4514,4523|false|false|false|||elevation
Procedure|Therapeutic or Preventive Procedure|General Exam|4514,4523|false|false|false|C0439775|Elevation procedure|elevation
Anatomy|Body Part, Organ, or Organ Component|General Exam|4525,4531|false|false|false|C0040408|Tongue|tongue
Disorder|Neoplastic Process|General Exam|4525,4531|false|false|false|C0153933|Benign neoplasm of tongue|tongue
Procedure|Health Care Activity|General Exam|4525,4531|false|false|false|C0872394|Procedure on tongue|tongue
Finding|Finding|General Exam|4525,4539|false|false|false|C3693372|tongue midline|tongue midline
Anatomy|Cell Component|General Exam|4532,4539|false|false|false|C1660780|midline cell component|midline
Anatomy|Body Location or Region|General Exam|4541,4545|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|General Exam|4541,4545|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|General Exam|4541,4545|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Anatomy|Body Location or Region|General Exam|4550,4558|false|false|false|C0027530|Neck|cervical
Anatomy|Body Part, Organ, or Organ Component|General Exam|4575,4578|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|General Exam|4575,4578|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|General Exam|4575,4578|false|false|false|||LAD
Finding|Gene or Genome|General Exam|4575,4578|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Event|General Exam|4591,4594|false|false|false|||JVD
Finding|Finding|General Exam|4591,4594|true|false|false|C0425687|Jugular venous engorgement|JVD
Event|Event|General Exam|4596,4605|false|false|false|||difficult
Finding|Finding|General Exam|4596,4605|false|false|false|C0332218|Difficult (qualifier value)|difficult
Event|Event|General Exam|4610,4616|false|false|false|||assess
Anatomy|Anatomical Structure|General Exam|4621,4625|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Anatomy|Body Part, Organ, or Organ Component|General Exam|4621,4625|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Finding|Intellectual Product|General Exam|4621,4625|false|false|false|C1551342|Document Body|body
Procedure|Diagnostic Procedure|General Exam|4621,4633|false|false|false|C1318474|Assessment of body build|body habitus
Event|Event|General Exam|4626,4633|false|false|false|||habitus
Event|Event|General Exam|4639,4642|false|false|false|||RRR
Disorder|Disease or Syndrome|General Exam|4644,4648|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|General Exam|4667,4674|false|false|false|||murmurs
Finding|Finding|General Exam|4667,4674|true|false|false|C0018808|Heart murmur|murmurs
Event|Event|General Exam|4675,4680|false|false|false|||noted
Anatomy|Body Part, Organ, or Organ Component|General Exam|4682,4687|false|false|false|C0024109|Lung|Lungs
Finding|Organism Function|General Exam|4697,4707|false|false|false|C0231800|Expiration, Respiratory|expiratory
Finding|Finding|General Exam|4697,4715|false|false|false|C2235504|expiratory rhonchi|expiratory rhonchi
Event|Event|General Exam|4708,4715|false|false|false|||rhonchi
Finding|Finding|General Exam|4708,4715|false|false|false|C0035508|Rhonchi|rhonchi
Event|Event|General Exam|4733,4741|false|false|false|||wheezing
Finding|Sign or Symptom|General Exam|4733,4741|true|false|false|C0043144|Wheezing|wheezing
Anatomy|Body Location or Region|General Exam|4746,4750|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|General Exam|4746,4750|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|General Exam|4746,4750|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|General Exam|4746,4750|false|false|false|C0740941|Lung Problem|lung
Procedure|Diagnostic Procedure|General Exam|4746,4755|false|false|false|C2228454|examination of lungs|lung exam
Event|Event|General Exam|4751,4755|false|false|false|||exam
Finding|Functional Concept|General Exam|4751,4755|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|General Exam|4751,4755|false|false|false|C0582103|Medical Examination|exam
Event|Event|General Exam|4762,4770|false|false|false|||crackles
Finding|Finding|General Exam|4762,4770|false|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Drug|Chemical Viewed Functionally|General Exam|4784,4789|false|false|false|C0178499|Base|bases
Event|Event|General Exam|4784,4789|false|false|false|||bases
Finding|Intellectual Product|General Exam|4806,4810|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|Poor
Drug|Inorganic Chemical|General Exam|4812,4815|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|General Exam|4812,4815|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|General Exam|4812,4815|false|false|false|C0001861;C3536832|Air (substance);air|air
Finding|Finding|General Exam|4812,4815|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|General Exam|4812,4815|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|General Exam|4812,4815|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Phenomenon|Natural Phenomenon or Process|General Exam|4812,4824|false|false|false|C0001868|Air Movements|air movement
Event|Event|General Exam|4816,4824|false|false|false|||movement
Finding|Organism Function|General Exam|4816,4824|false|false|false|C0026649|Movement|movement
Finding|Intellectual Product|General Exam|4825,4832|false|false|false|C0282416|Overall Publication Type|overall
Anatomy|Body Location or Region|General Exam|4834,4841|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|General Exam|4834,4841|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Event|Event|General Exam|4834,4841|false|false|false|||Abdomen
Finding|Finding|General Exam|4834,4841|false|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|General Exam|4843,4847|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|General Exam|4843,4847|false|false|false|||soft
Disorder|Disease or Syndrome|General Exam|4849,4854|false|false|false|C0028754|Obesity|obese
Event|Event|General Exam|4849,4854|false|false|false|||obese
Event|Event|General Exam|4856,4865|false|false|false|||nontender
Finding|Finding|General Exam|4886,4892|false|false|false|C1299582|Unable|Unable
Event|Event|General Exam|4908,4914|false|false|false|||assess
Event|Event|General Exam|4915,4927|false|false|false|||organomegaly
Finding|Finding|General Exam|4915,4927|false|false|false|C4054315|Organomegaly|organomegaly
Disorder|Congenital Abnormality|General Exam|4942,4945|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|General Exam|4942,4945|false|false|false|||Ext
Finding|Gene or Genome|General Exam|4942,4945|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Finding|Organ or Tissue Function|General Exam|4955,4972|false|false|false|C0232139|Peripheral pulse|peripheral pulses
Drug|Food|General Exam|4966,4972|false|false|false|C5890763||pulses
Event|Event|General Exam|4966,4972|false|false|false|||pulses
Finding|Physiologic Function|General Exam|4966,4972|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|4966,4972|false|false|false|C0034107|Pulse taking|pulses
Finding|Finding|General Exam|4974,4990|false|false|false|C1720001|3+ pitting edema|3+ pitting edema
Finding|Functional Concept|General Exam|4977,4984|false|false|false|C0205323|Pitting|pitting
Finding|Finding|General Exam|4977,4990|false|false|false|C0333243|Pitting edema|pitting edema
Attribute|Clinical Attribute|General Exam|4985,4990|false|false|false|C1717255||edema
Event|Event|General Exam|4985,4990|false|false|false|||edema
Finding|Pathologic Function|General Exam|4985,4990|false|false|false|C0013604|Edema|edema
Anatomy|Body Location or Region|General Exam|4994,4998|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Part, Organ, or Organ Component|General Exam|4994,4998|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Space or Junction|General Exam|4994,4998|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Procedure|Diagnostic Procedure|General Exam|4994,4998|false|false|false|C0562271|Examination of knee joint|knee
Finding|Finding|General Exam|5006,5022|false|false|false|C1720371|2+ pitting edema|2+ pitting edema
Finding|Functional Concept|General Exam|5009,5016|false|false|false|C0205323|Pitting|pitting
Finding|Finding|General Exam|5009,5022|false|false|false|C0333243|Pitting edema|pitting edema
Attribute|Clinical Attribute|General Exam|5017,5022|false|false|false|C1717255||edema
Event|Event|General Exam|5017,5022|false|false|false|||edema
Finding|Pathologic Function|General Exam|5017,5022|false|false|false|C0013604|Edema|edema
Anatomy|Body Part, Organ, or Organ Component|General Exam|5028,5031|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Gene or Genome|General Exam|5040,5043|false|false|false|C1539110|CNDP2 gene|CN2
Event|Event|General Exam|5047,5054|false|false|false|||notable
Finding|Finding|General Exam|5069,5073|false|false|false|C0553544|Gaze|gaze
Disorder|Disease or Syndrome|General Exam|5074,5083|false|false|false|C0028738|Nystagmus|nystagmus
Event|Event|General Exam|5074,5083|false|false|false|||nystagmus
Event|Event|General Exam|5107,5113|false|false|false|||intact
Finding|Finding|General Exam|5107,5113|false|false|false|C1554187|Gender Status - Intact|intact
Attribute|Clinical Attribute|General Exam|5122,5128|false|false|false|C5890614||person
Event|Event|General Exam|5122,5128|false|false|false|||person
Finding|Intellectual Product|General Exam|5122,5128|false|false|false|C1522390|Person Info|person
Event|Event|General Exam|5130,5138|false|false|false|||hospital
Finding|Idea or Concept|General Exam|5130,5138|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|General Exam|5140,5145|false|false|false|||month
Finding|Idea or Concept|General Exam|5140,5145|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|General Exam|5140,5145|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Idea or Concept|General Exam|5147,5151|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|General Exam|5147,5151|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|General Exam|5153,5157|false|false|false|||date
Event|Event|General Exam|5172,5180|false|false|false|||calendar
Event|Event|General Exam|5192,5196|false|false|false|||know
Finding|Pathologic Function|General Exam|5207,5221|true|false|false|C1504476|Pronator drift|pronator drift
Event|Event|General Exam|5216,5221|false|false|false|||drift
Finding|Finding|General Exam|5229,5239|false|false|false|C0240795|positional|positional
Event|Event|General Exam|5240,5246|false|false|false|||tremor
Finding|Sign or Symptom|General Exam|5240,5246|false|false|false|C0040822|Tremor|tremor
Anatomy|Body Part, Organ, or Organ Component|General Exam|5260,5265|false|false|false|C0018563|Hand|hands
Drug|Organic Chemical|General Exam|5267,5270|false|false|false|C0033228|fenofibrate|FNF
Drug|Pharmacologic Substance|General Exam|5267,5270|false|false|false|C0033228|fenofibrate|FNF
Event|Event|General Exam|5267,5270|false|false|false|||FNF
Event|Event|General Exam|5276,5285|false|false|false|||hesitancy
Finding|Finding|General Exam|5276,5285|false|false|false|C0152032;C5779516|Hesitancy (gait);Urinary hesitation|hesitancy
Finding|Sign or Symptom|General Exam|5276,5285|false|false|false|C0152032;C5779516|Hesitancy (gait);Urinary hesitation|hesitancy
Drug|Amino Acid, Peptide, or Protein|General Exam|5290,5293|false|false|false|C0082420|Endoglin, human|end
Drug|Immunologic Factor|General Exam|5290,5293|false|false|false|C0082420|Endoglin, human|end
Finding|Functional Concept|General Exam|5290,5293|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Finding|Gene or Genome|General Exam|5290,5293|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Event|Activity|General Exam|5294,5300|false|false|false|C3266814|Action|action
Event|Event|General Exam|5294,5300|false|false|false|||action
Finding|Functional Concept|General Exam|5294,5300|false|false|false|C0441472;C1552007|Clinical action|action
Finding|Idea or Concept|General Exam|5294,5300|false|false|false|C0441472;C1552007|Clinical action|action
Event|Event|General Exam|5305,5314|false|false|false|||asterixis
Finding|Sign or Symptom|General Exam|5305,5314|true|false|false|C0232766|Asterixis|asterixis
Event|Event|General Exam|5316,5325|false|false|false|||Sensation
Finding|Finding|General Exam|5316,5325|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Finding|Organ or Tissue Function|General Exam|5316,5325|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Procedure|Health Care Activity|General Exam|5316,5325|false|false|false|C2229507|sensory exam|Sensation
Drug|Amino Acid, Peptide, or Protein|General Exam|5329,5334|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|General Exam|5329,5334|false|false|false|C1570446|TNFSF14 protein, human|light
Finding|Finding|General Exam|5329,5334|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|General Exam|5329,5334|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|General Exam|5329,5334|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|General Exam|5329,5334|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|General Exam|5329,5334|false|false|false|C0031765|Phototherapy|light
Finding|Physiologic Function|General Exam|5329,5340|false|false|false|C0423553|Light touch|light touch
Event|Event|General Exam|5335,5340|false|false|false|||touch
Finding|Mental Process|General Exam|5335,5340|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Finding|Organ or Tissue Function|General Exam|5335,5340|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Procedure|Therapeutic or Preventive Procedure|General Exam|5335,5340|false|false|false|C0152054|Therapeutic Touch|touch
Event|Event|General Exam|5350,5356|false|false|false|||intact
Finding|Finding|General Exam|5350,5356|false|false|false|C1554187|Gender Status - Intact|intact
Anatomy|Body Part, Organ, or Organ Component|General Exam|5360,5375|false|false|false|C0278454|All extremities|all extremities
Anatomy|Body Part, Organ, or Organ Component|General Exam|5364,5375|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Finding|Sign or Symptom|General Exam|5380,5394|true|false|false|C0427190|Ataxia, Truncal|truncal ataxia
Disorder|Disease or Syndrome|General Exam|5388,5394|true|false|false|C0007758|Cerebellar Ataxia|ataxia
Event|Event|General Exam|5388,5394|false|false|false|||ataxia
Finding|Pathologic Function|General Exam|5388,5394|true|false|false|C0004134;C1135207|Ataxia;Ataxia as late effect of cerebrovascular disease|ataxia
Finding|Sign or Symptom|General Exam|5388,5394|true|false|false|C0004134;C1135207|Ataxia;Ataxia as late effect of cerebrovascular disease|ataxia
Event|Event|General Exam|5395,5402|false|false|false|||sitting
Finding|Finding|General Exam|5395,5410|false|false|false|C1280451|Sitting upright|sitting upright
Finding|Intellectual Product|General Exam|5403,5410|false|false|false|C1550127|Special Handling Code - Upright|upright
Phenomenon|Human-caused Phenomenon or Process|General Exam|5403,5410|false|false|false|C1550585|Entity Handling - upright|upright
Disorder|Disease or Syndrome|General Exam|5415,5418|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Event|Event|General Exam|5415,5418|false|false|false|||bed
Finding|Intellectual Product|General Exam|5415,5418|false|false|false|C2346952|Bachelor of Education|bed
Event|Event|General Exam|5426,5430|false|false|false|||exam
Finding|Functional Concept|General Exam|5426,5430|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|General Exam|5426,5430|false|false|false|C0582103|Medical Examination|exam
Finding|Finding|General Exam|5432,5436|false|false|false|C0016928|Gait|Gait
Event|Event|General Exam|5437,5444|false|false|false|||testing
Finding|Functional Concept|General Exam|5437,5444|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|testing
Finding|Intellectual Product|General Exam|5437,5444|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|testing
Event|Event|General Exam|5445,5453|false|false|false|||deferred
Event|Event|General Exam|5455,5460|false|false|false|||Noted
Event|Event|General Exam|5469,5479|false|false|false|||repetitive
Event|Event|General Exam|5481,5490|false|false|false|||movements
Finding|Organism Function|General Exam|5481,5490|false|false|false|C0026649|Movement|movements
Finding|Functional Concept|General Exam|5491,5498|false|false|false|C0443144|At rest (qualifier value)|at rest
Drug|Amino Acid, Peptide, or Protein|General Exam|5494,5498|false|false|false|C1742913|REST protein, human|rest
Drug|Biologically Active Substance|General Exam|5494,5498|false|false|false|C1742913|REST protein, human|rest
Event|Event|General Exam|5494,5498|false|false|false|||rest
Finding|Daily or Recreational Activity|General Exam|5494,5498|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Gene or Genome|General Exam|5494,5498|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Molecular Function|General Exam|5494,5498|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Anatomy|Body Part, Organ, or Organ Component|General Exam|5504,5510|false|false|false|C0230371|Structure of left hand|L hand
Anatomy|Body Part, Organ, or Organ Component|General Exam|5506,5510|false|false|false|C0018563;C4285005|Hand;Upper extremity>Hand|hand
Finding|Finding|General Exam|5506,5510|false|false|false|C0741992|Hand problem|hand
Event|Event|General Exam|5521,5527|false|false|false|||sheets
Event|Event|General Exam|5529,5536|false|false|false|||tapping
Finding|Idea or Concept|General Exam|5538,5541|false|false|false|C1548556|Etc.|etc
Finding|Body Substance|General Exam|5554,5561|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|General Exam|5554,5561|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|General Exam|5554,5561|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|General Exam|5562,5569|false|false|false|||unaware
Procedure|Research Activity|General Exam|5562,5569|false|false|false|C0150114|unaware|unaware
Anatomy|Body System|General Exam|5572,5576|false|false|false|C1123023;C4520765|Skin;Skin, Human|Skin
Disorder|Disease or Syndrome|General Exam|5572,5576|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Disorder|Neoplastic Process|General Exam|5572,5576|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Finding|Body Substance|General Exam|5572,5576|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Finding|Intellectual Product|General Exam|5572,5576|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Event|Event|General Exam|5589,5595|false|false|false|||rashes
Finding|Sign or Symptom|General Exam|5589,5595|false|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Disorder|Injury or Poisoning|General Exam|5596,5608|false|false|false|C0015256|Excoriation|excoriations
Event|Event|General Exam|5596,5608|false|false|false|||excoriations
Anatomy|Body Part, Organ, or Organ Component|General Exam|5612,5623|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Anatomy|Body Location or Region|General Exam|5629,5636|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|General Exam|5629,5636|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Event|Event|General Exam|5629,5636|false|false|false|||abdomen
Finding|Finding|General Exam|5629,5636|false|false|false|C0941288|Abdomen problem|abdomen
Finding|Body Substance|General Exam|5644,5653|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|5644,5653|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|5644,5653|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|5644,5653|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|General Exam|5654,5662|false|false|false|||PHYSICAL
Finding|Finding|General Exam|5654,5662|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|General Exam|5654,5662|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|General Exam|5654,5662|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|General Exam|5654,5667|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|General Exam|5654,5667|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Event|Event|General Exam|5663,5667|false|false|false|||EXAM
Finding|Functional Concept|General Exam|5663,5667|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|5663,5667|false|false|false|C0582103|Medical Examination|EXAM
Attribute|Clinical Attribute|General Exam|5722,5725|false|false|false|C0871470|Systolic Pressure|SBP
Drug|Amino Acid, Peptide, or Protein|General Exam|5722,5725|false|false|false|C0085805|Androgen Binding Protein|SBP
Drug|Biologically Active Substance|General Exam|5722,5725|false|false|false|C0085805|Androgen Binding Protein|SBP
Event|Event|General Exam|5722,5725|false|false|false|||SBP
Finding|Gene or Genome|General Exam|5722,5725|false|false|false|C1705296;C3274833|CCHCR1 wt Allele;SHBG wt Allele|SBP
Procedure|Diagnostic Procedure|General Exam|5722,5725|false|false|false|C1306620|Systolic blood pressure measurement|SBP
Attribute|Clinical Attribute|General Exam|5753,5759|false|false|false|C0944911||Weight
Event|Event|General Exam|5753,5759|false|false|false|||Weight
Finding|Finding|General Exam|5753,5759|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|Weight
Finding|Sign or Symptom|General Exam|5753,5759|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|Weight
Procedure|Health Care Activity|General Exam|5753,5759|false|false|false|C1305866|Weighing patient|Weight
Event|Event|General Exam|5769,5776|false|false|false|||General
Finding|Classification|General Exam|5769,5776|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|General Exam|5769,5776|false|false|false|C3812897|General medical service|General
Disorder|Disease or Syndrome|General Exam|5778,5783|false|false|false|C0028754|Obesity|Obese
Event|Event|General Exam|5778,5783|false|false|false|||Obese
Disorder|Disease or Syndrome|General Exam|5793,5796|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|5793,5796|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|5793,5796|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|5793,5796|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|5793,5796|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|General Exam|5793,5796|false|false|false|||NAD
Finding|Finding|General Exam|5793,5796|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|General Exam|5799,5804|false|false|false|C1512338|HEENT|HEENT
Event|Event|General Exam|5806,5811|false|false|false|||PERRL
Finding|Finding|General Exam|5806,5811|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Event|Event|General Exam|5813,5817|false|false|false|||EOMI
Disorder|Disease or Syndrome|General Exam|5836,5845|false|false|false|C0028738|Nystagmus|nystagmus
Event|Event|General Exam|5836,5845|false|false|false|||nystagmus
Event|Event|General Exam|5859,5863|false|false|false|||gaze
Finding|Finding|General Exam|5859,5863|false|false|false|C0553544|Gaze|gaze
Anatomy|Body Part, Organ, or Organ Component|General Exam|5868,5877|false|false|false|C0229118|Structure of both eyes|both eyes
Anatomy|Body Part, Organ, or Organ Component|General Exam|5873,5877|false|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|General Exam|5873,5877|false|false|false|C5848506||eyes
Disorder|Disease or Syndrome|General Exam|5888,5897|true|false|false|C0028738|Nystagmus|nystagmus
Event|Event|General Exam|5888,5897|false|false|false|||nystagmus
Anatomy|Body Part, Organ, or Organ Component|General Exam|5899,5905|false|false|false|C0036410|Sclera|sclera
Disorder|Disease or Syndrome|General Exam|5899,5905|false|false|false|C0036412|Scleral Diseases|sclera
Event|Event|General Exam|5899,5905|false|false|false|||sclera
Procedure|Health Care Activity|General Exam|5899,5905|false|false|false|C2228481|examination of sclera|sclera
Event|Event|General Exam|5906,5915|false|false|false|||anicteris
Event|Event|General Exam|5917,5921|false|false|false|||some
Event|Event|General Exam|5936,5942|false|false|false|||pallor
Finding|Finding|General Exam|5936,5942|false|false|false|C0241137|Pallor of skin|pallor
Anatomy|Body Part, Organ, or Organ Component|General Exam|5944,5947|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|General Exam|5944,5947|false|false|false|C0026987|Myelofibrosis|MMM
Finding|Idea or Concept|General Exam|5949,5954|false|false|false|C1550016|Remote control command - Clear|clear
Disorder|Disease or Syndrome|General Exam|5955,5964|false|false|false|C0751438|Posterior pituitary disease|posterior
Event|Event|General Exam|5972,5979|false|false|false|||lesions
Finding|Finding|General Exam|5972,5979|true|false|false|C0221198|Lesion|lesions
Finding|Conceptual Entity|General Exam|5982,5991|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|General Exam|5982,5991|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Anatomy|Body Part, Organ, or Organ Component|General Exam|5992,5998|false|false|false|C0700374|Palate|palate
Event|Event|General Exam|5999,6008|false|false|false|||elevation
Procedure|Therapeutic or Preventive Procedure|General Exam|5999,6008|false|false|false|C0439775|Elevation procedure|elevation
Anatomy|Body Part, Organ, or Organ Component|General Exam|6010,6016|false|false|false|C0040408|Tongue|tongue
Disorder|Neoplastic Process|General Exam|6010,6016|false|false|false|C0153933|Benign neoplasm of tongue|tongue
Procedure|Health Care Activity|General Exam|6010,6016|false|false|false|C0872394|Procedure on tongue|tongue
Finding|Finding|General Exam|6010,6024|false|false|false|C3693372|tongue midline|tongue midline
Anatomy|Cell Component|General Exam|6017,6024|false|false|false|C1660780|midline cell component|midline
Anatomy|Body Location or Region|General Exam|6028,6032|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|General Exam|6028,6032|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|General Exam|6028,6032|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|General Exam|6045,6048|false|false|false|||JVD
Finding|Finding|General Exam|6045,6048|true|false|false|C0425687|Jugular venous engorgement|JVD
Event|Event|General Exam|6050,6059|false|false|false|||difficult
Finding|Finding|General Exam|6050,6059|false|false|false|C0332218|Difficult (qualifier value)|difficult
Event|Event|General Exam|6063,6069|false|false|false|||assess
Anatomy|Anatomical Structure|General Exam|6074,6078|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Anatomy|Body Part, Organ, or Organ Component|General Exam|6074,6078|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Finding|Intellectual Product|General Exam|6074,6078|false|false|false|C1551342|Document Body|body
Procedure|Diagnostic Procedure|General Exam|6074,6086|false|false|false|C1318474|Assessment of body build|body habitus
Event|Event|General Exam|6079,6086|false|false|false|||habitus
Event|Event|General Exam|6092,6095|false|false|false|||RRR
Disorder|Disease or Syndrome|General Exam|6097,6101|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|General Exam|6120,6127|false|false|false|||murmurs
Finding|Finding|General Exam|6120,6127|true|false|false|C0018808|Heart murmur|murmurs
Event|Event|General Exam|6128,6133|false|false|false|||noted
Anatomy|Body Part, Organ, or Organ Component|General Exam|6135,6140|false|false|false|C0024109|Lung|Lungs
Drug|Organic Chemical|General Exam|6142,6146|false|false|false|C0951233|cetrimonium bromide|CTAB
Event|Event|General Exam|6142,6146|false|false|false|||CTAB
Anatomy|Body Location or Region|General Exam|6148,6155|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|General Exam|6148,6155|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Event|Event|General Exam|6148,6155|false|false|false|||Abdomen
Finding|Finding|General Exam|6148,6155|false|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|General Exam|6157,6161|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|General Exam|6157,6161|false|false|false|||soft
Disorder|Disease or Syndrome|General Exam|6163,6168|false|false|false|C0028754|Obesity|obese
Event|Event|General Exam|6163,6168|false|false|false|||obese
Event|Event|General Exam|6170,6179|false|false|false|||nontender
Finding|Finding|General Exam|6200,6206|false|false|false|C1299582|Unable|Unable
Event|Event|General Exam|6222,6228|false|false|false|||assess
Event|Event|General Exam|6229,6241|false|false|false|||organomegaly
Finding|Finding|General Exam|6229,6241|false|false|false|C4054315|Organomegaly|organomegaly
Disorder|Congenital Abnormality|General Exam|6243,6246|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|General Exam|6243,6246|false|false|false|||Ext
Finding|Gene or Genome|General Exam|6243,6246|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Finding|Organ or Tissue Function|General Exam|6256,6273|false|false|false|C0232139|Peripheral pulse|peripheral pulses
Drug|Food|General Exam|6267,6273|false|false|false|C5890763||pulses
Event|Event|General Exam|6267,6273|false|false|false|||pulses
Finding|Physiologic Function|General Exam|6267,6273|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|6267,6273|false|false|false|C0034107|Pulse taking|pulses
Finding|Functional Concept|General Exam|6278,6285|true|false|false|C0205323|Pitting|pitting
Finding|Finding|General Exam|6278,6291|true|false|false|C0333243|Pitting edema|pitting edema
Attribute|Clinical Attribute|General Exam|6286,6291|true|false|false|C1717255||edema
Event|Event|General Exam|6286,6291|false|false|false|||edema
Finding|Pathologic Function|General Exam|6286,6291|true|false|false|C0013604|Edema|edema
Procedure|Health Care Activity|General Exam|6318,6327|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|General Exam|6328,6332|false|false|false|||LABS
Lab|Laboratory or Test Result|General Exam|6328,6332|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|General Exam|6350,6355|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|6350,6355|false|false|false|||BLOOD
Finding|Body Substance|General Exam|6350,6355|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|6356,6359|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|6364,6367|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|6364,6367|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|6364,6367|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|6374,6377|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|6374,6377|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|6374,6377|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|6374,6377|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|6383,6386|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|6383,6386|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|6394,6397|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|6394,6397|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|6394,6397|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|6394,6397|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|6394,6397|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|6401,6404|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|6401,6404|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|6401,6404|false|false|false|||MCH
Finding|Gene or Genome|General Exam|6401,6404|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|6401,6404|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|6401,6404|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|6410,6414|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|6410,6414|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|6429,6432|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|6449,6454|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|6449,6454|false|false|false|||BLOOD
Finding|Body Substance|General Exam|6449,6454|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Antibiotic|General Exam|6471,6476|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|General Exam|6471,6476|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|General Exam|6471,6476|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|General Exam|6481,6484|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Event|Event|General Exam|6481,6484|false|false|false|||Eos
Finding|Gene or Genome|General Exam|6481,6484|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|General Exam|6511,6516|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|6511,6516|false|false|false|||BLOOD
Finding|Body Substance|General Exam|6511,6516|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|6521,6524|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|General Exam|6521,6524|false|false|false|||PTT
Procedure|Laboratory Procedure|General Exam|6521,6524|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|General Exam|6547,6552|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|6547,6552|false|false|false|||BLOOD
Finding|Body Substance|General Exam|6547,6552|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|6547,6560|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|6547,6560|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|6547,6560|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|6553,6560|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|6553,6560|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|6553,6560|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|6553,6560|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|6553,6560|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|6553,6560|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|6608,6612|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|6608,6612|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|6608,6612|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|6637,6642|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|6637,6642|false|false|false|||BLOOD
Finding|Body Substance|General Exam|6637,6642|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|6637,6650|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|General Exam|6643,6650|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|6643,6650|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|6643,6650|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|6643,6650|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|6643,6650|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|General Exam|6643,6650|false|false|false|||Calcium
Finding|Physiologic Function|General Exam|6643,6650|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|6643,6650|false|false|false|C0201925|Calcium measurement|Calcium
Finding|Body Substance|General Exam|6686,6691|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|6686,6691|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|6686,6691|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Finding|General Exam|6686,6697|false|false|false|C0278030|Color of urine|URINE Color
Drug|Biomedical or Dental Material|General Exam|6692,6697|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|Color
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|6692,6697|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|Color
Finding|Idea or Concept|General Exam|6712,6717|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Body Substance|General Exam|6737,6742|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|6737,6742|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|6737,6742|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Disorder|Disease or Syndrome|General Exam|6737,6748|false|false|false|C0018965|Hematuria|URINE Blood
Disorder|Disease or Syndrome|General Exam|6743,6748|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Finding|Body Substance|General Exam|6743,6748|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Event|Event|General Exam|6749,6752|false|false|false|||NEG
Finding|Finding|General Exam|6749,6752|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|General Exam|6753,6760|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Drug|Inorganic Chemical|General Exam|6753,6760|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Drug|Pharmacologic Substance|General Exam|6753,6760|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Finding|Finding|General Exam|6761,6764|false|false|false|C5848551|Neg - answer|NEG
Drug|Amino Acid, Peptide, or Protein|General Exam|6765,6772|false|false|false|C0033684|Proteins|Protein
Drug|Biologically Active Substance|General Exam|6765,6772|false|false|false|C0033684|Proteins|Protein
Event|Event|General Exam|6765,6772|false|false|false|||Protein
Finding|Conceptual Entity|General Exam|6765,6772|false|false|false|C1521746|Protein Info|Protein
Procedure|Laboratory Procedure|General Exam|6765,6772|false|false|false|C0202202|Protein measurement|Protein
Drug|Biologically Active Substance|General Exam|6778,6785|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|6778,6785|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|6778,6785|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|6778,6785|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|6778,6785|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|6778,6785|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Organic Chemical|General Exam|6790,6796|false|false|false|C0022634|Ketones|Ketone
Event|Event|General Exam|6797,6800|false|false|false|||NEG
Finding|Finding|General Exam|6797,6800|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|General Exam|6809,6812|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|General Exam|6821,6824|false|false|false|C5848551|Neg - answer|NEG
Finding|Body Substance|General Exam|6854,6859|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|6854,6859|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|6854,6859|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Lab|Laboratory or Test Result|General Exam|6854,6863|false|false|false|C0221752;C2188659|Red blood cells urine positive|URINE RBC
Anatomy|Cell|General Exam|6860,6863|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|6860,6863|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|6860,6863|false|false|false|C0014792|Erythrocytes|RBC
Anatomy|Cell|General Exam|6866,6869|false|false|false|C0023516|Leukocytes|WBC
Drug|Food|General Exam|6884,6889|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Immunologic Factor|General Exam|6884,6889|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|6884,6889|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Pharmacologic Substance|General Exam|6884,6889|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Disorder|Disease or Syndrome|General Exam|6895,6898|false|false|false|C0267963|Exocrine pancreatic insufficiency|Epi
Drug|Amino Acid, Peptide, or Protein|General Exam|6895,6898|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Biologically Active Substance|General Exam|6895,6898|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Hormone|General Exam|6895,6898|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Organic Chemical|General Exam|6895,6898|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Pharmacologic Substance|General Exam|6895,6898|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Event|Event|General Exam|6895,6898|false|false|false|||Epi
Finding|Gene or Genome|General Exam|6895,6898|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|Epi
Finding|Intellectual Product|General Exam|6895,6898|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|Epi
Procedure|Diagnostic Procedure|General Exam|6895,6898|false|false|false|C0162734;C3641909|Echo-Planar Imaging;Electronic Portal Imaging|Epi
Finding|Body Substance|General Exam|6913,6918|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|6913,6918|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|6913,6918|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Disorder|Disease or Syndrome|General Exam|6942,6947|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|6942,6947|false|false|false|||BLOOD
Finding|Body Substance|General Exam|6942,6947|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|6962,6968|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Drug|Hormone|General Exam|6962,6968|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Disorder|Disease or Syndrome|General Exam|6987,6992|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|6987,6992|false|false|false|||BLOOD
Finding|Body Substance|General Exam|6987,6992|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Event|General Exam|7013,7020|false|false|false|||IMAGING
Finding|Finding|General Exam|7013,7020|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|General Exam|7013,7020|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Anatomy|Body Location or Region|General Exam|7031,7036|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|CHEST
Finding|Finding|General Exam|7031,7036|false|false|false|C0741025|Chest problem|CHEST
Drug|Amino Acid, Peptide, or Protein|General Exam|7045,7048|false|false|false|C1366678;C1433371;C4049852|L-Type Amino Acid Transporter;LAT protein, human;ORC3 protein, human|LAT
Drug|Biologically Active Substance|General Exam|7045,7048|false|false|false|C1366678;C1433371;C4049852|L-Type Amino Acid Transporter;LAT protein, human;ORC3 protein, human|LAT
Drug|Immunologic Factor|General Exam|7045,7048|false|false|false|C1366678;C1433371;C4049852|L-Type Amino Acid Transporter;LAT protein, human;ORC3 protein, human|LAT
Event|Event|General Exam|7045,7048|false|false|false|||LAT
Finding|Gene or Genome|General Exam|7045,7048|false|false|false|C1335085;C1425844;C1705279;C2240043|LAT gene;ORC3 gene;ORC3 wt Allele;SPNS1 gene|LAT
Anatomy|Body Part, Organ, or Organ Component|General Exam|7055,7060|false|false|false|C0024109|Lung|lungs
Event|Event|General Exam|7065,7070|false|false|false|||clear
Finding|Idea or Concept|General Exam|7065,7070|false|false|false|C1550016|Remote control command - Clear|clear
Disorder|Disease or Syndrome|General Exam|7074,7087|false|false|false|C0521530|Lung consolidation|consolidation
Event|Event|General Exam|7074,7087|false|false|false|||consolidation
Event|Event|General Exam|7089,7097|false|false|false|||effusion
Finding|Body Substance|General Exam|7089,7097|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|General Exam|7089,7097|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|General Exam|7089,7097|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Attribute|Clinical Attribute|General Exam|7102,7107|false|false|false|C1717255||edema
Event|Event|General Exam|7102,7107|false|false|false|||edema
Finding|Pathologic Function|General Exam|7102,7107|false|false|false|C0013604|Edema|edema
Anatomy|Body Part, Organ, or Organ Component|General Exam|7110,7117|false|false|false|C0018787|Heart|Cardiac
Finding|Intellectual Product|General Exam|7110,7117|false|false|false|C1314974|Cardiac attachment|Cardiac
Anatomy|Body Location or Region|General Exam|7110,7128|false|false|false|C0507134|Cardiac shadow viewed radiologically|Cardiac silhouette
Event|Event|General Exam|7136,7142|false|false|false|||normal
Finding|Functional Concept|General Exam|7144,7154|false|false|false|C1547177|Sequencing - Descending|Descending
Anatomy|Body Part, Organ, or Organ Component|General Exam|7144,7169|false|false|false|C1522460;C3163626|Descending thoracic aorta;Thoracic aorta|Descending thoracic aorta
Anatomy|Body Location or Region|General Exam|7155,7163|false|false|false|C0817096|Chest|thoracic
Disorder|Disease or Syndrome|General Exam|7155,7163|false|false|false|C5779551|Dissecting Thoracic Aortic Aneurysm|thoracic
Anatomy|Body Part, Organ, or Organ Component|General Exam|7155,7169|false|false|false|C1522460;C4037977|Chest>Aorta.thoracic;Thoracic aorta|thoracic aorta
Anatomy|Body Part, Organ, or Organ Component|General Exam|7164,7169|false|false|false|C0003483;C4037978|Aorta;Chest+Abdomen>Aorta|aorta
Procedure|Health Care Activity|General Exam|7164,7169|false|false|false|C0869784|Procedure on aorta|aorta
Event|Event|General Exam|7174,7182|false|false|false|||tortuous
Finding|Finding|General Exam|7174,7182|true|false|false|C4068863|Tortuous|tortuous
Finding|Functional Concept|General Exam|7188,7203|false|false|false|C0333482|atherosclerotic|atherosclerotic
Event|Event|General Exam|7204,7217|false|false|false|||calcification
Finding|Organ or Tissue Function|General Exam|7204,7217|false|false|false|C0006660;C0006663;C1533591|Calcification;Calcinosis;Physiologic calcification|calcification
Finding|Pathologic Function|General Exam|7204,7217|false|false|false|C0006660;C0006663;C1533591|Calcification;Calcinosis;Physiologic calcification|calcification
Event|Event|General Exam|7218,7222|false|false|false|||seen
Anatomy|Body Location or Region|General Exam|7230,7234|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Anatomy|Body Part, Organ, or Organ Component|General Exam|7230,7234|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Anatomy|Body Space or Junction|General Exam|7230,7234|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Finding|Finding|General Exam|7230,7234|false|false|false|C1538146;C4722404|Age-Related Clonal Hematopoiesis;ZBTB8OS gene|arch
Finding|Gene or Genome|General Exam|7230,7234|false|false|false|C1538146;C4722404|Age-Related Clonal Hematopoiesis;ZBTB8OS gene|arch
Finding|Intellectual Product|General Exam|7240,7245|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Part, Organ, or Organ Component|General Exam|7246,7253|false|false|false|C0262950;C4520924|Bone Tissue, Human;Skeletal bone|osseous
Anatomy|Tissue|General Exam|7246,7253|false|false|false|C0262950;C4520924|Bone Tissue, Human;Skeletal bone|osseous
Disorder|Congenital Abnormality|General Exam|7254,7267|false|false|false|C0000768|Congenital Abnormality|abnormalities
Event|Event|General Exam|7254,7267|false|false|false|||abnormalities
Finding|Functional Concept|General Exam|7254,7267|false|false|false|C0000769|teratologic|abnormalities
Event|Event|General Exam|7268,7278|false|false|false|||identified
Finding|Intellectual Product|Impression|7298,7303|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Location or Region|Impression|7304,7319|false|false|false|C0553534|Cardiopulmonary|cardiopulmonary
Disorder|Disease or Syndrome|Impression|7304,7319|false|false|false|C4072686|Cardiovascular disease+Pulmonary disease|cardiopulmonary
Anatomy|Body Part, Organ, or Organ Component|Impression|7320,7327|false|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|Impression|7320,7327|true|false|false|C1951340|Process Pharmacologic Substance|process
Event|Event|Impression|7320,7327|false|false|false|||process
Finding|Functional Concept|Impression|7320,7327|true|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|Impression|7320,7327|true|false|false|C1522240|Process|process
Event|Event|Impression|7336,7340|false|false|false|||MIBI
Procedure|Laboratory Procedure|Impression|7336,7340|false|false|false|C5557372|Multiplexed Ion Beam Imaging|MIBI
Finding|Intellectual Product|Impression|7342,7350|false|false|false|C1315013|Clinical NEC (not elsewhere classified in LNC)|Clinical
Attribute|Clinical Attribute|Impression|7342,7361|false|false|false|C5890495||Clinical Indication
Finding|Functional Concept|Impression|7342,7361|false|false|false|C5670000|Clinical indication|Clinical Indication
Attribute|Clinical Attribute|Impression|7351,7361|false|false|false|C5890010||Indication
Event|Event|Impression|7351,7361|false|false|false|||Indication
Finding|Idea or Concept|Impression|7351,7361|false|false|false|C0392360;C3146298|Indication;Indication of (contextual qualifier)|Indication
Anatomy|Body Location or Region|Impression|7366,7371|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|CHEST
Finding|Finding|Impression|7366,7371|false|false|false|C0741025|Chest problem|CHEST
Finding|Sign or Symptom|Impression|7366,7381|false|false|false|C0232292|Chest tightness|CHEST TIGHTNESS
Event|Event|Impression|7382,7388|false|false|false|||ASSESS
Finding|Idea or Concept|Impression|7393,7401|false|false|false|C3887511|Evidence|EVIDENCE
Finding|Functional Concept|Impression|7393,7404|false|false|false|C0332120|Evidence of (contextual qualifier)|EVIDENCE OF
Event|Event|Impression|7402,7404|false|false|false|||OF
Event|Event|Impression|7406,7414|false|false|false|||ISCHEMIA
Finding|Pathologic Function|Impression|7406,7414|false|false|false|C0022116|Ischemia|ISCHEMIA
Procedure|Therapeutic or Preventive Procedure|Impression|7406,7414|false|false|false|C4321499|Ischemia Procedure|ISCHEMIA
Event|Event|Impression|7417,7424|false|false|false|||HISTORY
Finding|Conceptual Entity|Impression|7417,7424|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|HISTORY
Finding|Finding|Impression|7417,7424|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|HISTORY
Finding|Functional Concept|Impression|7417,7424|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|HISTORY
Event|Event|Impression|7446,7453|false|false|false|||history
Finding|Conceptual Entity|Impression|7446,7453|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Impression|7446,7453|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Impression|7446,7453|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Impression|7446,7456|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|Impression|7457,7460|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Impression|7457,7460|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Impression|7457,7460|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Impression|7457,7460|false|false|false|||CAD
Finding|Gene or Genome|Impression|7457,7460|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Impression|7457,7460|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Impression|7457,7460|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Impression|7457,7460|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Anatomy|Body Space or Junction|Impression|7465,7468|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|Impression|7465,7468|false|false|false|C0018802|Congestive heart failure|CHF
Event|Event|Impression|7465,7468|false|false|false|||CHF
Event|Event|Impression|7469,7477|false|false|false|||referred
Event|Event|Impression|7483,7493|false|false|false|||evaluation
Finding|Idea or Concept|Impression|7483,7493|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|Impression|7483,7493|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Anatomy|Body Location or Region|Impression|7497,7502|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Impression|7497,7502|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Impression|7497,7507|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Impression|7497,7507|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Impression|7503,7507|false|false|false|C2598155||pain
Event|Event|Impression|7503,7507|false|false|false|||pain
Finding|Functional Concept|Impression|7503,7507|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Impression|7503,7507|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Impression|7512,7519|false|false|false|||dyspnea
Finding|Finding|Impression|7512,7519|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|Impression|7512,7519|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Event|Event|Impression|7522,7529|false|false|false|||SUMMARY
Finding|Intellectual Product|Impression|7522,7529|false|false|false|C1552616;C1706244|Summary (document);summary - ActRelationshipSubset|SUMMARY
Event|Event|Impression|7539,7547|false|false|false|||EXERCISE
Finding|Daily or Recreational Activity|Impression|7539,7547|false|false|false|C0015259|Exercise|EXERCISE
Procedure|Therapeutic or Preventive Procedure|Impression|7539,7547|false|false|false|C1522704|Exercise Pain Management|EXERCISE
Event|Event|Impression|7548,7551|false|false|false|||LAB
Finding|Gene or Genome|Impression|7548,7551|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|LAB
Finding|Intellectual Product|Impression|7548,7551|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|LAB
Finding|Functional Concept|Impression|7558,7571|false|false|false|C0205464|pharmacological|pharmacologic
Anatomy|Body Part, Organ, or Organ Component|Impression|7572,7580|false|false|false|C0018787|Heart|coronary
Finding|Organ or Tissue Function|Impression|7581,7595|false|false|false|C0042401;C0595862|Vasodilation;Vasodilation disorder|vasodilatation
Finding|Pathologic Function|Impression|7581,7595|false|false|false|C0042401;C0595862|Vasodilation;Vasodilation disorder|vasodilatation
Drug|Organic Chemical|Impression|7596,7608|false|false|false|C0012582|dipyridamole|dipyridamole
Drug|Pharmacologic Substance|Impression|7596,7608|false|false|false|C0012582|dipyridamole|dipyridamole
Event|Event|Impression|7596,7608|false|false|false|||dipyridamole
Event|Event|Impression|7614,7621|false|false|false|||infused
Event|Event|Impression|7655,7659|false|false|false|||dose
Event|Event|Impression|7670,7679|false|false|false|||milligram
Event|Event|Impression|7713,7721|false|false|false|||symptoms
Finding|Functional Concept|Impression|7713,7721|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Impression|7713,7721|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|Impression|7725,7733|false|false|false|||ischemic
Finding|Functional Concept|Impression|7725,7733|true|false|false|C0475224|Ischemic|ischemic
Drug|Amino Acid, Peptide, or Protein|Impression|7735,7738|false|false|false|C0018064|Equine Gonadotropins|ECG
Drug|Hormone|Impression|7735,7738|false|false|false|C0018064|Equine Gonadotropins|ECG
Drug|Pharmacologic Substance|Impression|7735,7738|false|false|false|C0018064|Equine Gonadotropins|ECG
Event|Event|Impression|7735,7738|false|false|false|||ECG
Finding|Intellectual Product|Impression|7735,7738|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|ECG
Procedure|Diagnostic Procedure|Impression|7735,7738|false|false|false|C1623258|Electrocardiography|ECG
Event|Event|Impression|7739,7746|false|false|false|||changes
Finding|Functional Concept|Impression|7739,7746|false|false|false|C0392747|Changing|changes
Drug|Element, Ion, or Isotope|Technique|7761,7768|false|false|false|C0022262|Isotopes|ISOTOPE
Event|Event|Technique|7769,7773|false|false|false|||DATA
Finding|Idea or Concept|Technique|7769,7773|false|false|false|C1511726|Data|DATA
Disorder|Mental or Behavioral Dysfunction|Technique|7786,7789|false|false|false|C1270972|Mild cognitive disorder|mCi
Event|Event|Technique|7786,7789|false|false|false|||mCi
Finding|Gene or Genome|Technique|7786,7789|false|false|false|C3463911;C5890839|MCIDAS gene;MCIDAS wt Allele|mCi
Drug|Indicator, Reagent, or Diagnostic Aid|Technique|7790,7796|false|false|false|C0303611|technetium 99m|Tc-99m
Drug|Indicator, Reagent, or Diagnostic Aid|Technique|7790,7806|false|false|false|C0162680|technetium Tc 99m sestamibi|Tc-99m Sestamibi
Drug|Organic Chemical|Technique|7790,7806|false|false|false|C0162680|technetium Tc 99m sestamibi|Tc-99m Sestamibi
Event|Event|Technique|7793,7796|false|false|false|||99m
Drug|Organic Chemical|Technique|7797,7806|false|false|false|C1337333|SESTAMIBI|Sestamibi
Drug|Pharmacologic Substance|Technique|7797,7806|false|false|false|C1337333|SESTAMIBI|Sestamibi
Drug|Amino Acid, Peptide, or Protein|Technique|7807,7811|false|false|false|C1742913|REST protein, human|Rest
Drug|Biologically Active Substance|Technique|7807,7811|false|false|false|C1742913|REST protein, human|Rest
Event|Event|Technique|7807,7811|false|false|false|||Rest
Finding|Daily or Recreational Activity|Technique|7807,7811|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|Rest
Finding|Gene or Genome|Technique|7807,7811|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|Rest
Finding|Molecular Function|Technique|7807,7811|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|Rest
Disorder|Mental or Behavioral Dysfunction|Technique|7825,7828|false|false|false|C1270972|Mild cognitive disorder|mCi
Event|Event|Technique|7825,7828|false|false|false|||mCi
Finding|Gene or Genome|Technique|7825,7828|false|false|false|C3463911;C5890839|MCIDAS gene;MCIDAS wt Allele|mCi
Drug|Indicator, Reagent, or Diagnostic Aid|Technique|7829,7835|false|false|false|C0303611|technetium 99m|Tc-99m
Drug|Indicator, Reagent, or Diagnostic Aid|Technique|7829,7845|false|false|false|C0162680|technetium Tc 99m sestamibi|Tc-99m Sestamibi
Drug|Organic Chemical|Technique|7829,7845|false|false|false|C0162680|technetium Tc 99m sestamibi|Tc-99m Sestamibi
Event|Event|Technique|7832,7835|false|false|false|||99m
Drug|Organic Chemical|Technique|7836,7845|false|false|false|C1337333|SESTAMIBI|Sestamibi
Drug|Pharmacologic Substance|Technique|7836,7845|false|false|false|C1337333|SESTAMIBI|Sestamibi
Attribute|Clinical Attribute|Technique|7846,7852|false|false|false|C1718621|W stress|Stress
Drug|Organic Chemical|Technique|7846,7852|false|false|false|C0723460|Stress bismuth subsalicylate|Stress
Drug|Pharmacologic Substance|Technique|7846,7852|false|false|false|C0723460|Stress bismuth subsalicylate|Stress
Event|Event|Technique|7846,7852|false|false|false|||Stress
Finding|Finding|Technique|7846,7852|false|false|false|C0038435|Stress|Stress
Drug|Pharmacologic Substance|Technique|7854,7858|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|DRUG
Event|Event|Technique|7854,7858|false|false|false|||DRUG
Finding|Finding|Technique|7854,7858|false|false|false|C0740721|Drug problem|DRUG
Event|Event|Technique|7859,7863|false|false|false|||DATA
Finding|Idea or Concept|Technique|7859,7863|false|false|false|C1511726|Data|DATA
Event|Event|Technique|7874,7879|false|false|false|||admin
Event|Occupational Activity|Technique|7874,7879|false|false|false|C0001554|Administration occupational activities|admin
Finding|Intellectual Product|Technique|7874,7879|false|false|false|C4084955|Administrative - Clinical Class|admin
Drug|Organic Chemical|Technique|7881,7893|false|false|false|C0012582|dipyridamole|Dipyridamole
Drug|Pharmacologic Substance|Technique|7881,7893|false|false|false|C0012582|dipyridamole|Dipyridamole
Event|Event|Technique|7881,7893|false|false|false|||Dipyridamole
Event|Event|Technique|7896,7903|false|false|false|||IMAGING
Finding|Finding|Technique|7896,7903|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|Technique|7896,7903|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Finding|Functional Concept|Technique|7896,7910|false|false|false|C1275506|Imaging modality|IMAGING METHOD
Finding|Functional Concept|Technique|7904,7910|false|false|false|C0025663;C0449851;C2828387|Method, LOINC Axis 6;Methods;Techniques|METHOD
Finding|Intellectual Product|Technique|7904,7910|false|false|false|C0025663;C0449851;C2828387|Method, LOINC Axis 6;Methods;Techniques|METHOD
Finding|Daily or Recreational Activity|Technique|7912,7919|false|false|false|C0035253|Rest|Resting
Event|Event|Technique|7920,7929|false|false|false|||perfusion
Finding|Functional Concept|Technique|7920,7929|false|false|false|C4281794;C4723760|Perfusion (biological);Perfusion route|perfusion
Finding|Organism Function|Technique|7920,7929|false|false|false|C4281794;C4723760|Perfusion (biological);Perfusion route|perfusion
Procedure|Therapeutic or Preventive Procedure|Technique|7920,7929|false|false|false|C0031001;C4721534|Chemotherapeutic Perfusion;Perfusion (procedure)|perfusion
Event|Event|Technique|7930,7936|false|false|false|||images
Event|Event|Technique|7942,7950|false|false|false|||obtained
Drug|Indicator, Reagent, or Diagnostic Aid|Technique|7956,7962|false|false|false|C0303611|technetium 99m|Tc-99m
Drug|Indicator, Reagent, or Diagnostic Aid|Technique|7956,7972|false|false|false|C0162680|technetium Tc 99m sestamibi|Tc-99m sestamibi
Drug|Organic Chemical|Technique|7956,7972|false|false|false|C0162680|technetium Tc 99m sestamibi|Tc-99m sestamibi
Drug|Organic Chemical|Technique|7963,7972|false|false|false|C1337333|SESTAMIBI|sestamibi
Drug|Pharmacologic Substance|Technique|7963,7972|false|false|false|C1337333|SESTAMIBI|sestamibi
Event|Event|Technique|7963,7972|false|false|false|||sestamibi
Drug|Indicator, Reagent, or Diagnostic Aid|Technique|7975,7981|false|false|false|C1522485|Tracer|Tracer
Event|Event|Technique|7975,7981|false|false|false|||Tracer
Event|Event|Technique|7986,7994|false|false|false|||injected
Event|Event|Technique|8029,8038|false|false|false|||obtaining
Finding|Daily or Recreational Activity|Technique|8044,8051|false|false|false|C0035253|Rest|resting
Event|Event|Technique|8052,8058|false|false|false|||images
Event|Event|Technique|8079,8085|false|false|false|||images
Finding|Functional Concept|Technique|8100,8111|false|false|false|C1522726|Intravenous Route of Administration|intravenous
Drug|Biomedical or Dental Material|Technique|8100,8120|false|false|false|C1272892|Intravenous infusion (product)|intravenous infusion
Finding|Functional Concept|Technique|8100,8120|false|false|false|C1621368|Intravenous Drip Route of Administration|intravenous infusion
Procedure|Therapeutic or Preventive Procedure|Technique|8100,8120|false|false|false|C0021440|Intravenous infusion procedures|intravenous infusion
Event|Event|Technique|8112,8120|false|false|false|||infusion
Finding|Functional Concept|Technique|8112,8120|false|false|false|C1827465|Infusion route|infusion
Procedure|Therapeutic or Preventive Procedure|Technique|8112,8120|false|false|false|C0574032|Infusion procedures|infusion
Disorder|Disease or Syndrome|Technique|8143,8148|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Daily or Recreational Activity|Technique|8153,8160|false|false|false|C0035253|Rest|resting
Event|Event|Technique|8161,8165|false|false|false|||dose
Drug|Indicator, Reagent, or Diagnostic Aid|Technique|8169,8175|false|false|false|C0303611|technetium 99m|Tc-99m
Drug|Indicator, Reagent, or Diagnostic Aid|Technique|8169,8185|false|false|false|C0162680|technetium Tc 99m sestamibi|Tc-99m sestamibi
Drug|Organic Chemical|Technique|8169,8185|false|false|false|C0162680|technetium Tc 99m sestamibi|Tc-99m sestamibi
Drug|Organic Chemical|Technique|8176,8185|false|false|false|C1337333|SESTAMIBI|sestamibi
Drug|Pharmacologic Substance|Technique|8176,8185|false|false|false|C1337333|SESTAMIBI|sestamibi
Event|Event|Technique|8176,8185|false|false|false|||sestamibi
Event|Event|Technique|8191,8203|false|false|false|||administered
Procedure|Therapeutic or Preventive Procedure|Technique|8191,8217|false|false|false|C1737200|Administered intravenously|administered intravenously
Attribute|Clinical Attribute|Technique|8219,8225|false|false|false|C1718621|W stress|Stress
Drug|Organic Chemical|Technique|8219,8225|false|false|false|C0723460|Stress bismuth subsalicylate|Stress
Drug|Pharmacologic Substance|Technique|8219,8225|false|false|false|C0723460|Stress bismuth subsalicylate|Stress
Finding|Finding|Technique|8219,8225|false|false|false|C0038435|Stress|Stress
Event|Event|Technique|8226,8232|false|false|false|||images
Event|Event|Technique|8238,8246|false|false|false|||obtained
Drug|Indicator, Reagent, or Diagnostic Aid|Technique|8283,8289|false|false|false|C1522485|Tracer|tracer
Drug|Biomedical or Dental Material|Technique|8290,8299|false|false|false|C1272883|Injection|injection
Event|Event|Technique|8290,8299|false|false|false|||injection
Finding|Functional Concept|Technique|8290,8299|false|false|false|C1828121|Injection Route of Administration|injection
Procedure|Therapeutic or Preventive Procedure|Technique|8290,8299|false|false|false|C0021485;C1533685|Injection of therapeutic agent;Injection procedure|injection
Event|Event|Technique|8302,8309|false|false|false|||Imaging
Finding|Finding|Technique|8302,8309|false|false|false|C0740845|Imaging problem|Imaging
Procedure|Diagnostic Procedure|Technique|8302,8309|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|Imaging
Event|Event|Technique|8310,8318|false|false|false|||protocol
Finding|Finding|Technique|8310,8318|false|false|false|C0442711;C1507394;C1522729;C2348563;C3715209|Clinical trial protocol document;Library Protocol;Protocol - answer to question;Protocols documentation;Study Protocol|protocol
Finding|Intellectual Product|Technique|8310,8318|false|false|false|C0442711;C1507394;C1522729;C2348563;C3715209|Clinical trial protocol document;Library Protocol;Protocol - answer to question;Protocols documentation;Study Protocol|protocol
Finding|Finding|Technique|8320,8325|false|false|false|C4266464|Gated|Gated
Event|Event|Technique|8326,8331|false|false|false|||SPECT
Procedure|Diagnostic Procedure|Technique|8326,8331|false|false|false|C0040399|Tomography, Emission-Computed, Single-Photon|SPECT
Event|Event|Technique|8339,8344|false|false|false|||study
Finding|Intellectual Product|Technique|8339,8344|false|false|false|C1705923|Study Object|study
Procedure|Research Activity|Technique|8339,8344|false|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|study
Event|Event|Technique|8349,8360|false|false|false|||interpreted
Event|Event|Technique|8361,8366|false|false|false|||using
Anatomy|Tissue|Technique|8382,8392|false|false|false|C0027061|Myocardium|myocardial
Event|Event|Technique|8394,8403|false|false|false|||perfusion
Finding|Functional Concept|Technique|8394,8403|false|false|false|C4281794;C4723760|Perfusion (biological);Perfusion route|perfusion
Finding|Organism Function|Technique|8394,8403|false|false|false|C4281794;C4723760|Perfusion (biological);Perfusion route|perfusion
Procedure|Therapeutic or Preventive Procedure|Technique|8394,8403|false|false|false|C0031001;C4721534|Chemotherapeutic Perfusion;Perfusion (procedure)|perfusion
Event|Event|Technique|8404,8409|false|false|false|||model
Finding|Conceptual Entity|Technique|8404,8409|false|false|false|C3161035;C3714583;C3853906|Digital Model Attachment;Model;Model - style/design|model
Finding|Intellectual Product|Technique|8404,8409|false|false|false|C3161035;C3714583;C3853906|Digital Model Attachment;Model;Model - style/design|model
Disorder|Disease or Syndrome|Findings|8428,8433|false|false|false|C1846009|Intrauterine growth restriction, metaphyseal dysplasia, adrenal hypoplasia congenita, and genital anomaly syndrome|image
Event|Event|Findings|8428,8433|false|false|false|||image
Finding|Intellectual Product|Findings|8428,8433|false|false|false|C1696103;C1704254;C1704922;C3542466|Image;Image (foundation metadata concept);Medical Image;image - dosage form|image
Event|Event|Findings|8445,8453|false|false|false|||adequate
Event|Event|Findings|8458,8465|false|false|false|||limited
Finding|Functional Concept|Findings|8458,8465|false|false|false|C0439801;C3542948|Limited (extensiveness);Limited component (foundation metadata concept)|limited
Finding|Intellectual Product|Findings|8458,8465|false|false|false|C0439801;C3542948|Limited (extensiveness);Limited component (foundation metadata concept)|limited
Disorder|Disease or Syndrome|Findings|8473,8477|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Anatomy|Body Location or Region|Findings|8473,8484|false|false|false|C0225317;C4532079|Neck+Chest>Soft tissue;soft tissue|soft tissue
Anatomy|Tissue|Findings|8473,8484|false|false|false|C0225317;C4532079|Neck+Chest>Soft tissue;soft tissue|soft tissue
Anatomy|Tissue|Findings|8478,8484|false|false|false|C0040300|Body tissue|tissue
Finding|Intellectual Product|Findings|8478,8484|false|false|false|C1547928|Tissue Specimen Code|tissue
Anatomy|Body Part, Organ, or Organ Component|Findings|8490,8496|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|Findings|8490,8496|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Event|Event|Findings|8490,8496|false|false|false|||breast
Finding|Finding|Findings|8490,8496|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|Findings|8490,8496|false|false|false|C0191838|Procedures on breast|breast
Event|Activity|Findings|8497,8508|false|false|false|C0599946|Attenuation|attenuation
Event|Event|Findings|8497,8508|false|false|false|||attenuation
Finding|Functional Concept|Findings|8510,8514|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Space or Junction|Findings|8510,8533|false|false|false|C0503990|Cavity of left ventricle|Left ventricular cavity
Attribute|Clinical Attribute|Findings|8510,8538|false|false|false|C0455830|Left ventricular cavity size|Left ventricular cavity size
Anatomy|Body Part, Organ, or Organ Component|Findings|8515,8526|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Space or Junction|Findings|8515,8533|false|false|false|C0507083|Cavity of ventricle|ventricular cavity
Anatomy|Body Space or Junction|Findings|8527,8533|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|Findings|8527,8533|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|Findings|8527,8533|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Event|Event|Findings|8542,8551|false|false|false|||increased
Drug|Amino Acid, Peptide, or Protein|Findings|8553,8557|false|false|false|C1742913|REST protein, human|Rest
Drug|Biologically Active Substance|Findings|8553,8557|false|false|false|C1742913|REST protein, human|Rest
Event|Event|Findings|8553,8557|false|false|false|||Rest
Finding|Daily or Recreational Activity|Findings|8553,8557|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|Rest
Finding|Gene or Genome|Findings|8553,8557|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|Rest
Finding|Molecular Function|Findings|8553,8557|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|Rest
Attribute|Clinical Attribute|Findings|8562,8568|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|Findings|8562,8568|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|Findings|8562,8568|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Event|Event|Findings|8562,8568|false|false|false|||stress
Finding|Finding|Findings|8562,8568|false|false|false|C0038435|Stress|stress
Finding|Functional Concept|Findings|8569,8578|false|false|false|C4281794;C4723760|Perfusion (biological);Perfusion route|perfusion
Finding|Organism Function|Findings|8569,8578|false|false|false|C4281794;C4723760|Perfusion (biological);Perfusion route|perfusion
Procedure|Therapeutic or Preventive Procedure|Findings|8569,8578|false|false|false|C0031001;C4721534|Chemotherapeutic Perfusion;Perfusion (procedure)|perfusion
Event|Event|Findings|8579,8585|false|false|false|||images
Drug|Indicator, Reagent, or Diagnostic Aid|Findings|8601,8607|false|false|false|C1522485|Tracer|tracer
Event|Event|Findings|8608,8614|false|false|false|||uptake
Finding|Cell Function|Findings|8608,8614|false|false|false|C0243144;C3888108;C3893696|Import into cell;Uptake;import across plasma membrane|uptake
Finding|Physiologic Function|Findings|8608,8614|false|false|false|C0243144;C3888108;C3893696|Import into cell;Uptake;import across plasma membrane|uptake
Finding|Functional Concept|Findings|8631,8635|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Findings|8631,8658|false|false|false|C0225899|Myocardium of left ventricle|left ventricular myocardium
Anatomy|Body Part, Organ, or Organ Component|Findings|8636,8647|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Part, Organ, or Organ Component|Findings|8636,8658|false|false|false|C0225880|Structure of myocardium of ventricle|ventricular myocardium
Anatomy|Tissue|Findings|8648,8658|false|false|false|C0027061|Myocardium|myocardium
Finding|Finding|Findings|8661,8666|false|false|false|C4266464|Gated|Gated
Event|Event|Findings|8667,8673|false|false|false|||images
Attribute|Clinical Attribute|Findings|8688,8699|false|false|false|C1980023|Wall motion|wall motion
Event|Event|Findings|8693,8699|false|false|false|||motion
Phenomenon|Natural Phenomenon or Process|Findings|8693,8699|false|false|false|C0026597|Motion|motion
Procedure|Diagnostic Procedure|Findings|8706,8751|false|false|false|C4525750|Calculated Left Ventricular Ejection Fraction|calculated left ventricular ejection fraction
Finding|Functional Concept|Findings|8717,8721|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Physiologic Function|Findings|8717,8742|false|false|false|C2733342|Left ventricular ejection|left ventricular ejection
Attribute|Clinical Attribute|Findings|8717,8751|false|false|false|C0428772;C0488728|Left ventricular ejection fraction|left ventricular ejection fraction
Anatomy|Body Part, Organ, or Organ Component|Findings|8722,8733|false|false|false|C0018827|Heart Ventricle|ventricular
Finding|Physiologic Function|Findings|8722,8742|false|false|false|C2733340|Ventricular ejection|ventricular ejection
Lab|Laboratory or Test Result|Findings|8722,8751|false|false|false|C0042508|Ventricular Ejection Fraction|ventricular ejection fraction
Attribute|Clinical Attribute|Findings|8734,8742|false|false|false|C0812388|Ejection time|ejection
Finding|Daily or Recreational Activity|Findings|8734,8742|false|false|false|C0336969|Ejection as a Sports activity|ejection
Phenomenon|Phenomenon or Process|Findings|8734,8742|false|false|false|C0302131|Ejection as a Circumstance of Injury|ejection
Finding|Finding|Findings|8734,8751|false|false|false|C2020641;C2700378|Ejection fraction;stress echo measurements ejection fraction|ejection fraction
Procedure|Diagnostic Procedure|Findings|8734,8751|false|false|false|C0489482|Ejection fraction (procedure)|ejection fraction
Event|Event|Findings|8743,8751|false|false|false|||fraction
Finding|Intellectual Product|Findings|8743,8751|false|false|false|C1554103|MDFAttributeType - Fraction|fraction
Event|Event|Findings|8768,8771|false|false|false|||EDV
Procedure|Diagnostic Procedure|Findings|8768,8771|false|false|false|C2986747|End Diastolic Volume Imaging|EDV
Anatomy|Tissue|Impression|8806,8816|false|false|false|C0027061|Myocardium|myocardial
Event|Event|Impression|8817,8826|false|false|false|||perfusion
Finding|Functional Concept|Impression|8817,8826|false|false|false|C4281794;C4723760|Perfusion (biological);Perfusion route|perfusion
Finding|Organism Function|Impression|8817,8826|false|false|false|C4281794;C4723760|Perfusion (biological);Perfusion route|perfusion
Procedure|Therapeutic or Preventive Procedure|Impression|8817,8826|false|false|false|C0031001;C4721534|Chemotherapeutic Perfusion;Perfusion (procedure)|perfusion
Event|Event|Impression|8832,8841|false|false|false|||Increased
Finding|Functional Concept|Impression|8842,8846|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Space or Junction|Impression|8842,8865|false|false|false|C0503990|Cavity of left ventricle|left ventricular cavity
Attribute|Clinical Attribute|Impression|8842,8870|false|false|false|C0455830|Left ventricular cavity size|left ventricular cavity size
Anatomy|Body Part, Organ, or Organ Component|Impression|8847,8858|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Space or Junction|Impression|8847,8865|false|false|false|C0507083|Cavity of ventricle|ventricular cavity
Anatomy|Body Space or Junction|Impression|8859,8865|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|Impression|8859,8865|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|Impression|8859,8865|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Event|Event|Impression|8866,8870|false|false|false|||size
Event|Event|Impression|8883,8891|false|false|false|||systolic
Finding|Organ or Tissue Function|Impression|8883,8891|false|false|false|C0039155|Systole|systolic
Event|Event|Impression|8893,8901|false|false|false|||function
Finding|Finding|Impression|8893,8901|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|Impression|8893,8901|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|Impression|8893,8901|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|Impression|8893,8901|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Event|Event|Impression|8903,8911|false|false|false|||Compared
Event|Event|Impression|8923,8928|false|false|false|||study
Finding|Intellectual Product|Impression|8923,8928|false|false|false|C1705923|Study Object|study
Procedure|Research Activity|Impression|8923,8928|false|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|study
Anatomy|Body Space or Junction|Impression|8941,8947|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|Impression|8941,8947|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|Impression|8941,8947|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Finding|Idea or Concept|Hospital Course|8996,9000|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|Hospital Course|8996,9000|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|Hospital Course|9001,9004|false|false|false|||old
Event|Event|Hospital Course|9017,9024|false|false|false|||history
Finding|Conceptual Entity|Hospital Course|9017,9024|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|9017,9024|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|9017,9024|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|9017,9027|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|Hospital Course|9028,9031|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|Hospital Course|9028,9031|false|false|false|||HTN
Disorder|Disease or Syndrome|Hospital Course|9033,9036|false|false|false|C0001365;C0038454|Acute ill-defined cerebrovascular disease;Cerebrovascular accident|CVA
Drug|Pharmacologic Substance|Hospital Course|9033,9036|false|false|false|C5779650|Cyclophosphamide/Doxorubicin/Vincristine|CVA
Event|Event|Hospital Course|9033,9036|false|false|false|||CVA
Disorder|Disease or Syndrome|Hospital Course|9038,9041|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9038,9041|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|9038,9041|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Hospital Course|9038,9041|false|false|false|||CAD
Finding|Gene or Genome|Hospital Course|9038,9041|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|9038,9041|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|9038,9041|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9038,9041|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|Hospital Course|9047,9050|false|false|false|C0006430|Burning Mouth Syndrome|BMS
Event|Event|Hospital Course|9047,9050|false|false|false|||BMS
Event|Event|Hospital Course|9055,9065|false|false|false|||circumflex
Anatomy|Body Space or Junction|Hospital Course|9074,9077|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|Hospital Course|9074,9077|false|false|false|C0018802|Congestive heart failure|CHF
Event|Event|Hospital Course|9097,9106|false|false|false|||presented
Finding|Intellectual Product|Hospital Course|9113,9118|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Intellectual Product|Hospital Course|9113,9124|false|false|false|C1272517|Sudden onset (contextual qualifier) (qualifier value)|acute onset
Event|Event|Hospital Course|9125,9134|false|false|false|||shortness
Attribute|Clinical Attribute|Hospital Course|9125,9144|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|Hospital Course|9125,9144|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|Hospital Course|9138,9144|false|false|false|C0225386|Breath|breath
Anatomy|Body Location or Region|Hospital Course|9160,9165|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|9160,9165|false|false|false|C0741025|Chest problem|chest
Event|Event|Hospital Course|9167,9176|false|false|false|||tightness
Attribute|Clinical Attribute|Hospital Course|9181,9200|false|false|false|C2707305||Shortness of breath
Finding|Sign or Symptom|Hospital Course|9181,9200|false|false|false|C0013404|Dyspnea|Shortness of breath
Finding|Body Substance|Hospital Course|9194,9200|false|false|false|C0225386|Breath|breath
Finding|Body Substance|Hospital Course|9202,9209|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|9202,9209|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|9202,9209|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|9215,9220|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Intellectual Product|Hospital Course|9215,9226|false|false|false|C1272517|Sudden onset (contextual qualifier) (qualifier value)|acute onset
Event|Event|Hospital Course|9227,9230|false|false|false|||SOB
Finding|Sign or Symptom|Hospital Course|9227,9230|false|false|false|C0013404|Dyspnea|SOB
Drug|Food|Hospital Course|9241,9248|false|false|false|C0206208|Seafood|seafood
Event|Event|Hospital Course|9249,9253|false|false|false|||meal
Finding|Daily or Recreational Activity|Hospital Course|9249,9253|false|false|false|C1998602|Meal (occasion for eating)|meal
Anatomy|Body Location or Region|Hospital Course|9271,9276|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|9271,9276|false|false|false|C0741025|Chest problem|chest
Finding|Sign or Symptom|Hospital Course|9271,9286|false|false|false|C0232292|Chest tightness|chest tightness
Event|Event|Hospital Course|9277,9286|false|false|false|||tightness
Event|Event|Hospital Course|9288,9291|false|false|false|||see
Finding|Body Substance|Hospital Course|9300,9307|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|9300,9307|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|9300,9307|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|9313,9321|false|false|false|||crackles
Finding|Finding|Hospital Course|9313,9321|false|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Finding|Organism Function|Hospital Course|9327,9337|false|false|false|C0231800|Expiration, Respiratory|expiratory
Finding|Finding|Hospital Course|9327,9345|false|false|false|C2235504|expiratory rhonchi|expiratory rhonchi
Event|Event|Hospital Course|9338,9345|false|false|false|||rhonchi
Finding|Finding|Hospital Course|9338,9345|false|false|false|C0035508|Rhonchi|rhonchi
Anatomy|Body Location or Region|Hospital Course|9349,9353|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9349,9353|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Hospital Course|9349,9353|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Hospital Course|9349,9353|false|false|false|C0740941|Lung Problem|lung
Procedure|Diagnostic Procedure|Hospital Course|9349,9358|false|false|false|C2228454|examination of lungs|lung exam
Event|Event|Hospital Course|9354,9358|false|false|false|||exam
Finding|Functional Concept|Hospital Course|9354,9358|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|Hospital Course|9354,9358|false|false|false|C0582103|Medical Examination|exam
Event|Event|Hospital Course|9360,9363|false|false|false|||CXR
Procedure|Diagnostic Procedure|Hospital Course|9360,9363|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|Hospital Course|9372,9376|false|false|false|||show
Finding|Idea or Concept|Hospital Course|9378,9389|false|false|false|C0750502|Significant|significant
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9390,9399|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Hospital Course|9390,9399|false|false|false|C2707265||pulmonary
Finding|Finding|Hospital Course|9390,9399|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|Hospital Course|9390,9405|false|false|false|C0034063|Pulmonary Edema|pulmonary edema
Attribute|Clinical Attribute|Hospital Course|9400,9405|false|false|false|C1717255||edema
Event|Event|Hospital Course|9400,9405|false|false|false|||edema
Finding|Pathologic Function|Hospital Course|9400,9405|false|false|false|C0013604|Edema|edema
Anatomy|Tissue|Hospital Course|9407,9414|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|Hospital Course|9407,9414|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Pathologic Function|Hospital Course|9407,9424|false|false|false|C0032227|Pleural effusion (disorder)|pleural effusions
Event|Event|Hospital Course|9415,9424|false|false|false|||effusions
Finding|Pathologic Function|Hospital Course|9415,9424|false|false|false|C0013687|effusion|effusions
Disorder|Disease or Syndrome|Hospital Course|9429,9442|false|false|false|C0521530|Lung consolidation|consolidation
Event|Event|Hospital Course|9429,9442|false|false|false|||consolidation
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9457,9460|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Hormone|Hospital Course|9457,9460|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Pharmacologic Substance|Hospital Course|9457,9460|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Event|Event|Hospital Course|9457,9460|false|false|false|||BNP
Finding|Gene or Genome|Hospital Course|9457,9460|false|false|false|C1417808;C2982014|NPPB gene;NPPB wt Allele|BNP
Procedure|Laboratory Procedure|Hospital Course|9457,9460|false|false|false|C1095989|Brain natriuretic peptide measurement|BNP
Event|Event|Hospital Course|9465,9473|false|false|false|||elevated
Event|Event|Hospital Course|9479,9487|false|false|false|||pharmacy
Finding|Intellectual Product|Hospital Course|9479,9487|false|false|false|C1547997;C3244303|Diagnostic Service Section ID - Pharmacy;Pharmacy domain|pharmacy
Procedure|Health Care Activity|Hospital Course|9479,9487|false|false|false|C0031321|Pharmaceutical Services|pharmacy
Finding|Intellectual Product|Hospital Course|9479,9495|false|false|false|C2600053|Pharmacy records|pharmacy records
Event|Event|Hospital Course|9488,9495|false|false|false|||records
Finding|Idea or Concept|Hospital Course|9488,9495|false|false|false|C0034869;C1548330|Quantity limited request - Records;Records|records
Finding|Intellectual Product|Hospital Course|9488,9495|false|false|false|C0034869;C1548330|Quantity limited request - Records;Records|records
Finding|Body Substance|Hospital Course|9497,9504|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|9497,9504|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|9497,9504|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|9514,9522|false|false|false|||refilled
Drug|Organic Chemical|Hospital Course|9523,9528|false|false|false|C0699992|Lasix|lasix
Drug|Pharmacologic Substance|Hospital Course|9523,9528|false|false|false|C0699992|Lasix|lasix
Attribute|Clinical Attribute|Hospital Course|9529,9541|true|false|false|C5886759|Prescription (attribute)|prescription
Event|Event|Hospital Course|9529,9541|false|false|false|||prescription
Finding|Intellectual Product|Hospital Course|9529,9541|true|false|false|C1521941|prescription document|prescription
Procedure|Health Care Activity|Hospital Course|9529,9541|true|false|false|C0033080|Prescription (procedure)|prescription
Finding|Intellectual Product|Hospital Course|9553,9560|false|false|false|C0282416|Overall Publication Type|Overall
Event|Event|Hospital Course|9563,9575|false|false|false|||presentation
Finding|Idea or Concept|Hospital Course|9563,9575|false|false|false|C0449450|Presentation|presentation
Event|Event|Hospital Course|9585,9595|false|false|false|||consistent
Finding|Idea or Concept|Hospital Course|9585,9595|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|Hospital Course|9585,9600|false|false|false|C0332290|Consistent with|consistent with
Finding|Intellectual Product|Hospital Course|9603,9607|false|false|false|C1547225|Mild Severity of Illness Code|mild
Anatomy|Body Space or Junction|Hospital Course|9608,9611|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|Hospital Course|9608,9611|false|false|false|C0018802|Congestive heart failure|CHF
Event|Event|Hospital Course|9612,9624|false|false|false|||exacerbation
Finding|Finding|Hospital Course|9612,9624|false|false|false|C4086268|Exacerbation|exacerbation
Event|Event|Hospital Course|9640,9649|false|false|false|||treatment
Finding|Conceptual Entity|Hospital Course|9640,9649|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Hospital Course|9640,9649|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Hospital Course|9640,9649|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9640,9649|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Drug|Organic Chemical|Hospital Course|9658,9663|false|false|false|C0699992|Lasix|lasix
Drug|Pharmacologic Substance|Hospital Course|9658,9663|false|false|false|C0699992|Lasix|lasix
Event|Event|Hospital Course|9658,9663|false|false|false|||lasix
Event|Event|Hospital Course|9672,9681|false|false|false|||shortness
Attribute|Clinical Attribute|Hospital Course|9672,9691|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|Hospital Course|9672,9691|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|Hospital Course|9685,9691|false|false|false|C0225386|Breath|breath
Event|Event|Hospital Course|9706,9714|false|false|false|||improved
Event|Event|Hospital Course|9732,9736|false|false|false|||able
Finding|Finding|Hospital Course|9732,9736|false|false|false|C1299581|Able (qualifier value)|able
Event|Event|Hospital Course|9743,9755|false|false|false|||transitioned
Event|Event|Hospital Course|9765,9772|false|false|false|||regimen
Finding|Intellectual Product|Hospital Course|9765,9772|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9765,9772|false|false|false|C0040808|Treatment Protocols|regimen
Finding|Idea or Concept|Hospital Course|9800,9803|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|9800,9803|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|9807,9816|false|false|false|||discharge
Finding|Body Substance|Hospital Course|9807,9816|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|9807,9816|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|9807,9816|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|9807,9816|false|false|false|C0030685|Patient Discharge|discharge
Attribute|Clinical Attribute|Hospital Course|9824,9830|false|false|false|C0944911||weight
Event|Event|Hospital Course|9824,9830|false|false|false|||weight
Finding|Finding|Hospital Course|9824,9830|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|Hospital Course|9824,9830|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|Hospital Course|9824,9830|false|false|false|C1305866|Weighing patient|weight
Finding|Idea or Concept|Hospital Course|9834,9837|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|9834,9837|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|9841,9850|false|false|false|||discharge
Finding|Body Substance|Hospital Course|9841,9850|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|9841,9850|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|9841,9850|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|9841,9850|false|false|false|C0030685|Patient Discharge|discharge
Anatomy|Body Location or Region|Hospital Course|9866,9871|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|Hospital Course|9866,9871|false|false|false|C0741025|Chest problem|Chest
Finding|Sign or Symptom|Hospital Course|9866,9881|false|false|false|C0232292|Chest tightness|Chest Tightness
Event|Event|Hospital Course|9872,9881|false|false|false|||Tightness
Finding|Body Substance|Hospital Course|9883,9890|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|9883,9890|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|9883,9890|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|9891,9899|false|false|false|||reported
Anatomy|Body Location or Region|Hospital Course|9900,9905|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|9900,9905|false|false|false|C0741025|Chest problem|chest
Finding|Sign or Symptom|Hospital Course|9900,9915|false|false|false|C0232292|Chest tightness|chest tightness
Event|Event|Hospital Course|9906,9915|false|false|false|||tightness
Event|Event|Hospital Course|9936,9945|false|false|false|||shortness
Finding|Body Substance|Hospital Course|9950,9956|false|false|false|C0225386|Breath|breath
Drug|Organic Chemical|Hospital Course|9968,9975|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|Hospital Course|9968,9975|false|false|false|C0004057|aspirin|aspirin
Event|Event|Hospital Course|9968,9975|false|false|false|||aspirin
Drug|Organic Chemical|Hospital Course|9983,9996|false|false|false|C0017887|nitroglycerin|nitroglycerin
Drug|Pharmacologic Substance|Hospital Course|9983,9996|false|false|false|C0017887|nitroglycerin|nitroglycerin
Event|Event|Hospital Course|9983,9996|false|false|false|||nitroglycerin
Disorder|Disease or Syndrome|Hospital Course|10004,10007|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|Hospital Course|10004,10007|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|Hospital Course|10004,10007|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10004,10007|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|Hospital Course|10004,10007|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|Hospital Course|10004,10007|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|Hospital Course|10004,10007|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|Hospital Course|10004,10007|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|Hospital Course|10004,10007|false|false|false|||PCP
Finding|Gene or Genome|Hospital Course|10004,10007|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|Hospital Course|10004,10007|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|Hospital Course|10011,10017|false|false|false|||office
Finding|Idea or Concept|Hospital Course|10011,10017|false|false|false|C1549636|Address type - Office|office
Event|Event|Hospital Course|10033,10041|false|false|false|||directed
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10053,10061|false|false|false|C0041199|Troponin|Troponin
Drug|Biologically Active Substance|Hospital Course|10053,10061|false|false|false|C0041199|Troponin|Troponin
Event|Event|Hospital Course|10053,10061|false|false|false|||Troponin
Procedure|Laboratory Procedure|Hospital Course|10053,10061|false|false|false|C0523952|Troponin measurement|Troponin
Event|Event|Hospital Course|10066,10074|false|false|false|||negative
Finding|Classification|Hospital Course|10066,10074|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|10066,10074|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|10066,10074|false|false|false|C5237010|Expression Negative|negative
Event|Event|Hospital Course|10080,10083|false|false|false|||EKG
Finding|Intellectual Product|Hospital Course|10080,10083|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|Hospital Course|10080,10083|false|false|false|C1623258|Electrocardiography|EKG
Event|Event|Hospital Course|10092,10100|false|false|false|||evidence
Finding|Idea or Concept|Hospital Course|10092,10100|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Hospital Course|10092,10103|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Finding|Intellectual Product|Hospital Course|10104,10109|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Disease or Syndrome|Hospital Course|10104,10118|true|false|false|C0232353|Acute vascular insufficiency|acute ischemia
Event|Event|Hospital Course|10110,10118|false|false|false|||ischemia
Finding|Pathologic Function|Hospital Course|10110,10118|true|false|false|C0022116|Ischemia|ischemia
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10110,10118|true|false|false|C4321499|Ischemia Procedure|ischemia
Finding|Idea or Concept|Hospital Course|10132,10143|false|false|false|C0750502|Significant|significant
Disorder|Disease or Syndrome|Hospital Course|10144,10147|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10144,10147|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|10144,10147|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Hospital Course|10144,10147|false|false|false|||CAD
Finding|Gene or Genome|Hospital Course|10144,10147|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|10144,10147|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|10144,10147|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10144,10147|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|Hospital Course|10148,10155|false|false|false|||history
Finding|Conceptual Entity|Hospital Course|10148,10155|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|10148,10155|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|10148,10155|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Event|Event|Hospital Course|10161,10170|false|false|false|||underwent
Event|Event|Hospital Course|10175,10179|false|false|false|||MIBI
Procedure|Laboratory Procedure|Hospital Course|10175,10179|false|false|false|C5557372|Multiplexed Ion Beam Imaging|MIBI
Event|Event|Hospital Course|10198,10210|false|false|false|||unremarkable
Anatomy|Body Location or Region|Hospital Course|10216,10221|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|10216,10221|false|false|false|C0741025|Chest problem|chest
Finding|Sign or Symptom|Hospital Course|10216,10231|false|false|false|C0232292|Chest tightness|chest tightness
Event|Event|Hospital Course|10222,10231|false|false|false|||tightness
Event|Event|Hospital Course|10236,10243|false|false|false|||thought
Event|Event|Hospital Course|10266,10274|false|false|false|||etiology
Finding|Conceptual Entity|Hospital Course|10266,10274|false|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|etiology
Finding|Functional Concept|Hospital Course|10266,10274|false|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|etiology
Disorder|Disease or Syndrome|Hospital Course|10279,10282|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|Hospital Course|10279,10282|false|false|false|||HTN
Finding|Body Substance|Hospital Course|10284,10291|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|10284,10291|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|10284,10291|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|10292,10301|false|false|false|||presented
Attribute|Clinical Attribute|Hospital Course|10307,10310|false|false|false|C0871470|Systolic Pressure|SBP
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10307,10310|false|false|false|C0085805|Androgen Binding Protein|SBP
Drug|Biologically Active Substance|Hospital Course|10307,10310|false|false|false|C0085805|Androgen Binding Protein|SBP
Event|Event|Hospital Course|10307,10310|false|false|false|||SBP
Finding|Gene or Genome|Hospital Course|10307,10310|false|false|false|C1705296;C3274833|CCHCR1 wt Allele;SHBG wt Allele|SBP
Procedure|Diagnostic Procedure|Hospital Course|10307,10310|false|false|false|C1306620|Systolic blood pressure measurement|SBP
Anatomy|Body System|Hospital Course|10323,10333|false|false|false|C0007226|Cardiovascular system|Cardiology
Event|Event|Hospital Course|10338,10347|false|false|false|||consulted
Event|Event|Hospital Course|10353,10364|false|false|false|||recommended
Event|Event|Hospital Course|10365,10375|false|false|false|||increasing
Drug|Organic Chemical|Hospital Course|10380,10390|false|false|false|C0054836|carvedilol|carvedilol
Drug|Pharmacologic Substance|Hospital Course|10380,10390|false|false|false|C0054836|carvedilol|carvedilol
Event|Event|Hospital Course|10380,10390|false|false|false|||carvedilol
Disorder|Mental or Behavioral Dysfunction|Hospital Course|10403,10406|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10403,10406|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|10403,10406|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|10403,10406|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|10403,10406|false|false|false|C1332410|BID gene|BID
Disorder|Mental or Behavioral Dysfunction|Hospital Course|10418,10421|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10418,10421|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|10418,10421|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|10418,10421|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|10418,10421|false|false|false|C1332410|BID gene|BID
Event|Event|Hospital Course|10433,10439|false|false|false|||change
Finding|Functional Concept|Hospital Course|10433,10439|false|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10433,10439|false|false|false|C4319952|Change - procedure|change
Event|Event|Hospital Course|10445,10457|false|false|false|||continuation
Event|Event|Hospital Course|10471,10475|false|false|false|||home
Finding|Idea or Concept|Hospital Course|10471,10475|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|10471,10475|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|10471,10475|false|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|Hospital Course|10477,10488|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Hospital Course|10477,10488|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Hospital Course|10477,10488|false|false|false|||medications
Finding|Intellectual Product|Hospital Course|10477,10488|false|false|false|C4284232|Medications|medications
Disorder|Disease or Syndrome|Hospital Course|10494,10499|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Hospital Course|10494,10499|false|false|false|||blood
Finding|Body Substance|Hospital Course|10494,10499|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|Hospital Course|10494,10508|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Finding|Organism Function|Hospital Course|10494,10508|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Procedure|Health Care Activity|Hospital Course|10494,10508|false|false|false|C0005824|Blood pressure determination|blood pressure
Event|Event|Hospital Course|10500,10508|false|false|false|||pressure
Finding|Finding|Hospital Course|10500,10508|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|Hospital Course|10500,10508|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|Hospital Course|10500,10508|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|Hospital Course|10500,10508|false|false|false|C0033095||pressure
Event|Event|Hospital Course|10509,10518|false|false|false|||decreased
Event|Event|Hospital Course|10522,10531|false|false|false|||systolics
Event|Event|Hospital Course|10535,10540|false|false|false|||range
Finding|Intellectual Product|Hospital Course|10535,10540|false|false|false|C3542016|Concept model range (foundation metadata concept)|range
Finding|Idea or Concept|Hospital Course|10556,10559|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|10556,10559|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|10563,10572|false|false|false|||discharge
Finding|Body Substance|Hospital Course|10563,10572|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|10563,10572|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|10563,10572|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|10563,10572|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|Hospital Course|10580,10587|false|false|false|||unclear
Finding|Finding|Hospital Course|10606,10617|false|false|false|C0497247|Increase in blood pressure|elevated BP
Event|Event|Hospital Course|10615,10617|false|false|false|||BP
Event|Event|Hospital Course|10621,10630|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|10621,10630|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|Hospital Course|10635,10644|false|false|false|||occurring
Finding|Mental Process|Hospital Course|10652,10659|false|false|false|C0542559|contextual factors|setting
Drug|Pharmacologic Substance|Hospital Course|10664,10674|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Hospital Course|10664,10674|false|false|false|||medication
Finding|Intellectual Product|Hospital Course|10664,10674|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Finding|Individual Behavior|Hospital Course|10664,10689|false|false|false|C3489773|Medication Compliance|medication non-compliance
Event|Event|Hospital Course|10675,10689|false|false|false|||non-compliance
Drug|Organic Chemical|Hospital Course|10691,10701|false|false|false|C0028066|nifedipine|Nifedipine
Drug|Pharmacologic Substance|Hospital Course|10691,10701|false|false|false|C0028066|nifedipine|Nifedipine
Event|Event|Hospital Course|10691,10701|false|false|false|||Nifedipine
Event|Event|Hospital Course|10706,10715|false|false|false|||decreased
Disorder|Mental or Behavioral Dysfunction|Hospital Course|10721,10724|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10721,10724|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|10721,10724|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|10721,10724|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|10721,10724|false|false|false|C1332410|BID gene|BID
Event|Event|Hospital Course|10741,10750|false|false|false|||increased
Drug|Organic Chemical|Hospital Course|10751,10761|false|false|false|C0054836|carvedilol|carvedilol
Drug|Pharmacologic Substance|Hospital Course|10751,10761|false|false|false|C0054836|carvedilol|carvedilol
Event|Event|Hospital Course|10751,10761|false|false|false|||carvedilol
Event|Event|Hospital Course|10766,10774|false|false|false|||addition
Finding|Functional Concept|Hospital Course|10766,10774|false|false|false|C0332287;C1883712|Add - instruction imperative;In addition to|addition
Drug|Organic Chemical|Hospital Course|10778,10783|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|Hospital Course|10778,10783|false|false|false|C0699992|Lasix|Lasix
Event|Event|Hospital Course|10778,10783|false|false|false|||Lasix
Finding|Body Substance|Hospital Course|10792,10799|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|10792,10799|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|10792,10799|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|10804,10812|false|false|false|||believed
Event|Event|Hospital Course|10826,10839|false|false|false|||non-compliant
Event|Event|Hospital Course|10860,10869|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|10860,10869|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Idea or Concept|Hospital Course|10878,10890|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Anatomy|Body Space or Junction|Hospital Course|10906,10909|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|Hospital Course|10906,10909|false|false|false|C0018802|Congestive heart failure|CHF
Event|Event|Hospital Course|10906,10909|false|false|false|||CHF
Event|Event|Hospital Course|10917,10925|false|false|false|||services
Event|Occupational Activity|Hospital Course|10917,10925|false|false|false|C0557854|Services|services
Procedure|Health Care Activity|Hospital Course|10917,10925|false|false|false|C1704289|Clinical Service|services
Drug|Pharmacologic Substance|Hospital Course|10930,10940|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Hospital Course|10930,10940|false|false|false|||medication
Finding|Intellectual Product|Hospital Course|10930,10940|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Hospital Course|10941,10949|false|false|false|||teaching
Finding|Intellectual Product|Hospital Course|10941,10949|false|false|false|C1548344|Visit User Code - Teaching|teaching
Procedure|Educational Activity|Hospital Course|10941,10949|false|false|false|C0039401;C0220924|Education (procedure);Teaching aspects|teaching
Drug|Biomedical or Dental Material|Hospital Course|10954,10958|false|false|false|C0009905;C0994475|Contraceptives, Oral;Pills|pill
Drug|Pharmacologic Substance|Hospital Course|10954,10958|false|false|false|C0009905;C0994475|Contraceptives, Oral;Pills|pill
Event|Event|Hospital Course|10954,10958|false|false|false|||pill
Event|Event|Hospital Course|10959,10962|false|false|false|||box
Finding|Idea or Concept|Hospital Course|10959,10962|false|false|false|C1552831|Table Frame - box|box
Finding|Finding|Hospital Course|10967,10971|false|false|false|C5575035|Well (answer to question)|well
Event|Event|Hospital Course|10976,10983|false|false|false|||weights
Finding|Daily or Recreational Activity|Hospital Course|10976,10983|false|false|false|C3812400|Weights - exercise activity|weights
Finding|Functional Concept|Hospital Course|10986,10992|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|Follow
Finding|Intellectual Product|Hospital Course|10986,10992|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|Follow
Finding|Finding|Hospital Course|10986,10995|false|false|false|C0589120|Follow-up status|Follow up
Procedure|Health Care Activity|Hospital Course|10986,10995|false|false|false|C1522577|follow-up|Follow up
Event|Event|Hospital Course|10993,10995|false|false|false|||up
Event|Event|Hospital Course|11042,11047|false|false|false|||check
Finding|Functional Concept|Hospital Course|11048,11054|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Event|Event|Hospital Course|11055,11059|false|false|false|||Chem
Finding|Functional Concept|Hospital Course|11055,11059|false|false|false|C0079107|chemical aspects|Chem
Procedure|Laboratory Procedure|Hospital Course|11055,11059|false|false|false|C0201682|Chemical procedure|Chem
Anatomy|Cell Component|Hospital Course|11067,11070|false|false|false|C2263086|Nuclear cap binding complex location|CBC
Procedure|Laboratory Procedure|Hospital Course|11067,11070|false|false|false|C0009555|Complete Blood Count|CBC
Event|Event|Hospital Course|11080,11088|false|false|false|||Continue
Drug|Organic Chemical|Hospital Course|11089,11099|false|false|false|C0016860|furosemide|furosemide
Drug|Pharmacologic Substance|Hospital Course|11089,11099|false|false|false|C0016860|furosemide|furosemide
Procedure|Laboratory Procedure|Hospital Course|11113,11116|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11113,11116|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Drug|Biomedical or Dental Material|Hospital Course|11117,11121|false|false|false|C0991568|Drops - Drug Form|Drop
Event|Activity|Hospital Course|11117,11121|false|false|false|C1705648|Dropping|Drop
Event|Event|Hospital Course|11117,11121|false|false|false|||Drop
Finding|Body Substance|Hospital Course|11123,11130|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|11123,11130|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|11123,11130|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|11136,11143|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Hospital Course|11136,11143|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|Hospital Course|11136,11150|false|false|false|C0581384|Chronic anemia|chronic anemia
Disorder|Disease or Syndrome|Hospital Course|11144,11150|false|false|false|C0002871|Anemia|anemia
Event|Event|Hospital Course|11144,11150|false|false|false|||anemia
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11155,11158|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Hospital Course|11155,11158|false|false|false|C0019046|Hemoglobin|Hgb
Event|Event|Hospital Course|11155,11158|false|false|false|||Hgb
Finding|Gene or Genome|Hospital Course|11155,11158|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Hospital Course|11155,11158|false|false|false|C0019029|Hemoglobin concentration|Hgb
Drug|Biomedical or Dental Material|Hospital Course|11159,11163|false|false|false|C0991568|Drops - Drug Form|drop
Event|Activity|Hospital Course|11159,11163|false|false|false|C1705648|Dropping|drop
Finding|Idea or Concept|Hospital Course|11167,11170|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|11167,11170|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|11175,11184|false|false|false|||discharge
Finding|Body Substance|Hospital Course|11175,11184|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|11175,11184|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|11175,11184|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|11175,11184|false|false|false|C0030685|Patient Discharge|discharge
Finding|Functional Concept|Hospital Course|11204,11210|false|false|false|C0205341;C1705914|Repeat;Repeat Object|Repeat
Anatomy|Cell Component|Hospital Course|11211,11214|false|false|false|C2263086|Nuclear cap binding complex location|CBC
Procedure|Laboratory Procedure|Hospital Course|11211,11214|false|false|false|C0009555|Complete Blood Count|CBC
Event|Activity|Hospital Course|11215,11220|false|false|false|C1283174||check
Event|Event|Hospital Course|11215,11220|false|false|false|||check
Finding|Functional Concept|Hospital Course|11215,11220|false|false|false|C4321547|Check|check
Disorder|Disease or Syndrome|Hospital Course|11231,11234|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|Hospital Course|11231,11234|false|false|false|||HTN
Event|Event|Hospital Course|11238,11247|false|false|false|||Increased
Drug|Organic Chemical|Hospital Course|11248,11258|false|false|false|C0054836|carvedilol|carvedilol
Drug|Pharmacologic Substance|Hospital Course|11248,11258|false|false|false|C0054836|carvedilol|carvedilol
Event|Event|Hospital Course|11248,11258|false|false|false|||carvedilol
Disorder|Mental or Behavioral Dysfunction|Hospital Course|11269,11272|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11269,11272|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|11269,11272|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|11269,11272|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|11269,11272|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|11275,11285|false|false|false|C0028066|nifedipine|Nifedipine
Drug|Pharmacologic Substance|Hospital Course|11275,11285|false|false|false|C0028066|nifedipine|Nifedipine
Event|Event|Hospital Course|11275,11285|false|false|false|||Nifedipine
Event|Event|Hospital Course|11290,11299|false|false|false|||decreased
Disorder|Mental or Behavioral Dysfunction|Hospital Course|11305,11308|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11305,11308|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|11305,11308|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|11305,11308|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|11305,11308|false|false|false|C1332410|BID gene|BID
Event|Event|Hospital Course|11324,11333|false|false|false|||increased
Drug|Organic Chemical|Hospital Course|11335,11345|false|false|false|C0054836|carvedilol|carvedilol
Drug|Pharmacologic Substance|Hospital Course|11335,11345|false|false|false|C0054836|carvedilol|carvedilol
Event|Event|Hospital Course|11335,11345|false|false|false|||carvedilol
Event|Event|Hospital Course|11350,11358|false|false|false|||addition
Finding|Functional Concept|Hospital Course|11350,11358|false|false|false|C0332287;C1883712|Add - instruction imperative;In addition to|addition
Drug|Organic Chemical|Hospital Course|11362,11367|false|false|false|C0699992|Lasix|lasix
Drug|Pharmacologic Substance|Hospital Course|11362,11367|false|false|false|C0699992|Lasix|lasix
Event|Event|Hospital Course|11362,11367|false|false|false|||lasix
Finding|Body Substance|Hospital Course|11380,11387|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|11380,11387|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|11380,11387|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|Hospital Course|11392,11398|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|11392,11398|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|Hospital Course|11428,11437|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|11428,11437|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Idea or Concept|Hospital Course|11443,11449|false|false|false|C0018684|Health|Health
Procedure|Diagnostic Procedure|Hospital Course|11443,11459|false|false|false|C0220908|Screening procedure|Health Screening
Event|Event|Hospital Course|11450,11459|false|false|false|||Screening
Finding|Finding|Hospital Course|11450,11459|false|false|false|C0220909;C1305399;C1409616|Aspects of disease screening;Screening - procedure intent;Special screening finding|Screening
Finding|Functional Concept|Hospital Course|11450,11459|false|false|false|C0220909;C1305399;C1409616|Aspects of disease screening;Screening - procedure intent;Special screening finding|Screening
Procedure|Diagnostic Procedure|Hospital Course|11450,11459|false|false|false|C0199230;C0220908;C1698960;C1710031;C1710032|Disease Screening;Screening;Screening for cancer;Screening procedure;research subject screening|Screening
Procedure|Health Care Activity|Hospital Course|11450,11459|false|false|false|C0199230;C0220908;C1698960;C1710031;C1710032|Disease Screening;Screening;Screening for cancer;Screening procedure;research subject screening|Screening
Procedure|Research Activity|Hospital Course|11450,11459|false|false|false|C0199230;C0220908;C1698960;C1710031;C1710032|Disease Screening;Screening;Screening for cancer;Screening procedure;research subject screening|Screening
Finding|Body Substance|Hospital Course|11462,11469|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|11462,11469|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|11462,11469|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|11481,11492|false|false|false|||colonoscopy
Procedure|Diagnostic Procedure|Hospital Course|11481,11492|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Procedure|Health Care Activity|Hospital Course|11481,11492|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Finding|Idea or Concept|Hospital Course|11498,11502|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|Hospital Course|11498,11502|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Disorder|Disease or Syndrome|Hospital Course|11506,11509|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|Hospital Course|11506,11509|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|Hospital Course|11506,11509|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11506,11509|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|Hospital Course|11506,11509|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|Hospital Course|11506,11509|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|Hospital Course|11506,11509|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|Hospital Course|11506,11509|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|Hospital Course|11506,11509|false|false|false|||PCP
Finding|Gene or Genome|Hospital Course|11506,11509|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|Hospital Course|11506,11509|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|Hospital Course|11510,11516|false|false|false|||follow
Finding|Functional Concept|Hospital Course|11510,11516|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|Hospital Course|11510,11516|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|Hospital Course|11510,11519|false|false|false|C0589120|Follow-up status|follow up
Procedure|Health Care Activity|Hospital Course|11510,11519|false|false|false|C1522577|follow-up|follow up
Event|Event|Hospital Course|11517,11519|false|false|false|||up
Attribute|Clinical Attribute|Hospital Course|11543,11549|false|false|false|C0944911||Weight
Event|Event|Hospital Course|11543,11549|false|false|false|||Weight
Finding|Finding|Hospital Course|11543,11549|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|Weight
Finding|Sign or Symptom|Hospital Course|11543,11549|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|Weight
Procedure|Health Care Activity|Hospital Course|11543,11549|false|false|false|C1305866|Weighing patient|Weight
Event|Event|Hospital Course|11553,11562|false|false|false|||discharge
Finding|Body Substance|Hospital Course|11553,11562|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|11553,11562|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|11553,11562|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|11553,11562|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|Hospital Course|11575,11579|false|false|false|||Code
Event|Occupational Activity|Hospital Course|11575,11579|false|false|false|C0009219|Coding|Code
Finding|Intellectual Product|Hospital Course|11575,11579|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|Code
Event|Event|Hospital Course|11587,11596|false|false|false|||confirmed
Finding|Body Substance|Hospital Course|11602,11609|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|11602,11609|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|11602,11609|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|11613,11622|false|false|false|||Emergency
Finding|Finding|Hospital Course|11613,11622|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Idea or Concept|Hospital Course|11613,11622|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Intellectual Product|Hospital Course|11613,11622|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Pathologic Function|Hospital Course|11613,11622|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Phenomenon|Phenomenon or Process|Hospital Course|11613,11622|false|false|false|C0013956|Emergency Situation|Emergency
Procedure|Health Care Activity|Hospital Course|11613,11622|false|false|false|C1553500|emergency encounter|Emergency
Event|Event|Hospital Course|11623,11631|false|false|false|||Contacts
Procedure|Health Care Activity|Hospital Course|11623,11631|false|false|false|C4036459|Contacts|Contacts
Finding|Functional Concept|Hospital Course|11652,11661|false|false|false|C0332270;C1552848|Alternating;alternate - HtmlLinkType|Alternate
Finding|Idea or Concept|Hospital Course|11652,11661|false|false|false|C0332270;C1552848|Alternating;alternate - HtmlLinkType|Alternate
Disorder|Disease or Syndrome|Hospital Course|11662,11665|false|false|false|C0162531|Hereditary Coproporphyria|HCP
Event|Event|Hospital Course|11662,11665|false|false|false|||HCP
Finding|Gene or Genome|Hospital Course|11662,11665|false|false|false|C1335283;C1412376;C1413681;C1705637;C5780748|AMBP gene;AMBP wt Allele;CPOX gene;PTPN6 gene;PTPN6 wt Allele|HCP
Attribute|Clinical Attribute|Hospital Course|11676,11687|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|11676,11687|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|11676,11687|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|11676,11687|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|11676,11700|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|11691,11700|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|11691,11700|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|Hospital Course|11719,11729|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Hospital Course|11719,11729|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|Hospital Course|11719,11734|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|Hospital Course|11730,11734|false|false|false|||list
Finding|Intellectual Product|Hospital Course|11730,11734|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|Hospital Course|11738,11746|false|false|false|||accurate
Drug|Organic Chemical|Hospital Course|11751,11759|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Hospital Course|11751,11759|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Hospital Course|11751,11759|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|Hospital Course|11751,11759|false|false|false|||complete
Finding|Functional Concept|Hospital Course|11751,11759|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|11751,11759|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|Hospital Course|11764,11771|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Hospital Course|11764,11771|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|Hospital Course|11791,11802|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Pharmacologic Substance|Hospital Course|11791,11802|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Organic Chemical|Hospital Course|11822,11832|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|Hospital Course|11822,11832|false|false|false|C0016860|furosemide|Furosemide
Drug|Organic Chemical|Hospital Course|11852,11865|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|Hospital Course|11852,11865|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|Hospital Course|11852,11865|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Event|Event|Hospital Course|11852,11865|false|false|false|||Multivitamins
Drug|Biomedical or Dental Material|Hospital Course|11868,11871|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|Hospital Course|11868,11871|false|false|false|||TAB
Drug|Organic Chemical|Hospital Course|11885,11895|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Pharmacologic Substance|Hospital Course|11885,11895|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Organic Chemical|Hospital Course|11916,11928|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|11916,11928|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11948,11955|false|false|false|C0020171;C0020172;C3538423|Humulin;Humulin S;Humulin insulin|HumuLIN
Drug|Hormone|Hospital Course|11948,11955|false|false|false|C0020171;C0020172;C3538423|Humulin;Humulin S;Humulin insulin|HumuLIN
Drug|Pharmacologic Substance|Hospital Course|11948,11955|false|false|false|C0020171;C0020172;C3538423|Humulin;Humulin S;Humulin insulin|HumuLIN
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11948,11961|false|false|false|C0306367|HumuLIN 70/30|HumuLIN 70/30
Drug|Hormone|Hospital Course|11948,11961|false|false|false|C0306367|HumuLIN 70/30|HumuLIN 70/30
Drug|Pharmacologic Substance|Hospital Course|11948,11961|false|false|false|C0306367|HumuLIN 70/30|HumuLIN 70/30
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11963,11970|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|Hospital Course|11963,11970|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|Hospital Course|11963,11970|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|Hospital Course|11963,11970|false|false|false|||insulin
Finding|Gene or Genome|Hospital Course|11963,11970|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|Hospital Course|11963,11970|false|false|false|C0202098|Insulin measurement|insulin
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11963,11974|false|false|false|C0021658|insulin isophane|insulin NPH
Drug|Hormone|Hospital Course|11963,11974|false|false|false|C0021658|insulin isophane|insulin NPH
Drug|Pharmacologic Substance|Hospital Course|11963,11974|false|false|false|C0021658|insulin isophane|insulin NPH
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11971,11974|false|false|false|C0027442|Nasopharynx|NPH
Disorder|Disease or Syndrome|Hospital Course|11971,11974|false|false|false|C0020258|Hydrocephalus, Normal Pressure|NPH
Event|Event|Hospital Course|11971,11974|false|false|false|||NPH
Finding|Functional Concept|Hospital Course|12004,12016|false|false|false|C1522438|Subcutaneous Route of Administration|subcutaneous
Drug|Organic Chemical|Hospital Course|12027,12040|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Pharmacologic Substance|Hospital Course|12027,12040|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Event|Event|Hospital Course|12027,12040|false|false|false|||Nitroglycerin
Finding|Gene or Genome|Hospital Course|12054,12057|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Location or Region|Hospital Course|12058,12063|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|12058,12063|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|12058,12068|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Hospital Course|12058,12068|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Hospital Course|12064,12068|false|true|false|C2598155||pain
Event|Event|Hospital Course|12064,12068|false|false|false|||pain
Finding|Functional Concept|Hospital Course|12064,12068|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|12064,12068|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|12073,12080|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|12073,12080|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|12073,12080|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|Hospital Course|12073,12082|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|Hospital Course|12073,12082|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|Hospital Course|12073,12082|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|Hospital Course|12073,12082|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|Hospital Course|12073,12082|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|Hospital Course|12081,12082|false|false|false|||D
Event|Event|Hospital Course|12087,12091|false|false|false|||UNIT
Drug|Organic Chemical|Hospital Course|12106,12116|false|false|false|C0028066|nifedipine|NIFEdipine
Drug|Pharmacologic Substance|Hospital Course|12106,12116|false|false|false|C0028066|nifedipine|NIFEdipine
Event|Event|Hospital Course|12106,12116|false|false|false|||NIFEdipine
Disorder|Mental or Behavioral Dysfunction|Hospital Course|12129,12132|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12129,12132|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|12129,12132|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|12129,12132|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|12129,12132|false|false|false|C1332410|BID gene|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12138,12148|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|Hospital Course|12138,12148|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Organic Chemical|Hospital Course|12169,12180|false|false|false|C0002144|allopurinol|Allopurinol
Drug|Pharmacologic Substance|Hospital Course|12169,12180|false|false|false|C0002144|allopurinol|Allopurinol
Drug|Element, Ion, or Isotope|Hospital Course|12202,12209|false|false|false|C2346592|Ferrous|Ferrous
Drug|Inorganic Chemical|Hospital Course|12202,12217|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Pharmacologic Substance|Hospital Course|12202,12217|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Element, Ion, or Isotope|Hospital Course|12210,12217|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Inorganic Chemical|Hospital Course|12210,12217|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Pharmacologic Substance|Hospital Course|12210,12217|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Event|Event|Hospital Course|12210,12217|false|false|false|||Sulfate
Drug|Organic Chemical|Hospital Course|12239,12249|false|false|false|C0054836|carvedilol|Carvedilol
Drug|Pharmacologic Substance|Hospital Course|12239,12249|false|false|false|C0054836|carvedilol|Carvedilol
Disorder|Mental or Behavioral Dysfunction|Hospital Course|12261,12264|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12261,12264|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|12261,12264|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|12261,12264|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|12261,12264|false|false|false|C1332410|BID gene|BID
Event|Event|Hospital Course|12269,12278|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|12269,12278|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|12269,12278|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|12269,12278|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|12269,12278|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|12269,12290|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|12279,12290|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|12279,12290|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|12279,12290|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|12279,12290|false|false|false|C4284232|Medications|Medications
Finding|Classification|Hospital Course|12295,12305|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|Outpatient
Finding|Idea or Concept|Hospital Course|12295,12305|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|Outpatient
Finding|Gene or Genome|Hospital Course|12306,12309|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|Lab
Finding|Intellectual Product|Hospital Course|12306,12309|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|Lab
Event|Event|Hospital Course|12310,12314|false|false|false|||Work
Event|Occupational Activity|Hospital Course|12310,12314|false|false|false|C0043227|Work|Work
Event|Event|Hospital Course|12327,12331|false|false|false|||Chem
Finding|Functional Concept|Hospital Course|12327,12331|false|false|false|C0079107|chemical aspects|Chem
Procedure|Laboratory Procedure|Hospital Course|12327,12331|false|false|false|C0201682|Chemical procedure|Chem
Anatomy|Cell Component|Hospital Course|12339,12342|false|false|false|C2263086|Nuclear cap binding complex location|CBC
Procedure|Laboratory Procedure|Hospital Course|12339,12342|false|false|false|C0009555|Complete Blood Count|CBC
Attribute|Clinical Attribute|Hospital Course|12351,12361|false|false|false|C5890010||Indication
Event|Event|Hospital Course|12351,12361|false|false|false|||Indication
Finding|Idea or Concept|Hospital Course|12351,12361|false|false|false|C0392360;C3146298|Indication;Indication of (contextual qualifier)|Indication
Anatomy|Body Space or Junction|Hospital Course|12370,12373|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|Hospital Course|12370,12373|false|false|false|C0018802|Congestive heart failure|CHF
Disorder|Disease or Syndrome|Hospital Course|12379,12385|false|false|false|C0002871|Anemia|anemia
Event|Event|Hospital Course|12379,12385|false|false|false|||anemia
Event|Event|Hospital Course|12399,12406|false|false|false|||results
Finding|Idea or Concept|Hospital Course|12419,12422|false|false|false|C1547563;C1549619|Authorization Mode - Fax;Fax Number|fax
Finding|Intellectual Product|Hospital Course|12419,12422|false|false|false|C1547563;C1549619|Authorization Mode - Fax;Fax Number|fax
Drug|Organic Chemical|Hospital Course|12431,12444|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Pharmacologic Substance|Hospital Course|12431,12444|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Event|Event|Hospital Course|12431,12444|false|false|false|||Nitroglycerin
Finding|Gene or Genome|Hospital Course|12458,12461|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Location or Region|Hospital Course|12462,12467|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|12462,12467|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|12462,12472|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Hospital Course|12462,12472|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Hospital Course|12468,12472|false|true|false|C2598155||pain
Event|Event|Hospital Course|12468,12472|false|false|false|||pain
Finding|Functional Concept|Hospital Course|12468,12472|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|12468,12472|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|12477,12484|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|12477,12484|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|12477,12484|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|Hospital Course|12477,12486|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|Hospital Course|12477,12486|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|Hospital Course|12477,12486|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|Hospital Course|12477,12486|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|Hospital Course|12477,12486|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|Hospital Course|12485,12486|false|false|false|||D
Event|Event|Hospital Course|12491,12495|false|false|false|||UNIT
Drug|Organic Chemical|Hospital Course|12509,12519|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Pharmacologic Substance|Hospital Course|12509,12519|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Organic Chemical|Hospital Course|12540,12550|false|false|false|C0028066|nifedipine|NIFEdipine
Drug|Pharmacologic Substance|Hospital Course|12540,12550|false|false|false|C0028066|nifedipine|NIFEdipine
Event|Event|Hospital Course|12540,12550|false|false|false|||NIFEdipine
Drug|Organic Chemical|Hospital Course|12573,12586|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|Hospital Course|12573,12586|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|Hospital Course|12573,12586|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Event|Event|Hospital Course|12573,12586|false|false|false|||Multivitamins
Drug|Biomedical or Dental Material|Hospital Course|12589,12592|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|Hospital Course|12589,12592|false|false|false|||TAB
Drug|Organic Chemical|Hospital Course|12606,12617|false|false|false|C0002144|allopurinol|Allopurinol
Drug|Pharmacologic Substance|Hospital Course|12606,12617|false|false|false|C0002144|allopurinol|Allopurinol
Drug|Organic Chemical|Hospital Course|12638,12645|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Hospital Course|12638,12645|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|Hospital Course|12665,12677|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|12665,12677|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|Hospital Course|12698,12709|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Pharmacologic Substance|Hospital Course|12698,12709|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Element, Ion, or Isotope|Hospital Course|12730,12737|false|false|false|C2346592|Ferrous|Ferrous
Drug|Inorganic Chemical|Hospital Course|12730,12745|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Pharmacologic Substance|Hospital Course|12730,12745|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Element, Ion, or Isotope|Hospital Course|12738,12745|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Inorganic Chemical|Hospital Course|12738,12745|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Pharmacologic Substance|Hospital Course|12738,12745|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Event|Event|Hospital Course|12738,12745|false|false|false|||Sulfate
Drug|Organic Chemical|Hospital Course|12767,12777|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|Hospital Course|12767,12777|false|false|false|C0016860|furosemide|Furosemide
Event|Event|Hospital Course|12794,12796|false|false|false|||RX
Drug|Organic Chemical|Hospital Course|12798,12808|false|false|false|C0016860|furosemide|furosemide
Drug|Pharmacologic Substance|Hospital Course|12798,12808|false|false|false|C0016860|furosemide|furosemide
Event|Event|Hospital Course|12798,12808|false|false|false|||furosemide
Drug|Biomedical or Dental Material|Hospital Course|12817,12823|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|12827,12835|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|12830,12835|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|12830,12835|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Biomedical or Dental Material|Hospital Course|12851,12857|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|12851,12857|false|false|false|||Tablet
Event|Event|Hospital Course|12859,12866|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|12859,12866|false|false|false|C0807726|refill|Refills
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12874,12881|false|false|false|C0020171;C0020172;C3538423|Humulin;Humulin S;Humulin insulin|HumuLIN
Drug|Hormone|Hospital Course|12874,12881|false|false|false|C0020171;C0020172;C3538423|Humulin;Humulin S;Humulin insulin|HumuLIN
Drug|Pharmacologic Substance|Hospital Course|12874,12881|false|false|false|C0020171;C0020172;C3538423|Humulin;Humulin S;Humulin insulin|HumuLIN
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12874,12887|false|false|false|C0306367|HumuLIN 70/30|HumuLIN 70/30
Drug|Hormone|Hospital Course|12874,12887|false|false|false|C0306367|HumuLIN 70/30|HumuLIN 70/30
Drug|Pharmacologic Substance|Hospital Course|12874,12887|false|false|false|C0306367|HumuLIN 70/30|HumuLIN 70/30
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12889,12896|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|Hospital Course|12889,12896|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|Hospital Course|12889,12896|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|Hospital Course|12889,12896|false|false|false|||insulin
Finding|Gene or Genome|Hospital Course|12889,12896|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|Hospital Course|12889,12896|false|false|false|C0202098|Insulin measurement|insulin
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12889,12900|false|false|false|C0021658|insulin isophane|insulin NPH
Drug|Hormone|Hospital Course|12889,12900|false|false|false|C0021658|insulin isophane|insulin NPH
Drug|Pharmacologic Substance|Hospital Course|12889,12900|false|false|false|C0021658|insulin isophane|insulin NPH
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12897,12900|false|false|false|C0027442|Nasopharynx|NPH
Disorder|Disease or Syndrome|Hospital Course|12897,12900|false|false|false|C0020258|Hydrocephalus, Normal Pressure|NPH
Event|Event|Hospital Course|12897,12900|false|false|false|||NPH
Finding|Functional Concept|Hospital Course|12930,12942|false|false|false|C1522438|Subcutaneous Route of Administration|subcutaneous
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12954,12964|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|Hospital Course|12954,12964|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Organic Chemical|Hospital Course|12985,12995|false|false|false|C0054836|carvedilol|Carvedilol
Drug|Pharmacologic Substance|Hospital Course|12985,12995|false|false|false|C0054836|carvedilol|Carvedilol
Disorder|Mental or Behavioral Dysfunction|Hospital Course|13007,13010|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|13007,13010|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|13007,13010|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|13007,13010|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|13007,13010|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|13016,13026|false|false|false|C0054836|carvedilol|carvedilol
Drug|Pharmacologic Substance|Hospital Course|13016,13026|false|false|false|C0054836|carvedilol|carvedilol
Event|Event|Hospital Course|13016,13026|false|false|false|||carvedilol
Drug|Biomedical or Dental Material|Hospital Course|13037,13043|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|13047,13055|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|13050,13055|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|13050,13055|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|Hospital Course|13064,13067|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|13064,13067|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Activity|Hospital Course|13068,13072|false|false|false|C1880359|Dispense (activity)|Disp
Finding|Gene or Genome|Hospital Course|13068,13072|false|false|false|C2828567|PRSS30P gene|Disp
Drug|Biomedical or Dental Material|Hospital Course|13079,13085|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|13086,13093|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|13086,13093|false|false|false|C0807726|refill|Refills
Event|Event|Hospital Course|13100,13109|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|13100,13109|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|13100,13109|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|13100,13109|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|13100,13109|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|13100,13121|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|13100,13121|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|13110,13121|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|13110,13121|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|13110,13121|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|Hospital Course|13123,13127|false|false|false|||Home
Finding|Idea or Concept|Hospital Course|13123,13127|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|13123,13127|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|13123,13127|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|Hospital Course|13133,13140|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|Hospital Course|13133,13140|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|Hospital Course|13143,13151|false|false|false|||Facility
Finding|Intellectual Product|Hospital Course|13143,13151|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|Hospital Course|13159,13168|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|13159,13168|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|13159,13168|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|13159,13168|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|13159,13168|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|13159,13178|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|13169,13178|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|13169,13178|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|13169,13178|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|13169,13178|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|13169,13178|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Intellectual Product|Principle Diagnosis|13201,13206|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Finding|Intellectual Product|Principle Diagnosis|13210,13217|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Principle Diagnosis|13210,13217|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Finding|Organ or Tissue Function|Principle Diagnosis|13232,13240|false|false|false|C0039155|Systole|systolic
Disorder|Disease or Syndrome|Principle Diagnosis|13232,13254|false|false|false|C1135191|Heart Failure, Systolic|systolic heart failure
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|13241,13246|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Principle Diagnosis|13241,13246|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Principle Diagnosis|13241,13246|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|Principle Diagnosis|13241,13254|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Event|Event|Principle Diagnosis|13247,13254|false|false|false|||failure
Finding|Functional Concept|Principle Diagnosis|13247,13254|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|Principle Diagnosis|13247,13254|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|Principle Diagnosis|13247,13254|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Mental Process|Discharge Condition|13279,13285|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|13279,13292|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|13279,13292|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|13286,13292|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|13286,13292|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|13294,13299|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|13294,13299|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|13304,13312|false|false|false|||coherent
Finding|Finding|Discharge Condition|13304,13312|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|13314,13319|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|13314,13336|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|13314,13336|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|13323,13336|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|13323,13336|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|13323,13336|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|13338,13343|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|13338,13343|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|13338,13343|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|13338,13343|false|false|false|||Alert
Finding|Finding|Discharge Condition|13338,13343|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|13338,13343|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|13338,13343|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|13348,13359|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|13348,13359|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|13361,13369|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|13361,13369|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|13361,13369|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|13370,13376|false|false|false|C5889824||Status
Event|Event|Discharge Condition|13370,13376|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|13370,13376|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|13378,13388|false|false|false|||Ambulatory
Finding|Functional Concept|Discharge Condition|13378,13388|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|13378,13388|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|13378,13388|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|13378,13388|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|13391,13402|false|false|false|||Independent
Finding|Finding|Discharge Condition|13391,13402|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Condition|13391,13402|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Gene or Genome|Discharge Instructions|13431,13435|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|Discharge Instructions|13451,13459|false|false|false|||admitted
Event|Event|Discharge Instructions|13479,13488|false|false|false|||shortness
Attribute|Clinical Attribute|Discharge Instructions|13479,13498|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|Discharge Instructions|13479,13498|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|Discharge Instructions|13492,13498|false|false|false|C0225386|Breath|breath
Event|Event|Discharge Instructions|13510,13519|false|false|false|||diagnosed
Event|Event|Discharge Instructions|13528,13540|false|false|false|||exacerbation
Finding|Finding|Discharge Instructions|13528,13540|false|false|false|C4086268|Exacerbation|exacerbation
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|13549,13554|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|13549,13554|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Discharge Instructions|13549,13554|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|Discharge Instructions|13549,13562|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Event|Event|Discharge Instructions|13555,13562|false|false|false|||failure
Finding|Functional Concept|Discharge Instructions|13555,13562|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|Discharge Instructions|13555,13562|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|Discharge Instructions|13555,13562|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|Discharge Instructions|13567,13573|false|false|false|||result
Finding|Finding|Discharge Instructions|13567,13573|false|false|false|C1274040;C1546471;C2825142|Experimental Result;Result;What subject filter - Result|result
Finding|Functional Concept|Discharge Instructions|13567,13573|false|false|false|C1274040;C1546471;C2825142|Experimental Result;Result;What subject filter - Result|result
Finding|Idea or Concept|Discharge Instructions|13567,13573|false|false|false|C1274040;C1546471;C2825142|Experimental Result;Result;What subject filter - Result|result
Event|Event|Discharge Instructions|13577,13586|false|false|false|||retaining
Finding|Finding|Discharge Instructions|13587,13595|false|false|false|C3843660|Too much|too much
Finding|Finding|Discharge Instructions|13591,13595|false|false|false|C4281574|Much|much
Drug|Substance|Discharge Instructions|13596,13601|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|Discharge Instructions|13596,13601|false|false|false|||fluid
Finding|Intellectual Product|Discharge Instructions|13596,13601|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|Discharge Instructions|13612,13619|false|false|false|||treated
Drug|Pharmacologic Substance|Discharge Instructions|13626,13635|false|false|false|C0012798|Diuretics|diuretics
Event|Event|Discharge Instructions|13626,13635|false|false|false|||diuretics
Event|Activity|Discharge Instructions|13640,13647|false|false|false|C1883720|Removing (action)|removal
Event|Event|Discharge Instructions|13640,13647|false|false|false|||removal
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|13640,13647|false|false|false|C0015252;C0185115;C0728940|Excision;Extraction;removal technique|removal
Drug|Substance|Discharge Instructions|13656,13661|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|Discharge Instructions|13656,13661|false|false|false|||fluid
Finding|Intellectual Product|Discharge Instructions|13656,13661|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|Discharge Instructions|13678,13689|false|false|false|||improvement
Finding|Conceptual Entity|Discharge Instructions|13678,13689|false|false|false|C2986411|Improvement|improvement
Event|Event|Discharge Instructions|13699,13707|false|false|false|||symptoms
Finding|Functional Concept|Discharge Instructions|13699,13707|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Discharge Instructions|13699,13707|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|Discharge Instructions|13717,13726|false|false|false|||increased
Drug|Organic Chemical|Discharge Instructions|13732,13742|false|false|false|C0054836|carvedilol|carvedilol
Drug|Pharmacologic Substance|Discharge Instructions|13732,13742|false|false|false|C0054836|carvedilol|carvedilol
Event|Event|Discharge Instructions|13743,13747|false|false|false|||dose
Finding|Idea or Concept|Discharge Instructions|13753,13759|false|false|false|C1550462|Observation Interpretation - better|better
Disorder|Disease or Syndrome|Discharge Instructions|13760,13765|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Discharge Instructions|13760,13765|false|false|false|||blood
Finding|Body Substance|Discharge Instructions|13760,13765|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|Discharge Instructions|13760,13774|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Finding|Organism Function|Discharge Instructions|13760,13774|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Procedure|Health Care Activity|Discharge Instructions|13760,13774|false|false|false|C0005824|Blood pressure determination|blood pressure
Event|Event|Discharge Instructions|13766,13774|false|false|false|||pressure
Finding|Finding|Discharge Instructions|13766,13774|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|Discharge Instructions|13766,13774|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|Discharge Instructions|13766,13774|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|Discharge Instructions|13766,13774|false|false|false|C0033095||pressure
Drug|Organic Chemical|Discharge Instructions|13775,13782|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|Discharge Instructions|13775,13782|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|Discharge Instructions|13775,13782|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Event|Event|Discharge Instructions|13775,13782|false|false|false|||control
Finding|Conceptual Entity|Discharge Instructions|13775,13782|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|Discharge Instructions|13775,13782|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|Discharge Instructions|13775,13782|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Finding|Discharge Instructions|13791,13805|false|false|false|C3844729|Very Important|very important
Event|Event|Discharge Instructions|13796,13805|false|false|false|||important
Event|Event|Discharge Instructions|13845,13849|false|false|false|||call
Finding|Functional Concept|Discharge Instructions|13845,13849|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Gene or Genome|Discharge Instructions|13845,13849|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Intellectual Product|Discharge Instructions|13845,13849|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Mental Process|Discharge Instructions|13845,13849|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Attribute|Clinical Attribute|Discharge Instructions|13857,13863|false|false|false|C0944911||weight
Event|Event|Discharge Instructions|13857,13863|false|false|false|||weight
Finding|Finding|Discharge Instructions|13857,13863|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|Discharge Instructions|13857,13863|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|Discharge Instructions|13857,13863|false|false|false|C1305866|Weighing patient|weight
Event|Event|Discharge Instructions|13864,13868|false|false|false|||goes
Procedure|Laboratory Procedure|Discharge Instructions|13884,13887|false|false|false|C3161851|liquid-based cytology (procedure)|lbs
Event|Event|Discharge Instructions|13889,13895|false|false|false|||Taking
Drug|Organic Chemical|Discharge Instructions|13901,13911|false|false|false|C0016860|furosemide|furosemide
Drug|Pharmacologic Substance|Discharge Instructions|13901,13911|false|false|false|C0016860|furosemide|furosemide
Event|Event|Discharge Instructions|13901,13911|false|false|false|||furosemide
Event|Event|Discharge Instructions|13918,13922|false|false|false|||keep
Drug|Substance|Discharge Instructions|13942,13947|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|Discharge Instructions|13942,13947|false|false|false|||fluid
Finding|Intellectual Product|Discharge Instructions|13942,13947|false|false|false|C1546638|Fluid Specimen Code|fluid
Procedure|Health Care Activity|Discharge Instructions|13977,13985|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|13986,13998|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|13986,13998|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|13986,13998|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

