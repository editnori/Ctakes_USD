 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|22,26
No|27,29
:|29,30
_|33,34
_|34,35
_|35,36
<EOL>|36,37
<EOL>|38,39
Admission|39,48
Date|49,53
:|53,54
_|56,57
_|57,58
_|58,59
Discharge|73,82
Date|83,87
:|87,88
_|91,92
_|92,93
_|93,94
<EOL>|94,95
<EOL>|96,97
Date|97,101
of|102,104
Birth|105,110
:|110,111
_|113,114
_|114,115
_|115,116
Sex|129,132
:|132,133
F|136,137
<EOL>|137,138
<EOL>|139,140
Service|140,147
:|147,148
MEDICINE|149,157
<EOL>|157,158
<EOL>|159,160
No|172,174
Known|175,180
Allergies|181,190
/|191,192
Adverse|193,200
Drug|201,205
Reactions|206,215
<EOL>|215,216
<EOL>|217,218
Attending|218,227
:|227,228
_|229,230
_|230,231
_|231,232
.|232,233
<EOL>|233,234
<EOL>|235,236
dyspnea|253,260
<EOL>|260,261
<EOL>|262,263
Major|263,268
Surgical|269,277
or|278,280
Invasive|281,289
Procedure|290,299
:|299,300
<EOL>|300,301
Cardiac|301,308
catheterization|309,324
_|325,326
_|326,327
_|327,328
<EOL>|328,329
<EOL>|329,330
<EOL>|331,332
This|360,364
is|365,367
a|368,369
_|370,371
_|371,372
_|372,373
M|374,375
with|376,380
history|381,388
of|389,391
diabetes|392,400
,|400,401
diastolic|402,411
CHF|412,415
,|415,416
<EOL>|417,418
hypertension|418,430
,|430,431
?|432,433
CAD|433,436
,|436,437
peripheral|438,448
vascular|449,457
disease|458,465
,|465,466
CKD|467,470
presenting|471,481
<EOL>|482,483
with|483,487
_|488,489
_|489,490
_|490,491
days|492,496
of|497,499
increasing|500,510
dyspnea|511,518
and|519,522
non-productive|523,537
cough|538,543
.|543,544
<EOL>|545,546
She|546,549
denies|550,556
fevers|557,563
,|563,564
chills|565,571
,|571,572
chest|573,578
pain|579,583
,|583,584
nausea|585,591
,|591,592
vomiting|593,601
.|601,602
Did|603,606
<EOL>|607,608
report|608,614
feeling|615,622
somewhat|623,631
wheezy|632,638
.|638,639
Denies|640,646
leg|647,650
swelling|651,659
,|659,660
has|661,664
<EOL>|665,666
possibly|666,674
had|675,678
a|679,680
2|681,682
lb|683,685
weight|686,692
gain|693,697
.|697,698
Denies|699,705
missed|706,712
medication|713,723
doses|724,729
.|729,730
<EOL>|731,732
Does|732,736
report|737,743
2|744,745
pillow|746,752
orthopnea|753,762
last|763,767
night|768,773
.|773,774
Her|775,778
husband|779,786
has|787,790
also|791,795
<EOL>|796,797
been|797,801
sick|802,806
with|807,811
a|812,813
cough|814,819
for|820,823
the|824,827
past|828,832
day|833,836
or|837,839
so|840,842
.|842,843
She|844,847
is|848,850
a|851,852
<EOL>|853,854
non-smoker|854,864
.|864,865
She|866,869
lives|870,875
at|876,878
home|879,883
and|884,887
has|888,891
had|892,895
no|896,898
recent|899,905
<EOL>|906,907
hospitalizations|907,923
or|924,926
courses|927,934
of|935,937
antibiotics|938,949
.|949,950
<EOL>|950,951
<EOL>|951,952
In|952,954
the|955,958
ED|959,961
,|961,962
initial|963,970
vitals|971,977
:|977,978
97.8|980,984
80|985,987
132|988,991
/|991,992
83|992,994
25|995,997
97|998,1000
%|1000,1001
ra|1002,1004
.|1004,1005
CXR|1006,1009
showed|1010,1016
<EOL>|1017,1018
probable|1018,1026
RUL|1027,1030
PNA|1031,1034
.|1034,1035
Normal|1036,1042
WBC|1043,1046
and|1047,1050
lactate|1051,1058
,|1058,1059
Cr|1060,1062
at|1063,1065
baseline|1066,1074
.|1074,1075
<EOL>|1077,1078
Troponin|1078,1086
0.09|1087,1091
with|1092,1096
normal|1097,1103
CK|1104,1106
-|1106,1107
MB|1107,1109
.|1109,1110
BNP|1111,1114
2826|1115,1119
.|1119,1120
She|1121,1124
was|1125,1128
started|1129,1136
on|1137,1139
<EOL>|1140,1141
bipap|1141,1146
due|1147,1150
to|1151,1153
tachypnea|1154,1163
and|1164,1167
increased|1168,1177
work|1178,1182
of|1183,1185
breathing|1186,1195
.|1195,1196
She|1197,1200
was|1201,1204
<EOL>|1205,1206
given|1206,1211
40mg|1212,1216
IV|1217,1219
lasix|1220,1225
and|1226,1229
started|1230,1237
on|1238,1240
vancomycin|1241,1251
,|1251,1252
cefepime|1253,1261
and|1262,1265
<EOL>|1266,1267
levofloxacin|1267,1279
.|1279,1280
<EOL>|1280,1281
<EOL>|1282,1283
On|1283,1285
transfer|1286,1294
,|1294,1295
vitals|1296,1302
were|1303,1307
:|1307,1308
69|1310,1312
141|1313,1316
/|1316,1317
82|1317,1319
28|1320,1322
100|1323,1326
%|1326,1327
bipap|1328,1333
<EOL>|1334,1335
<EOL>|1335,1336
On|1336,1338
arrival|1339,1346
to|1347,1349
the|1350,1353
MICU|1354,1358
,|1358,1359
patient|1360,1367
reports|1368,1375
improved|1376,1384
breathing|1385,1394
on|1395,1397
<EOL>|1398,1399
bipap|1399,1404
.|1404,1405
<EOL>|1407,1408
<EOL>|1408,1409
Review|1409,1415
of|1416,1418
systems|1419,1426
:|1426,1427
<EOL>|1429,1430
(|1430,1431
+|1431,1432
)|1432,1433
Per|1434,1437
HPI|1438,1441
<EOL>|1443,1444
<EOL>|1445,1446
-|1468,1469
hypertension|1470,1482
<EOL>|1482,1483
-|1483,1484
diabetes|1485,1493
<EOL>|1493,1494
-|1494,1495
hx|1496,1498
CVA|1499,1502
(|1503,1504
cerebellar|1504,1514
-|1514,1515
medullary|1515,1524
stroke|1525,1531
in|1532,1534
_|1535,1536
_|1536,1537
_|1537,1538
<EOL>|1538,1539
-|1539,1540
CAD|1541,1544
(|1545,1546
has|1546,1549
never|1550,1555
been|1556,1560
cathed|1561,1567
,|1567,1568
hx|1569,1571
of|1572,1574
MI|1575,1577
in|1578,1580
_|1581,1582
_|1582,1583
_|1583,1584
<EOL>|1584,1585
-|1585,1586
peripheral|1587,1597
arterial|1598,1606
disease|1607,1614
-|1614,1615
claudication|1616,1628
,|1628,1629
followed|1630,1638
by|1639,1641
<EOL>|1642,1643
vascular|1643,1651
,|1651,1652
managed|1653,1660
conservatively|1661,1675
<EOL>|1675,1676
-|1676,1677
stage|1678,1683
IV|1684,1686
CKD|1687,1690
(|1691,1692
baseline|1692,1700
2.5|1701,1704
-|1704,1705
2.8|1705,1708
)|1708,1709
<EOL>|1709,1710
-|1710,1711
GERD|1712,1716
/|1716,1717
esophageal|1717,1727
rings|1728,1733
<EOL>|1733,1734
<EOL>|1735,1736
:|1750,1751
<EOL>|1751,1752
_|1752,1753
_|1753,1754
_|1754,1755
<EOL>|1755,1756
:|1770,1771
<EOL>|1771,1772
Niece|1772,1777
had|1778,1781
some|1782,1786
sort|1787,1791
of|1792,1794
cancer|1795,1801
.|1801,1802
Otherwise|1803,1812
,|1812,1813
no|1814,1816
family|1817,1823
history|1824,1831
of|1832,1834
<EOL>|1835,1836
cancer|1836,1842
or|1843,1845
early|1846,1851
heart|1852,1857
disease|1858,1865
.|1865,1866
<EOL>|1866,1867
<EOL>|1868,1869
ADMISSION|1884,1893
EXAM|1894,1898
:|1898,1899
<EOL>|1899,1900
General|1900,1907
-|1907,1908
appears|1910,1917
comfortable|1918,1929
on|1930,1932
BiPap|1933,1938
<EOL>|1938,1939
HEENT|1939,1944
-|1944,1945
PERRL|1946,1951
,|1951,1952
EOMI|1953,1957
<EOL>|1958,1959
Neck|1959,1963
-|1963,1964
difficult|1965,1974
to|1975,1977
assess|1978,1984
JVP|1985,1988
due|1989,1992
to|1993,1995
habitus|1996,2003
and|2004,2007
presence|2008,2016
of|2017,2019
<EOL>|2020,2021
BiPap|2021,2026
strap|2027,2032
<EOL>|2033,2034
CV|2034,2036
-|2036,2037
RRR|2039,2042
,|2042,2043
no|2044,2046
gallops|2047,2054
<EOL>|2054,2055
Lungs|2055,2060
-|2060,2061
good|2063,2067
air|2068,2071
entry|2072,2077
.|2077,2078
diffuse|2079,2086
crackles|2087,2095
R|2096,2097
>|2097,2098
L|2098,2099
,|2099,2100
rhonchi|2101,2108
in|2109,2111
RUL|2112,2115
.|2115,2116
<EOL>|2117,2118
scattered|2118,2127
inspiratory|2128,2139
wheezing|2140,2148
<EOL>|2148,2149
Abdomen|2149,2156
-|2156,2157
soft|2159,2163
,|2163,2164
NTND|2165,2169
<EOL>|2169,2170
Ext|2170,2173
-|2173,2174
trace|2176,2181
edema|2182,2187
,|2187,2188
faint|2189,2194
peripheral|2195,2205
pulses|2206,2212
<EOL>|2212,2213
Neuro|2213,2218
-|2218,2219
A|2221,2222
and|2223,2226
O|2227,2228
x|2229,2230
3|2231,2232
,|2232,2233
moving|2234,2240
all|2241,2244
4|2245,2246
extremities|2247,2258
.|2258,2259
mildly|2260,2266
decreased|2267,2276
<EOL>|2277,2278
strength|2278,2286
in|2287,2289
LLL|2290,2293
<EOL>|2293,2294
<EOL>|2294,2295
DISCHARGE|2295,2304
EXAM|2305,2309
:|2309,2310
<EOL>|2310,2311
VS|2311,2313
:|2313,2314
T98|2315,2318
.9|2318,2320
BP144|2321,2326
/|2326,2327
83|2327,2329
P66|2330,2333
RR18|2334,2338
99RA|2339,2343
76|2344,2346
.|2346,2347
1kg|2347,2350
<EOL>|2350,2351
GENERAL|2351,2358
:|2358,2359
Laying|2360,2366
in|2367,2369
bed|2370,2373
,|2373,2374
sleeping|2375,2383
.|2383,2384
No|2385,2387
acute|2388,2393
distress|2394,2402
.|2402,2403
<EOL>|2405,2406
HEENT|2406,2411
:|2411,2412
Moist|2413,2418
mucous|2419,2425
membranes|2426,2435
.|2435,2436
<EOL>|2437,2438
NECK|2438,2442
:|2442,2443
Supple|2444,2450
,|2450,2451
unable|2452,2458
to|2459,2461
visualize|2462,2471
JVP|2472,2475
.|2475,2476
<EOL>|2476,2477
CARDIAC|2477,2484
:|2484,2485
Regular|2486,2493
rate|2494,2498
and|2499,2502
rhythm|2503,2509
.|2509,2510
Normal|2511,2517
S1|2518,2520
,|2520,2521
S2|2522,2524
.|2524,2525
No|2526,2528
S3|2529,2531
,|2531,2532
S4|2533,2535
.|2535,2536
_|2537,2538
_|2538,2539
_|2539,2540
<EOL>|2541,2542
systolic|2542,2550
murmur|2551,2557
.|2557,2558
<EOL>|2558,2559
LUNGS|2559,2564
:|2564,2565
Clear|2566,2571
to|2572,2574
auscultation|2575,2587
bilaterally|2588,2599
.|2599,2600
No|2601,2603
crackles|2604,2612
,|2612,2613
wheezes|2614,2621
,|2621,2622
<EOL>|2623,2624
rhonchi|2624,2631
.|2631,2632
<EOL>|2634,2635
ABDOMEN|2635,2642
:|2642,2643
+|2644,2645
BS|2645,2647
,|2647,2648
soft|2649,2653
,|2653,2654
nondistended|2655,2667
,|2667,2668
nontender|2669,2678
to|2679,2681
palpation|2682,2691
.|2691,2692
<EOL>|2695,2696
EXTREMITIES|2696,2707
:|2707,2708
Warm|2709,2713
and|2714,2717
well|2718,2722
perfused|2723,2731
.|2731,2732
Pulses|2733,2739
2|2740,2741
+|2741,2742
.|2742,2743
Trace|2744,2749
peripheral|2750,2760
<EOL>|2761,2762
edema|2762,2767
.|2767,2768
<EOL>|2769,2770
<EOL>|2771,2772
Pertinent|2772,2781
Results|2782,2789
:|2789,2790
<EOL>|2790,2791
ON|2791,2793
ADMISSION|2794,2803
:|2803,2804
<EOL>|2804,2805
<EOL>|2805,2806
_|2806,2807
_|2807,2808
_|2808,2809
06|2810,2812
:|2812,2813
48AM|2813,2817
BLOOD|2818,2823
WBC|2824,2827
-|2827,2828
5.3|2828,2831
RBC|2832,2835
-|2835,2836
2|2836,2837
.|2837,2838
94|2838,2840
*|2840,2841
Hgb|2842,2845
-|2845,2846
9|2846,2847
.|2847,2848
5|2848,2849
*|2849,2850
Hct|2851,2854
-|2854,2855
27|2855,2857
.|2857,2858
3|2858,2859
*|2859,2860
<EOL>|2861,2862
MCV|2862,2865
-|2865,2866
93|2866,2868
MCH|2869,2872
-|2872,2873
32|2873,2875
.|2875,2876
4|2876,2877
*|2877,2878
MCHC|2879,2883
-|2883,2884
34.9|2884,2888
RDW|2889,2892
-|2892,2893
13.5|2893,2897
Plt|2898,2901
_|2902,2903
_|2903,2904
_|2904,2905
<EOL>|2905,2906
_|2906,2907
_|2907,2908
_|2908,2909
06|2910,2912
:|2912,2913
48AM|2913,2917
BLOOD|2918,2923
Neuts|2924,2929
-|2929,2930
65.6|2930,2934
_|2935,2936
_|2936,2937
_|2937,2938
Monos|2939,2944
-|2944,2945
5.2|2945,2948
Eos|2949,2952
-|2952,2953
2.7|2953,2956
<EOL>|2957,2958
Baso|2958,2962
-|2962,2963
0.4|2963,2966
<EOL>|2966,2967
_|2967,2968
_|2968,2969
_|2969,2970
08|2971,2973
:|2973,2974
03PM|2974,2978
BLOOD|2979,2984
_|2985,2986
_|2986,2987
_|2987,2988
PTT|2989,2992
-|2992,2993
69|2993,2995
.|2995,2996
6|2996,2997
*|2997,2998
_|2999,3000
_|3000,3001
_|3001,3002
<EOL>|3002,3003
_|3003,3004
_|3004,3005
_|3005,3006
06|3007,3009
:|3009,3010
48AM|3010,3014
BLOOD|3015,3020
Glucose|3021,3028
-|3028,3029
89|3029,3031
UreaN|3032,3037
-|3037,3038
37|3038,3040
*|3040,3041
Creat|3042,3047
-|3047,3048
2|3048,3049
.|3049,3050
3|3050,3051
*|3051,3052
Na|3053,3055
-|3055,3056
144|3056,3059
<EOL>|3060,3061
K|3061,3062
-|3062,3063
3.9|3063,3066
Cl|3067,3069
-|3069,3070
109|3070,3073
*|3073,3074
HCO3|3075,3079
-|3079,3080
21|3080,3082
*|3082,3083
AnGap|3084,3089
-|3089,3090
18|3090,3092
<EOL>|3092,3093
_|3093,3094
_|3094,3095
_|3095,3096
06|3097,3099
:|3099,3100
48AM|3100,3104
BLOOD|3105,3110
CK|3111,3113
-|3113,3114
MB|3114,3116
-|3116,3117
6|3117,3118
proBNP|3119,3125
-|3125,3126
2826|3126,3130
*|3130,3131
<EOL>|3131,3132
_|3132,3133
_|3133,3134
_|3134,3135
06|3136,3138
:|3138,3139
48AM|3139,3143
BLOOD|3144,3149
cTropnT|3150,3157
-|3157,3158
0|3158,3159
.|3159,3160
09|3160,3162
*|3162,3163
<EOL>|3163,3164
_|3164,3165
_|3165,3166
_|3166,3167
12|3168,3170
:|3170,3171
58PM|3171,3175
BLOOD|3176,3181
CK|3182,3184
-|3184,3185
MB|3185,3187
-|3187,3188
9|3188,3189
cTropnT|3190,3197
-|3197,3198
0|3198,3199
.|3199,3200
11|3200,3202
*|3202,3203
<EOL>|3203,3204
_|3204,3205
_|3205,3206
_|3206,3207
07|3208,3210
:|3210,3211
52AM|3211,3215
BLOOD|3216,3221
Lactate|3222,3229
-|3229,3230
1.7|3230,3233
<EOL>|3233,3234
_|3234,3235
_|3235,3236
_|3236,3237
07|3238,3240
:|3240,3241
40AM|3241,3245
URINE|3246,3251
Color|3252,3257
-|3257,3258
Straw|3258,3263
Appear|3264,3270
-|3270,3271
Clear|3271,3276
Sp|3277,3279
_|3280,3281
_|3281,3282
_|3282,3283
<EOL>|3283,3284
_|3284,3285
_|3285,3286
_|3286,3287
07|3288,3290
:|3290,3291
40AM|3291,3295
URINE|3296,3301
Blood|3302,3307
-|3307,3308
NEG|3308,3311
Nitrite|3312,3319
-|3319,3320
NEG|3320,3323
Protein|3324,3331
-|3331,3332
NEG|3332,3335
<EOL>|3336,3337
Glucose|3337,3344
-|3344,3345
NEG|3345,3348
Ketone|3349,3355
-|3355,3356
NEG|3356,3359
Bilirub|3360,3367
-|3367,3368
NEG|3368,3371
Urobiln|3372,3379
-|3379,3380
NEG|3380,3383
pH|3384,3386
-|3386,3387
6.0|3387,3390
Leuks|3391,3396
-|3396,3397
NEG|3397,3400
<EOL>|3400,3401
<EOL>|3401,3402
ON|3402,3404
DISCHARGE|3405,3414
:|3414,3415
<EOL>|3415,3416
<EOL>|3416,3417
_|3417,3418
_|3418,3419
_|3419,3420
09|3421,3423
:|3423,3424
00AM|3424,3428
BLOOD|3429,3434
WBC|3435,3438
-|3438,3439
4.8|3439,3442
RBC|3443,3446
-|3446,3447
2|3447,3448
.|3448,3449
53|3449,3451
*|3451,3452
Hgb|3453,3456
-|3456,3457
8|3457,3458
.|3458,3459
0|3459,3460
*|3460,3461
Hct|3462,3465
-|3465,3466
23|3466,3468
.|3468,3469
6|3469,3470
*|3470,3471
<EOL>|3472,3473
MCV|3473,3476
-|3476,3477
94|3477,3479
MCH|3480,3483
-|3483,3484
31.5|3484,3488
MCHC|3489,3493
-|3493,3494
33.7|3494,3498
RDW|3499,3502
-|3502,3503
12.9|3503,3507
Plt|3508,3511
_|3512,3513
_|3513,3514
_|3514,3515
<EOL>|3515,3516
_|3516,3517
_|3517,3518
_|3518,3519
09|3520,3522
:|3522,3523
26AM|3523,3527
BLOOD|3528,3533
Glucose|3534,3541
-|3541,3542
121|3542,3545
*|3545,3546
UreaN|3547,3552
-|3552,3553
52|3553,3555
*|3555,3556
Creat|3557,3562
-|3562,3563
2|3563,3564
.|3564,3565
2|3565,3566
*|3566,3567
Na|3568,3570
-|3570,3571
142|3571,3574
<EOL>|3575,3576
K|3576,3577
-|3577,3578
4.5|3578,3581
Cl|3582,3584
-|3584,3585
108|3585,3588
HCO3|3589,3593
-|3593,3594
24|3594,3596
AnGap|3597,3602
-|3602,3603
15|3603,3605
<EOL>|3605,3606
_|3606,3607
_|3607,3608
_|3608,3609
09|3610,3612
:|3612,3613
26AM|3613,3617
BLOOD|3618,3623
Calcium|3624,3631
-|3631,3632
9.9|3632,3635
Phos|3636,3640
-|3640,3641
4|3641,3642
.|3642,3643
8|3643,3644
*|3644,3645
Mg|3646,3648
-|3648,3649
2.5|3649,3652
<EOL>|3652,3653
<EOL>|3653,3654
CXR|3654,3657
:|3657,3658
_|3659,3660
_|3660,3661
_|3661,3662
<EOL>|3662,3663
Right|3663,3668
upper|3669,3674
lobe|3675,3679
pneumonia|3680,3689
or|3690,3692
mass|3693,3697
.|3697,3698
However|3700,3707
,|3707,3708
given|3709,3714
right|3715,3720
hilar|3721,3726
<EOL>|3727,3728
fullness|3728,3736
,|3736,3737
a|3738,3739
mass|3740,3744
resulting|3745,3754
in|3755,3757
post-obstructive|3758,3774
pneumonia|3775,3784
is|3785,3787
<EOL>|3788,3789
within|3789,3795
the|3796,3799
<EOL>|3800,3801
differential|3801,3813
.|3813,3814
Recommend|3816,3825
chest|3826,3831
CT|3832,3834
with|3835,3839
intravenous|3840,3851
contrast|3852,3860
for|3861,3864
<EOL>|3865,3866
further|3866,3873
<EOL>|3874,3875
assessment|3875,3885
.|3885,3886
<EOL>|3887,3888
<EOL>|3888,3889
TTE|3889,3892
:|3892,3893
_|3894,3895
_|3895,3896
_|3896,3897
<EOL>|3897,3898
The|3898,3901
left|3902,3906
atrium|3907,3913
is|3914,3916
elongated|3917,3926
.|3926,3927
There|3928,3933
is|3934,3936
mild|3937,3941
symmetric|3942,3951
left|3952,3956
<EOL>|3957,3958
ventricular|3958,3969
hypertrophy|3970,3981
with|3982,3986
normal|3987,3993
cavity|3994,4000
size|4001,4005
.|4005,4006
There|4007,4012
is|4013,4015
mild|4016,4020
<EOL>|4021,4022
to|4022,4024
moderate|4025,4033
regional|4034,4042
left|4043,4047
ventricular|4048,4059
systolic|4060,4068
dysfunction|4069,4080
with|4081,4085
<EOL>|4086,4087
near|4087,4091
-|4091,4092
akinesis|4092,4100
of|4101,4103
the|4104,4107
inferior|4108,4116
,|4116,4117
inferolateral|4118,4131
and|4132,4135
basal|4136,4141
lateral|4142,4149
<EOL>|4150,4151
segments|4151,4159
.|4159,4160
The|4161,4164
remaining|4165,4174
segments|4175,4183
contract|4184,4192
normally|4193,4201
(|4202,4203
LVEF|4203,4207
=|4208,4209
<EOL>|4210,4211
35|4211,4213
-|4213,4214
40|4214,4216
%|4216,4217
)|4217,4218
.|4218,4219
Right|4220,4225
ventricular|4226,4237
chamber|4238,4245
size|4246,4250
and|4251,4254
free|4255,4259
wall|4260,4264
motion|4265,4271
are|4272,4275
<EOL>|4276,4277
normal|4277,4283
.|4283,4284
The|4285,4288
aortic|4289,4295
valve|4296,4301
leaflets|4302,4310
(|4311,4312
3|4312,4313
)|4313,4314
are|4315,4318
mildly|4319,4325
thickened|4326,4335
but|4336,4339
<EOL>|4340,4341
aortic|4341,4347
stenosis|4348,4356
is|4357,4359
not|4360,4363
present|4364,4371
.|4371,4372
No|4373,4375
aortic|4376,4382
regurgitation|4383,4396
is|4397,4399
seen|4400,4404
.|4404,4405
<EOL>|4406,4407
The|4407,4410
mitral|4411,4417
valve|4418,4423
leaflets|4424,4432
are|4433,4436
mildly|4437,4443
thickened|4444,4453
.|4453,4454
An|4455,4457
eccentric|4458,4467
jet|4468,4471
<EOL>|4472,4473
of|4473,4475
moderate|4476,4484
to|4485,4487
severe|4488,4494
(|4495,4496
3|4496,4497
+|4497,4498
)|4498,4499
mitral|4500,4506
regurgitation|4507,4520
is|4521,4523
seen|4524,4528
.|4528,4529
There|4530,4535
<EOL>|4536,4537
is|4537,4539
moderate|4540,4548
pulmonary|4549,4558
artery|4559,4565
systolic|4566,4574
hypertension|4575,4587
.|4587,4588
There|4589,4594
is|4595,4597
no|4598,4600
<EOL>|4601,4602
pericardial|4602,4613
effusion|4614,4622
.|4622,4623
<EOL>|4623,4624
<EOL>|4624,4625
IMPRESSION|4625,4635
:|4635,4636
Mild|4637,4641
to|4642,4644
moderate|4645,4653
regional|4654,4662
left|4663,4667
ventricular|4668,4679
systolic|4680,4688
<EOL>|4689,4690
dysfunction|4690,4701
,|4701,4702
c|4703,4704
/|4704,4705
w|4705,4706
CAD|4707,4710
.|4710,4711
Moderate|4712,4720
to|4721,4723
severe|4724,4730
mitral|4731,4737
regurgitation|4738,4751
.|4751,4752
<EOL>|4753,4754
Moderate|4754,4762
pulmonary|4763,4772
hypertension|4773,4785
.|4785,4786
<EOL>|4786,4787
<EOL>|4787,4788
Compared|4788,4796
with|4797,4801
the|4802,4805
prior|4806,4811
study|4812,4817
(|4818,4819
images|4819,4825
reviewed|4826,4834
)|4834,4835
of|4836,4838
_|4839,4840
_|4840,4841
_|4841,4842
,|4842,4843
<EOL>|4844,4845
regional|4845,4853
LV|4854,4856
wall|4857,4861
motion|4862,4868
abnormalities|4869,4882
are|4883,4886
new|4887,4890
.|4890,4891
Severity|4892,4900
of|4901,4903
<EOL>|4904,4905
mitral|4905,4911
regurgitation|4912,4925
has|4926,4929
increased|4930,4939
.|4939,4940
<EOL>|4940,4941
<EOL>|4941,4942
CARDIAC|4942,4949
CATH|4950,4954
:|4954,4955
_|4956,4957
_|4957,4958
_|4958,4959
<EOL>|4959,4960
1.|4960,4962
Selective|4963,4972
coronary|4973,4981
angiography|4982,4993
of|4994,4996
this|4997,5001
right|5002,5007
dominant|5008,5016
system|5017,5023
<EOL>|5024,5025
revealed|5025,5033
three|5034,5039
vessel|5040,5046
coronary|5047,5055
artery|5056,5062
disease|5063,5070
.|5070,5071
The|5073,5076
LMCA|5077,5081
had|5082,5085
no|5086,5088
<EOL>|5089,5090
obstructive|5090,5101
disease|5102,5109
.|5109,5110
The|5112,5115
LAD|5116,5119
had|5120,5123
a|5124,5125
moderate|5126,5134
disease|5135,5142
in|5143,5145
the|5146,5149
mid|5150,5153
<EOL>|5154,5155
artery|5155,5161
and|5162,5165
a|5166,5167
diagonal|5168,5176
branch|5177,5183
had|5184,5187
an|5188,5190
80|5191,5193
%|5193,5194
proximal|5195,5203
lesion|5204,5210
.|5210,5211
The|5213,5216
<EOL>|5217,5218
Lcx|5218,5221
had|5222,5225
a|5226,5227
70|5228,5230
%|5230,5231
proximal|5232,5240
lesion|5241,5247
.|5247,5248
The|5250,5253
RCA|5254,5257
was|5258,5261
totally|5262,5269
occluded|5270,5278
<EOL>|5279,5280
mid-vessel|5280,5290
.|5290,5291
<EOL>|5292,5293
<EOL>|5295,5296
1.|5318,5320
Three|5321,5326
vessel|5327,5333
coronary|5334,5342
artery|5343,5349
disease|5350,5357
.|5357,5358
<EOL>|5359,5360
2.|5360,5362
Recommend|5363,5372
CABG|5373,5377
evaluation|5378,5388
<EOL>|5388,5389
<EOL>|5389,5390
CT|5390,5392
CHEST|5393,5398
:|5398,5399
_|5400,5401
_|5401,5402
_|5402,5403
<EOL>|5403,5404
1.|5404,5406
Diffuse|5408,5415
confluent|5416,5425
ground|5426,5432
-|5432,5433
glass|5433,5438
opacities|5439,5448
predominantly|5449,5462
in|5463,5465
<EOL>|5466,5467
the|5467,5470
right|5471,5476
upper|5477,5482
lobe|5483,5487
and|5488,5491
right|5492,5497
lower|5498,5503
lobe|5504,5508
most|5509,5513
likely|5514,5520
represent|5521,5530
<EOL>|5531,5532
residual|5532,5540
pulmonary|5541,5550
edema|5551,5556
,|5556,5557
localized|5558,5567
to|5568,5570
the|5571,5574
right|5575,5580
lung|5581,5585
because|5586,5593
of|5594,5596
<EOL>|5597,5598
direction|5598,5607
of|5608,5610
jet|5611,5614
in|5615,5617
mitral|5618,5624
<EOL>|5625,5626
regurgitation|5626,5639
.|5639,5640
<EOL>|5642,5643
2|5643,5644
.|5644,5645
Possible|5647,5655
pulmonary|5656,5665
hypertension|5666,5678
.|5678,5679
<EOL>|5680,5681
3.|5681,5683
Moderate|5685,5693
coronary|5694,5702
artery|5703,5709
disease|5710,5717
.|5717,5718
<EOL>|5719,5720
<EOL>|5720,5721
CAROTID|5721,5728
US|5729,5731
:|5731,5732
_|5733,5734
_|5734,5735
_|5735,5736
<EOL>|5736,5737
No|5737,5739
evidence|5740,5748
of|5749,5751
hemodynamically|5752,5767
significant|5768,5779
internal|5780,5788
carotid|5789,5796
<EOL>|5797,5798
stenosis|5798,5806
on|5807,5809
either|5810,5816
side|5817,5821
.|5821,5822
<EOL>|5823,5824
<EOL>|5824,5825
ECHO|5825,5829
_|5830,5831
_|5831,5832
_|5832,5833
-|5833,5834
PCI|5835,5838
)|5838,5839
<EOL>|5839,5840
There|5840,5845
is|5846,5848
mild|5849,5853
symmetric|5854,5863
left|5864,5868
ventricular|5869,5880
hypertrophy|5881,5892
with|5893,5897
normal|5898,5904
<EOL>|5905,5906
cavity|5906,5912
size|5913,5917
.|5917,5918
There|5919,5924
is|5925,5927
mild|5928,5932
regional|5933,5941
left|5942,5946
ventricular|5947,5958
systolic|5959,5967
<EOL>|5968,5969
dysfunction|5969,5980
with|5981,5985
inferior|5986,5994
and|5995,5998
infero|5999,6005
-|6005,6006
lateral|6006,6013
hypokinesis|6014,6025
.|6025,6026
No|6027,6029
<EOL>|6030,6031
masses|6031,6037
or|6038,6040
thrombi|6041,6048
are|6049,6052
seen|6053,6057
in|6058,6060
the|6061,6064
left|6065,6069
ventricle|6070,6079
.|6079,6080
There|6081,6086
is|6087,6089
no|6090,6092
<EOL>|6093,6094
ventricular|6094,6105
septal|6106,6112
defect|6113,6119
.|6119,6120
Right|6121,6126
ventricular|6127,6138
chamber|6139,6146
size|6147,6151
and|6152,6155
<EOL>|6156,6157
free|6157,6161
wall|6162,6166
motion|6167,6173
are|6174,6177
normal|6178,6184
.|6184,6185
The|6186,6189
mitral|6190,6196
valve|6197,6202
leaflets|6203,6211
are|6212,6215
<EOL>|6216,6217
mildly|6217,6223
thickened|6224,6233
.|6233,6234
An|6235,6237
eccentric|6238,6247
jet|6248,6251
of|6252,6254
mild|6255,6259
(|6260,6261
1|6261,6262
+|6262,6263
)|6263,6264
mitral|6265,6271
<EOL>|6272,6273
regurgitation|6273,6286
is|6287,6289
seen|6290,6294
.|6294,6295
There|6296,6301
is|6302,6304
no|6305,6307
pericardial|6308,6319
effusion|6320,6328
.|6328,6329
<EOL>|6330,6331
<EOL>|6331,6332
Compared|6332,6340
with|6341,6345
the|6346,6349
prior|6350,6355
study|6356,6361
(|6362,6363
images|6363,6369
reviewed|6370,6378
)|6378,6379
of|6380,6382
_|6383,6384
_|6384,6385
_|6385,6386
,|6386,6387
<EOL>|6388,6389
the|6389,6392
LVEF|6393,6397
has|6398,6401
increased|6402,6411
.|6411,6412
The|6413,6416
degree|6417,6423
of|6424,6426
MR|6427,6429
seen|6430,6434
has|6435,6438
decreased|6439,6448
.|6448,6449
<EOL>|6450,6451
<EOL>|6451,6452
<EOL>|6453,6454
_|6477,6478
_|6478,6479
_|6479,6480
female|6481,6487
with|6488,6492
_|6493,6494
_|6494,6495
_|6495,6496
,|6496,6497
HTN|6498,6501
,|6501,6502
diabetes|6503,6511
,|6511,6512
CKD|6513,6516
presented|6517,6526
with|6527,6531
<EOL>|6532,6533
increased|6533,6542
dyspnea|6543,6550
and|6551,6554
non-productive|6555,6569
cough|6570,6575
without|6576,6583
fevers|6584,6590
or|6591,6593
<EOL>|6594,6595
elevated|6595,6603
white|6604,6609
count|6610,6615
,|6615,6616
initially|6617,6626
admitted|6627,6635
to|6636,6638
_|6639,6640
_|6640,6641
_|6641,6642
with|6643,6647
concern|6648,6655
<EOL>|6656,6657
for|6657,6660
pneumonia|6661,6670
.|6670,6671
However|6672,6679
,|6679,6680
was|6681,6684
found|6685,6690
to|6691,6693
have|6694,6698
ST|6699,6701
-|6701,6702
changes|6702,6709
,|6709,6710
enzyme|6711,6717
<EOL>|6718,6719
leak|6719,6723
,|6723,6724
new|6725,6728
wall|6729,6733
motion|6734,6740
abnormality|6741,6752
consistent|6753,6763
with|6764,6768
a|6769,6770
recent|6771,6777
<EOL>|6778,6779
cardiac|6779,6786
event|6787,6792
and|6793,6796
had|6797,6800
no|6801,6803
evidence|6804,6812
of|6813,6815
pneumonia|6816,6825
(|6826,6827
no|6827,6829
fevers|6830,6836
,|6836,6837
wbc|6838,6841
,|6841,6842
<EOL>|6843,6844
lactate|6844,6851
,|6851,6852
normal|6853,6859
vitals|6860,6866
,|6866,6867
CXR|6868,6871
with|6872,6876
likely|6877,6883
one|6884,6887
sided|6888,6893
pulmonary|6894,6903
<EOL>|6904,6905
edema|6905,6910
from|6911,6915
mitral|6916,6922
regurgitation|6923,6936
)|6936,6937
.|6937,6938
She|6939,6942
was|6943,6946
seen|6947,6951
by|6952,6954
cardiology|6955,6965
who|6966,6969
<EOL>|6970,6971
transferred|6971,6982
the|6983,6986
patient|6987,6994
to|6995,6997
cardiology|6998,7008
floor|7009,7014
.|7014,7015
<EOL>|7015,7016
<EOL>|7016,7017
#|7017,7018
Acute|7019,7024
systolic|7025,7033
CHF|7034,7037
exacerbation|7038,7050
/|7050,7051
mitral|7051,7057
regurgitation|7058,7071
:|7071,7072
<EOL>|7073,7074
Likely|7074,7080
secondary|7081,7090
to|7091,7093
ischemic|7094,7102
valvular|7103,7111
disease|7112,7119
resulting|7120,7129
in|7130,7132
<EOL>|7133,7134
worsening|7134,7143
mitral|7144,7150
regurgitation|7151,7164
.|7164,7165
ECHO|7166,7170
also|7171,7175
with|7176,7180
akinetic|7181,7189
inferior|7190,7198
<EOL>|7199,7200
wall|7200,7204
segments|7205,7213
,|7213,7214
which|7215,7220
also|7221,7225
supports|7226,7234
an|7235,7237
ischemic|7238,7246
event|7247,7252
.|7252,7253
Cardiac|7254,7261
<EOL>|7262,7263
cath|7263,7267
revealed|7268,7276
3|7277,7278
vessel|7279,7285
disease|7286,7293
.|7293,7294
Patient|7295,7302
was|7303,7306
managed|7307,7314
medically|7315,7324
<EOL>|7325,7326
with|7326,7330
lasix|7331,7336
,|7336,7337
lisinopril|7338,7348
,|7348,7349
and|7350,7353
metoprolol|7354,7364
.|7364,7365
Cardiac|7366,7373
surgery|7374,7381
was|7382,7385
<EOL>|7386,7387
consulted|7387,7396
for|7397,7400
possible|7401,7409
CABG|7410,7414
and|7415,7418
mitral|7419,7425
valve|7426,7431
repair|7432,7438
/|7438,7439
replacement|7439,7450
.|7450,7451
<EOL>|7452,7453
However|7453,7460
,|7460,7461
given|7462,7467
her|7468,7471
multiple|7472,7480
comorbidities|7481,7494
,|7494,7495
she|7496,7499
is|7500,7502
extremely|7503,7512
high|7513,7517
<EOL>|7518,7519
risk|7519,7523
and|7524,7527
surgery|7528,7535
was|7536,7539
deferred|7540,7548
.|7548,7549
Therefore|7550,7559
,|7559,7560
the|7561,7564
decision|7565,7573
was|7574,7577
made|7578,7582
<EOL>|7583,7584
to|7584,7586
revascularize|7587,7600
the|7601,7604
patient|7605,7612
with|7613,7617
PCI|7618,7621
to|7622,7624
see|7625,7628
if|7629,7631
the|7632,7635
patient|7636,7643
<EOL>|7644,7645
would|7645,7650
regain|7651,7657
function|7658,7666
of|7667,7669
her|7670,7673
mitral|7674,7680
valve|7681,7686
.|7686,7687
Patient|7688,7695
received|7696,7704
a|7705,7706
<EOL>|7707,7708
bare|7708,7712
metal|7713,7718
stent|7719,7724
in|7725,7727
the|7728,7731
LCx|7732,7735
and|7736,7739
plain|7740,7745
old|7746,7749
balloon|7750,7757
angioplasty|7758,7769
in|7770,7772
<EOL>|7773,7774
the|7774,7777
diagonal|7778,7786
artery|7787,7793
.|7793,7794
Repeat|7795,7801
echo|7802,7806
showed|7807,7813
improvement|7814,7825
of|7826,7828
her|7829,7832
<EOL>|7833,7834
mitral|7834,7840
regurgitation|7841,7854
.|7854,7855
<EOL>|7856,7857
<EOL>|7857,7858
#|7858,7859
NSTEMI|7860,7866
/|7866,7867
CAD|7867,7870
:|7870,7871
<EOL>|7871,7872
As|7872,7874
evidenced|7875,7884
by|7885,7887
EKG|7888,7891
changes|7892,7899
and|7900,7903
troponin|7904,7912
leak|7913,7917
.|7917,7918
Patient|7919,7926
was|7927,7930
<EOL>|7931,7932
briefly|7932,7939
started|7940,7947
on|7948,7950
a|7951,7952
heparin|7953,7960
drip|7961,7965
prior|7966,7971
to|7972,7974
her|7975,7978
first|7979,7984
cardiac|7985,7992
<EOL>|7993,7994
catheterization|7994,8009
.|8009,8010
As|8011,8013
above|8014,8019
,|8019,8020
cardiac|8021,8028
catheterization|8029,8044
revealed|8045,8053
<EOL>|8054,8055
3|8055,8056
-|8056,8057
vessel|8057,8063
disease|8064,8071
.|8071,8072
Patient|8073,8080
was|8081,8084
initially|8085,8094
medically|8095,8104
managed|8105,8112
with|8113,8117
<EOL>|8118,8119
aspirin|8119,8126
,|8126,8127
plavix|8128,8134
,|8134,8135
metoprolol|8136,8146
,|8146,8147
lisinopril|8148,8158
,|8158,8159
and|8160,8163
atorvastatin|8164,8176
.|8176,8177
As|8178,8180
<EOL>|8181,8182
the|8182,8185
patient|8186,8193
would|8194,8199
be|8200,8202
too|8203,8206
high|8207,8211
risk|8212,8216
for|8217,8220
CABG|8221,8225
,|8225,8226
patient|8227,8234
returned|8235,8243
to|8244,8246
<EOL>|8247,8248
the|8248,8251
cath|8252,8256
lab|8257,8260
and|8261,8264
had|8265,8268
a|8269,8270
bare|8271,8275
metal|8276,8281
stent|8282,8287
and|8288,8291
POBA|8292,8296
.|8296,8297
She|8298,8301
will|8302,8306
<EOL>|8307,8308
require|8308,8315
plavix|8316,8322
for|8323,8326
at|8327,8329
least|8330,8335
1|8336,8337
month|8338,8343
.|8343,8344
<EOL>|8344,8345
<EOL>|8345,8346
#|8346,8347
Hypertension|8348,8360
:|8360,8361
Patient|8362,8369
remained|8370,8378
normotensive|8379,8391
.|8391,8392
Continued|8393,8402
<EOL>|8403,8404
nifedipine|8404,8414
at|8415,8417
half|8418,8422
of|8423,8425
her|8426,8429
home|8430,8434
dose|8435,8439
.|8439,8440
Continued|8441,8450
on|8451,8453
lisinopril|8454,8464
.|8464,8465
<EOL>|8466,8467
She|8467,8470
was|8471,8474
also|8475,8479
started|8480,8487
on|8488,8490
metoprolol|8491,8501
as|8502,8504
above|8505,8510
for|8511,8514
CHF|8515,8518
.|8518,8519
<EOL>|8519,8520
<EOL>|8520,8521
#|8521,8522
Diabetes|8523,8531
:|8531,8532
Continued|8533,8542
home|8543,8547
insulin|8548,8555
regime|8556,8562
.|8562,8563
<EOL>|8564,8565
<EOL>|8566,8567
#|8567,8568
CKD|8569,8572
stage|8573,8578
IV|8579,8581
:|8581,8582
Baseline|8583,8591
Cr|8592,8594
2.5|8595,8598
-|8598,8599
2.8|8599,8602
per|8603,8606
renal|8607,8612
notes|8613,8618
.|8618,8619
Currently|8620,8629
<EOL>|8630,8631
at|8631,8633
baseline|8634,8642
.|8642,8643
<EOL>|8644,8645
<EOL>|8645,8646
#|8646,8647
History|8648,8655
of|8656,8658
CVA|8659,8662
:|8662,8663
Continued|8664,8673
home|8674,8678
aspirin|8679,8686
and|8687,8690
clopidogrel|8691,8702
.|8702,8703
<EOL>|8704,8705
<EOL>|8705,8706
#|8706,8707
GERD|8708,8712
:|8712,8713
Continued|8714,8723
home|8724,8728
ranitidine|8729,8739
.|8739,8740
<EOL>|8740,8741
<EOL>|8741,8742
TRANSITIONAL|8742,8754
ISSUES|8755,8761
:|8761,8762
<EOL>|8763,8764
*|8764,8765
Will|8766,8770
need|8771,8775
follow|8776,8782
up|8783,8785
with|8786,8790
a|8791,8792
cardiologist|8793,8805
.|8805,8806
Patient|8807,8814
will|8815,8819
be|8820,8822
<EOL>|8823,8824
scheduled|8824,8833
to|8834,8836
follow|8837,8843
up|8844,8846
with|8847,8851
the|8852,8855
first|8856,8861
available|8862,8871
CMED|8872,8876
<EOL>|8877,8878
cardiologist|8878,8890
.|8890,8891
<EOL>|8892,8893
*|8893,8894
Will|8895,8899
need|8900,8904
plavix|8905,8911
for|8912,8915
at|8916,8918
least|8919,8924
one|8925,8928
month|8929,8934
(|8935,8936
day|8936,8939
of|8940,8942
bare|8943,8947
metal|8948,8953
<EOL>|8954,8955
stent|8955,8960
placement|8961,8970
=|8971,8972
_|8973,8974
_|8974,8975
_|8975,8976
.|8976,8977
<EOL>|8977,8978
*|8978,8979
Atorvastatin|8980,8992
dose|8993,8997
increased|8998,9007
to|9008,9010
80mg|9011,9015
(|9016,9017
per|9017,9020
pharmacy|9021,9029
,|9029,9030
her|9031,9034
<EOL>|9035,9036
insurance|9036,9045
will|9046,9050
cover|9051,9056
.|9056,9057
Her|9058,9061
co-pay|9062,9068
will|9069,9073
be|9074,9076
$|9077,9078
10|9078,9080
/|9080,9081
month|9081,9086
)|9086,9087
.|9087,9088
<EOL>|9088,9089
*|9089,9090
Consider|9091,9099
titrating|9100,9109
nifedipine|9110,9120
dose|9121,9125
back|9126,9130
to|9131,9133
120mg|9134,9139
if|9140,9142
still|9143,9148
<EOL>|9149,9150
hypertensive|9150,9162
.|9162,9163
<EOL>|9164,9165
*|9165,9166
Please|9167,9173
recheck|9174,9181
Chem7|9182,9187
at|9188,9190
next|9191,9195
appointment|9196,9207
to|9208,9210
evaluate|9211,9219
for|9220,9223
_|9224,9225
_|9225,9226
_|9226,9227
<EOL>|9228,9229
secondary|9229,9238
to|9239,9241
dye|9242,9245
received|9246,9254
during|9255,9261
cardiac|9262,9269
catheterization|9270,9285
.|9285,9286
<EOL>|9286,9287
<EOL>|9288,9289
Medications|9289,9300
on|9301,9303
Admission|9304,9313
:|9313,9314
<EOL>|9314,9315
The|9315,9318
Preadmission|9319,9331
Medication|9332,9342
list|9343,9347
is|9348,9350
accurate|9351,9359
and|9360,9363
complete|9364,9372
.|9372,9373
<EOL>|9373,9374
1.|9374,9376
Lisinopril|9377,9387
30|9388,9390
mg|9391,9393
PO|9394,9396
DAILY|9397,9402
<EOL>|9403,9404
2.|9404,9406
NIFEdipine|9407,9417
CR|9418,9420
60|9421,9423
mg|9424,9426
PO|9427,9429
DAILY|9430,9435
<EOL>|9436,9437
3.|9437,9439
Ranitidine|9440,9450
300|9451,9454
mg|9455,9457
PO|9458,9460
DAILY|9461,9466
<EOL>|9467,9468
4.|9468,9470
Pravastatin|9471,9482
80|9483,9485
mg|9486,9488
PO|9489,9491
DAILY|9492,9497
<EOL>|9498,9499
5.|9499,9501
HumuLIN|9502,9509
70|9510,9512
/|9512,9513
30|9513,9515
(|9516,9517
insulin|9517,9524
NPH|9525,9528
and|9529,9532
regular|9533,9540
human|9541,9546
)|9546,9547
30|9548,9550
units|9551,9556
<EOL>|9557,9558
subcutaneous|9558,9570
daily|9571,9576
<EOL>|9577,9578
6.|9578,9580
Ferrous|9581,9588
Sulfate|9589,9596
325|9597,9600
mg|9601,9603
PO|9604,9606
BID|9607,9610
<EOL>|9611,9612
7.|9612,9614
Furosemide|9615,9625
40|9626,9628
mg|9629,9631
PO|9632,9634
DAILY|9635,9640
<EOL>|9641,9642
8.|9642,9644
Multivitamins|9645,9658
1|9659,9660
TAB|9661,9664
PO|9665,9667
DAILY|9668,9673
<EOL>|9674,9675
9.|9675,9677
Nitroglycerin|9678,9691
SL|9692,9694
0.3|9695,9698
mg|9699,9701
SL|9702,9704
PRN|9705,9708
chest|9709,9714
pain|9715,9719
<EOL>|9720,9721
10|9721,9723
.|9723,9724
DiphenhydrAMINE|9725,9740
25|9741,9743
mg|9744,9746
PO|9747,9749
HS|9750,9752
:|9752,9753
PRN|9753,9756
insomnia|9757,9765
<EOL>|9766,9767
11.|9767,9770
sevelamer|9771,9780
CARBONATE|9781,9790
800|9791,9794
mg|9795,9797
PO|9798,9800
TID|9801,9804
W|9805,9806
/|9806,9807
MEALS|9807,9812
<EOL>|9813,9814
12.|9814,9817
Clopidogrel|9818,9829
75|9830,9832
mg|9833,9835
PO|9836,9838
DAILY|9839,9844
(|9845,9846
was|9846,9849
not|9850,9853
taking|9854,9860
regularly|9861,9870
)|9870,9871
<EOL>|9871,9872
13.|9872,9875
Aspirin|9876,9883
81|9884,9886
mg|9887,9889
PO|9890,9892
DAILY|9893,9898
<EOL>|9899,9900
14.|9900,9903
Vitamin|9904,9911
D|9912,9913
_|9914,9915
_|9915,9916
_|9916,9917
UNIT|9918,9922
PO|9923,9925
DAILY|9926,9931
<EOL>|9932,9933
<EOL>|9933,9934
<EOL>|9935,9936
Discharge|9936,9945
Medications|9946,9957
:|9957,9958
<EOL>|9958,9959
1.|9959,9961
Aspirin|9962,9969
81|9970,9972
mg|9973,9975
PO|9976,9978
DAILY|9979,9984
<EOL>|9985,9986
2.|9986,9988
Clopidogrel|9989,10000
75|10001,10003
mg|10004,10006
PO|10007,10009
DAILY|10010,10015
<EOL>|10016,10017
3.|10017,10019
Furosemide|10020,10030
40|10031,10033
mg|10034,10036
PO|10037,10039
DAILY|10040,10045
<EOL>|10046,10047
4.|10047,10049
Lisinopril|10050,10060
30|10061,10063
mg|10064,10066
PO|10067,10069
DAILY|10070,10075
<EOL>|10076,10077
5.|10077,10079
Multivitamins|10080,10093
1|10094,10095
TAB|10096,10099
PO|10100,10102
DAILY|10103,10108
<EOL>|10109,10110
6.|10110,10112
Ranitidine|10113,10123
300|10124,10127
mg|10128,10130
PO|10131,10133
DAILY|10134,10139
<EOL>|10140,10141
7.|10141,10143
sevelamer|10144,10153
CARBONATE|10154,10163
800|10164,10167
mg|10168,10170
PO|10171,10173
TID|10174,10177
W|10178,10179
/|10179,10180
MEALS|10180,10185
<EOL>|10186,10187
8.|10187,10189
Atorvastatin|10190,10202
80|10203,10205
mg|10206,10208
PO|10209,10211
DAILY|10212,10217
<EOL>|10218,10219
RX|10219,10221
*|10222,10223
atorvastatin|10223,10235
80|10236,10238
mg|10239,10241
1|10242,10243
tablet|10244,10250
(|10250,10251
s|10251,10252
)|10252,10253
by|10254,10256
mouth|10257,10262
daily|10263,10268
Disp|10269,10273
#|10274,10275
*|10275,10276
30|10276,10278
<EOL>|10279,10280
Tablet|10280,10286
Refills|10287,10294
:|10294,10295
*|10295,10296
0|10296,10297
<EOL>|10297,10298
9.|10298,10300
Metoprolol|10301,10311
Succinate|10312,10321
XL|10322,10324
25|10325,10327
mg|10328,10330
PO|10331,10333
DAILY|10334,10339
<EOL>|10340,10341
RX|10341,10343
*|10344,10345
metoprolol|10345,10355
succinate|10356,10365
25|10366,10368
mg|10369,10371
1|10372,10373
tablet|10374,10380
extended|10381,10389
release|10390,10397
24|10398,10400
<EOL>|10401,10402
hr|10402,10404
(|10404,10405
s|10405,10406
)|10406,10407
by|10408,10410
mouth|10411,10416
daily|10417,10422
Disp|10423,10427
#|10428,10429
*|10429,10430
30|10430,10432
Tablet|10433,10439
Refills|10440,10447
:|10447,10448
*|10448,10449
0|10449,10450
<EOL>|10450,10451
10.|10451,10454
DiphenhydrAMINE|10455,10470
25|10471,10473
mg|10474,10476
PO|10477,10479
HS|10480,10482
:|10482,10483
PRN|10483,10486
insomnia|10487,10495
<EOL>|10496,10497
11|10497,10499
.|10499,10500
HumuLIN|10501,10508
70|10509,10511
/|10511,10512
30|10512,10514
(|10515,10516
insulin|10516,10523
NPH|10524,10527
and|10528,10531
regular|10532,10539
human|10540,10545
)|10545,10546
30|10547,10549
units|10550,10555
<EOL>|10556,10557
subcutaneous|10557,10569
daily|10570,10575
<EOL>|10576,10577
12.|10577,10580
Nitroglycerin|10581,10594
SL|10595,10597
0.3|10598,10601
mg|10602,10604
SL|10605,10607
PRN|10608,10611
chest|10612,10617
pain|10618,10622
<EOL>|10623,10624
13|10624,10626
.|10626,10627
Vitamin|10628,10635
D|10636,10637
_|10638,10639
_|10639,10640
_|10640,10641
UNIT|10642,10646
PO|10647,10649
DAILY|10650,10655
<EOL>|10656,10657
14.|10657,10660
NIFEdipine|10661,10671
CR|10672,10674
60|10675,10677
mg|10678,10680
PO|10681,10683
DAILY|10684,10689
<EOL>|10690,10691
<EOL>|10691,10692
<EOL>|10693,10694
Discharge|10694,10703
Disposition|10704,10715
:|10715,10716
<EOL>|10716,10717
Home|10717,10721
With|10722,10726
Service|10727,10734
<EOL>|10734,10735
<EOL>|10736,10737
Facility|10737,10745
:|10745,10746
<EOL>|10746,10747
_|10747,10748
_|10748,10749
_|10749,10750
<EOL>|10750,10751
<EOL>|10752,10753
Discharge|10753,10762
Diagnosis|10763,10772
:|10772,10773
<EOL>|10773,10774
Severe|10793,10799
mitral|10800,10806
regurgitation|10807,10820
<EOL>|10820,10821
Coronary|10821,10829
artery|10830,10836
disease|10837,10844
<EOL>|10844,10845
<EOL>|10845,10846
SECONDARY|10846,10855
DIAGNOSIS|10856,10865
:|10865,10866
<EOL>|10866,10867
Hypertension|10867,10879
<EOL>|10879,10880
Diabetes|10880,10888
<EOL>|10888,10889
<EOL>|10889,10890
<EOL>|10891,10892
Mental|10913,10919
Status|10920,10926
:|10926,10927
Clear|10928,10933
and|10934,10937
coherent|10938,10946
.|10946,10947
<EOL>|10947,10948
Level|10948,10953
of|10954,10956
Consciousness|10957,10970
:|10970,10971
Alert|10972,10977
and|10978,10981
interactive|10982,10993
.|10993,10994
<EOL>|10994,10995
Activity|10995,11003
Status|11004,11010
:|11010,11011
Ambulatory|11012,11022
-|11023,11024
Independent|11025,11036
.|11036,11037
<EOL>|11037,11038
<EOL>|11038,11039
<EOL>|11040,11041
Dear|11065,11069
Ms.|11070,11073
_|11074,11075
_|11075,11076
_|11076,11077
,|11077,11078
<EOL>|11078,11079
<EOL>|11079,11080
It|11080,11082
was|11083,11086
a|11087,11088
pleasure|11089,11097
caring|11098,11104
for|11105,11108
you|11109,11112
at|11113,11115
_|11116,11117
_|11117,11118
_|11118,11119
<EOL>|11120,11121
_|11121,11122
_|11122,11123
_|11123,11124
.|11124,11125
As|11126,11128
you|11129,11132
recall|11133,11139
,|11139,11140
you|11141,11144
were|11145,11149
admitted|11150,11158
for|11159,11162
shortness|11163,11172
<EOL>|11173,11174
of|11174,11176
breath|11177,11183
.|11183,11184
This|11185,11189
was|11190,11193
because|11194,11201
one|11202,11205
of|11206,11208
your|11209,11213
heart|11214,11219
valves|11220,11226
was|11227,11230
weak|11231,11235
,|11235,11236
<EOL>|11237,11238
which|11238,11243
caused|11244,11250
fluid|11251,11256
to|11257,11259
build|11260,11265
up|11266,11268
in|11269,11271
your|11272,11276
lungs|11277,11282
.|11282,11283
Your|11284,11288
heart|11289,11294
valve|11295,11300
<EOL>|11301,11302
was|11302,11305
weak|11306,11310
because|11311,11318
there|11319,11324
was|11325,11328
a|11329,11330
blockage|11331,11339
in|11340,11342
one|11343,11346
of|11347,11349
your|11350,11354
heart|11355,11360
<EOL>|11361,11362
arteries|11362,11370
.|11370,11371
You|11372,11375
underwent|11376,11385
a|11386,11387
procedure|11388,11397
,|11397,11398
called|11399,11405
cardiac|11406,11413
<EOL>|11414,11415
catheterization|11415,11430
,|11430,11431
which|11432,11437
opened|11438,11444
up|11445,11447
the|11448,11451
blocked|11452,11459
arteries|11460,11468
.|11468,11469
Your|11470,11474
<EOL>|11475,11476
valve|11476,11481
and|11482,11485
heart|11486,11491
are|11492,11495
pumping|11496,11503
much|11504,11508
more|11509,11513
efficiently|11514,11525
now|11526,11529
.|11529,11530
We|11531,11533
are|11534,11537
<EOL>|11538,11539
glad|11539,11543
you|11544,11547
are|11548,11551
feeling|11552,11559
better|11560,11566
.|11566,11567
Please|11568,11574
weigh|11575,11580
yourself|11581,11589
every|11590,11595
<EOL>|11596,11597
morning|11597,11604
,|11604,11605
and|11606,11609
call|11610,11614
your|11615,11619
MD|11620,11622
if|11623,11625
your|11626,11630
weight|11631,11637
goes|11638,11642
up|11643,11645
more|11646,11650
than|11651,11655
3|11656,11657
lbs|11658,11661
<EOL>|11662,11663
over|11663,11667
24|11668,11670
hours|11671,11676
.|11676,11677
<EOL>|11677,11678
<EOL>|11679,11680
Followup|11680,11688
Instructions|11689,11701
:|11701,11702
<EOL>|11702,11703
_|11703,11704
_|11704,11705
_|11705,11706
<EOL>|11706,11707

