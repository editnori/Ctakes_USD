CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|true|false||Unit
null|Unit device|Device|true|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|true|false||Unit
null|Unit of Measure|LabModifier|true|false||Unit
null|Unit|LabModifier|true|false||Unit
null|Enzyme Unit|LabModifier|true|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Neurosurgical Procedures|Procedure|false|false||NEUROSURGERYnull|Science of neurosurgery|Title|false|false||NEUROSURGERYnull|penicillins|Drug|false|false||Penicillins
null|penicillins|Drug|false|false||Penicillinsnull|Poisoning by, adverse effect of and underdosing of penicillins|Disorder|false|false||Penicillins
null|Poisoning by penicillin|Disorder|false|false||Penicillinsnull|Adverse reaction to penicillins|Finding|false|false||Penicillinsnull|Paxil|Drug|false|false||Paxil
null|Paxil|Drug|false|false||Paxilnull|Wellbutrin|Drug|false|false||Wellbutrin
null|Wellbutrin|Drug|false|false||Wellbutrinnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Computer Hardware Device|Device|false|false||hardware
null|Diagnostic, Therapeutic, and Research Equipment|Device|false|false||hardwarenull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Hardware Removal|Procedure|false|false||hardware removalnull|Computer Hardware Device|Device|false|false||hardware
null|Diagnostic, Therapeutic, and Research Equipment|Device|false|false||hardwarenull|removal technique|Procedure|false|false||removal
null|Excision|Procedure|false|false||removal
null|Extraction|Procedure|false|false||removalnull|Removing (action)|Event|false|false||removalnull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Old|Time|false|false||oldnull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|History of surgery|Finding|false|false||prior surgerynull|null|Time|false|false||priornull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Possible|Finding|false|false||possiblenull|Possible diagnosis|Modifier|false|false||possible
null|Possibly Related to Intervention|Modifier|false|false||possiblenull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Parietal|Modifier|false|false||parietalnull|Anaplastic astrocytoma|Disorder|false|false||anaplastic astrocytomanull|Undifferentiated|Modifier|false|false||anaplasticnull|Astrocytoma|Disorder|false|false||astrocytomanull|Craniotomy|Procedure|false|false||craniotomynull|removal technique|Procedure|false|false||resection
null|Excision|Procedure|false|false||resectionnull|Involvement with|Finding|false|false||involvednull|Involved Anatomy|Modifier|false|false||involvednull|Knowledge Field|Finding|false|false||field
null|Force Field|Finding|false|false||field
null|Field|Finding|false|false||fieldnull|field - patient encounter|Procedure|false|false||fieldnull|Radiation therapy (procedure)|Procedure|false|false||irradiationnull|Irradiation (physical force)|Phenomenon|false|false||irradiation
null|Radiation|Phenomenon|false|false||irradiationnull|cGy|LabModifier|false|false||cGynull|event cycle|Time|false|false||cyclesnull|Temodar|Drug|false|false||Temodar
null|Temodar|Drug|false|false||Temodarnull|Precision - second|Finding|false|false||second
null|metastatic qualifier|Finding|false|false||second
null|Second Suffix|Finding|false|false||secondnull|seconds|Time|false|false||secondnull|Second Unit of Plane Angle|LabModifier|false|false||second
null|second (number)|LabModifier|false|false||secondnull|Craniotomy|Procedure|false|false||craniotomynull|Recurrent tumor|Disorder|false|false||tumor recurrencenull|Neoplasms|Disorder|false|false||tumornull|Tumor Mass|Finding|false|false||tumor
null|null|Finding|false|false||tumornull|Recurrent Malignant Neoplasm|Disorder|false|false||recurrencenull|Recurrence (disease attribute)|Finding|false|false||recurrencenull|Recurrence|Phenomenon|false|false||recurrencenull|penciclovir|Drug|false|false||PCV
null|penciclovir|Drug|false|false||PCVnull|Porcine circovirus|Disorder|false|false||PCVnull|Procarbazine-Lomustine-Vincristine (PCV) Regimen|Procedure|false|false||PCV
null|lomustine/procarbazine/vincristine|Procedure|false|false||PCV
null|Hematocrit Measurement|Procedure|false|false||PCVnull|area PCV|Anatomy|false|false||PCVnull|After Dinner|Time|false|false||PCVnull|Combid|Drug|false|false||comb
null|Combid|Drug|false|false||combnull|bleomycin/cyclophosphamide/methotrexate/vincristine protocol|Procedure|false|false||comb
null|bleomycin/cyclophosphamide/semustine/vincristine protocol|Procedure|false|false||combnull|Comb (body structure)|Anatomy|false|false||combnull|Comb (physical object)|Device|false|false||combnull|Chemotherapy Regimen|Procedure|false|false||chemo
null|Chemotherapy|Procedure|false|false||chemonull|Diagnostic, Therapeutic, and Research Equipment|Device|false|false||hardware
null|Computer Hardware Device|Device|false|false||hardwarenull|Address type - Office|Finding|false|false||officenull|Office|Device|false|false||officenull|Organization unit type - Office|Entity|false|false||officenull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|complex (molecular entity)|Drug|false|false||complexnull|Complex|Modifier|false|false||complexnull|Revision procedure|Procedure|false|false||revision
null|Surgical revision|Procedure|false|false||revisionnull|Revision|Time|false|false||revisionnull|Plate Device|Device|false|false||plate
null|Bone plates|Device|false|false||plate
null|Device Plate|Device|false|false||platenull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false||skinnull|Skin Specimen Source Code|Finding|false|false||skin
null|Skin Specimen|Finding|false|false||skinnull|Skin, Human|Anatomy|false|false||skin
null|Skin|Anatomy|false|false||skinnull|Plastics|Drug|false|false||Plasticsnull|Scalp structure|Anatomy|false|false||scalpnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Pruritus|Finding|false|false||pruritusnull|sensory perception of itch|Modifier|false|false||pruritusnull|Problems with head|Disorder|false|false||headnull|Procedure on head|Procedure|false|false||headnull|Structure of head of caudate nucleus|Anatomy|false|false||head
null|Head|Anatomy|false|false||headnull|Head Device|Device|false|false||headnull|Newly Diagnosed|Modifier|false|false||newly diagnosednull|newly|Finding|false|false||newlynull|Diagnostic, Therapeutic, and Research Equipment|Device|false|false||hardware
null|Computer Hardware Device|Device|false|false||hardwarenull|husband|Subject|false|false||husbandnull|Problems with head|Disorder|false|false||headnull|Procedure on head|Procedure|false|false||headnull|Structure of head of caudate nucleus|Anatomy|false|false||head
null|Head|Anatomy|false|false||headnull|Head Device|Device|false|false||headnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|Metals|Drug|false|false||metalnull|Diagnostic, Therapeutic, and Research Equipment|Device|false|false||hardware
null|Computer Hardware Device|Device|false|false||hardwarenull|History of surgery|Finding|false|false||prior surgerynull|null|Time|false|false||priornull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Parietal|Modifier|false|false||parietalnull|Anaplastic astrocytoma|Disorder|false|false||anaplastic astrocytomanull|Undifferentiated|Modifier|false|false||anaplasticnull|Astrocytoma|Disorder|false|false||astrocytomanull|Craniotomy|Procedure|false|false||Craniotomynull|Radiation therapy (procedure)|Procedure|false|false||irradiationnull|Irradiation (physical force)|Phenomenon|false|false||irradiation
null|Radiation|Phenomenon|false|false||irradiationnull|cGy|LabModifier|false|false||cGynull|event cycle|Time|false|false||cyclesnull|Temodar|Drug|false|false||Temodar
null|Temodar|Drug|false|false||Temodarnull|Craniotomy|Procedure|false|false||craniotomynull|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic Wound|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|Revision procedure|Procedure|false|false||revision
null|Surgical revision|Procedure|false|false||revisionnull|Revision|Time|false|false||revisionnull|removal technique|Procedure|false|false||removal
null|Excision|Procedure|false|false||removal
null|Extraction|Procedure|false|false||removalnull|Removing (action)|Event|false|false||removalnull|Computer Hardware Device|Device|false|false||hardware
null|Diagnostic, Therapeutic, and Research Equipment|Device|false|false||hardwarenull|Accutane|Drug|false|false||Accutane
null|Accutane|Drug|false|false||Accutanenull|2 Weeks|Time|false|false||2 weeksnull|week|Time|false|false||weeksnull|Disease|Disorder|false|false||diseasenull|Tubal Ligation|Procedure|false|false||tubal ligationnull|Ligation|Procedure|false|false||ligationnull|Tonsillectomy|Procedure|false|false||tonsillectomynull|Acute bronchitis|Disorder|false|false||bronchitis
null|Bronchitis|Disorder|false|false||bronchitisnull|Cancer patients and suicide and depression|Disorder|false|false||depression
null|Mental Depression|Disorder|false|false||depression
null|Depressive disorder|Disorder|false|false||depression
null|Depressed mood|Disorder|false|false||depressionnull|Depression - motion|Finding|false|false||depression
null|null|Finding|false|false||depressionnull|Depression - recess|Modifier|false|false||depressionnull|Seizures|Finding|false|false||seizuresnull|Obesity|Disorder|false|false||obesenull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Gen
null|GEN1 wt Allele|Finding|false|false||Gen
null|GEN1 gene|Finding|false|false||Gennull|Feeling comfortable|Finding|false|false||comfortablenull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|HEENT|Anatomy|false|false||HEENTnull|Extraocular|Finding|false|false||EOMsnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Passive joint movement of neck (finding)|Finding|false|false||Neck
null|Neck problem|Finding|false|false||Necknull|dendritic spine neck|Anatomy|false|false||Neck
null|Neck|Anatomy|false|false||Necknull|Supple|Finding|false|false||Supplenull|Dyspnea|Finding|true|false||SOBnull|Obesity|Disorder|true|false||obesenull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|Mental state|Finding|false|false||Mental statusnull|null|Attribute|false|false||Mental status
null|null|Attribute|false|false||Mental statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|Alert brand of caffeine|Drug|false|false||alert
null|Alert brand of caffeine|Drug|false|false||alertnull|Mentally alert|Finding|false|false||alert
null|Consciousness clear|Finding|false|false||alert
null|Alert note|Finding|false|false||alert
null|Alert|Finding|false|false||alertnull|null|Attribute|false|false||alertnull|cooperative|Entity|false|false||cooperativenull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Affect (mental function)|Finding|false|false||affectnull|assessment of affect|Procedure|false|false||affectnull|LITAF gene|Finding|false|false||simplenull|Simple|Modifier|false|false||simplenull|Recombinant DNA|Drug|false|false||constructnull|Construct|Finding|false|false||constructnull|Mental Orientation|Finding|false|false||Orientationnull|Orientation, Spatial|Modifier|false|false||Orientation
null|Genomic Orientation|Modifier|false|false||Orientation
null|Orientation|Modifier|false|false||Orientationnull|Oriented to person|Finding|false|false||Oriented to personnull|Oriented to place|Finding|false|false||Orientednull|Orientation, Spatial|Modifier|false|false||Orientednull|Person Info|Finding|false|false||personnull|null|Attribute|false|false||personnull|Persons|Subject|false|false||personnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Mental Recall|Finding|false|false||Recallnull|Recall (activity)|Event|false|false||Recallnull|Physical object|Entity|false|false||objectsnull|5 minutes Office visit|Procedure|false|false||5 minutesnull|5 minutes|Time|false|false||5 minutesnull|Minute of time|Time|false|false||minutesnull|Minute Unit of Plane Angle|LabModifier|false|false||minutes
null|Minute (diminutive)|LabModifier|false|false||minutes
null|Small|LabModifier|false|false||minutesnull|Programming Languages|Finding|false|false||Languagenull|null|Attribute|false|false||Languagenull|Languages|Entity|false|false||Languagenull|Speech|Finding|false|false||Speechnull|Speech assessment|Procedure|false|false||Speechnull|Language Ability Proficiency - Good|Finding|false|false||good
null|Language Proficiency - Good|Finding|false|false||goodnull|Specimen Quality - Good|Modifier|false|false||good
null|Good|Modifier|false|false||goodnull|Comprehension|Finding|false|false||comprehensionnull|speech fluency repetition (physical finding)|Finding|false|false||repetition
null|Repeat|Finding|false|false||repetitionnull|Naming (function)|Finding|false|false||Namingnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Dysarthria|Disorder|true|false||dysarthrianull|error|Modifier|true|false||errorsnull|Neoplasm of uncertain or unknown behavior of cranial nerves|Disorder|false|false||Cranial Nerves
null|Benign neoplasm of cranial nerves|Disorder|false|false||Cranial Nervesnull|Cranial Nerves|Anatomy|false|false||Cranial Nervesnull|Bone structure of cranium|Anatomy|false|false||Cranialnull|Cranial|Modifier|false|false||Cranialnull|Nerve|Anatomy|false|false||Nervesnull|Pupil|Anatomy|false|false||Pupilsnull|Round shape|Modifier|false|false||roundnull|Reactive to light|Finding|false|false||reactive to lightnull|Reactive Therapy|Procedure|false|false||reactivenull|Reactive|Modifier|false|false||reactivenull|TNFSF14 protein, human|Drug|false|false||light
null|TNFSF14 protein, human|Drug|false|false||lightnull|Light - subjective measurement|Finding|false|false||light
null|TNFSF14 wt Allele|Finding|false|false||light
null|TNFSF14 gene|Finding|false|false||light
null|Light color|Finding|false|false||lightnull|Phototherapy|Procedure|false|false||lightnull|Light|Phenomenon|false|false||lightnull|Light (qualifier)|Modifier|false|false||lightnull|Visual Fields|Modifier|false|false||Visual fieldsnull|Visual|Finding|false|false||Visualnull|Full|Modifier|false|false||fullnull|Social confrontation skill|Finding|false|false||confrontationnull|Confrontation visual field test|Procedure|false|false||confrontation
null|Confrontation|Procedure|false|false||confrontationnull|examination of extraocular movements|Procedure|true|false||Extraocular movementsnull|Extraocular|Finding|true|false||Extraocularnull|Movement|Finding|true|false||movementsnull|Gender Status - Intact|Finding|true|false||intactnull|Intact|Modifier|true|false||intactnull|Nystagmus|Disorder|true|false||nystagmusnull|Roman numeral VII|Finding|false|false||VIInull|Lamina VII of gray matter of spinal cord|Anatomy|false|false||VII
null|lobule VII|Anatomy|false|false||VII
null|layer VII (Cajal)|Anatomy|false|false||VIInull|Face|Anatomy|false|false||Facialnull|Facial|Modifier|false|false||Facialnull|Strength (attribute)|Finding|false|false||strengthnull|Pharmaceutical Strength|LabModifier|false|false||strength
null|Physical Strength|LabModifier|false|false||strengthnull|Observation of Sensation|Finding|false|false||sensation
null|Sensory perception|Finding|false|false||sensationnull|sensory exam|Procedure|false|false||sensationnull|Sensation quality|Modifier|false|false||sensationnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Symmetric Relationship|Finding|false|false||symmetric
null|Symmetrical|Finding|false|false||symmetricnull|Roman numeral VIII|Finding|false|false||VIII
null|COX8A gene|Finding|false|false||VIIInull|Lamina VIII of gray matter of spinal cord|Anatomy|false|false||VIII
null|Cerebellar pyramis|Anatomy|false|false||VIIInull|outcomes otolaryngology hearing|Finding|false|false||Hearing
null|Hearing finding|Finding|false|false||Hearing
null|Hearing|Finding|false|false||Hearingnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Authorization Mode - Voice|Finding|false|false||voice
null|Voice G-code|Finding|false|false||voice
null|Voice|Finding|false|false||voicenull|TelecommunicationCapabilities - voice|Modifier|false|false||voicenull|Palate|Anatomy|false|false||Palatalnull|Elevation procedure|Procedure|false|false||elevationnull|Elevation|Modifier|false|false||elevationnull|Symmetrical|Finding|false|false||symmetricalnull|Structure of sternocleidomastoid muscle|Anatomy|false|false||Sternocleidomastoidnull|Structure of trapezius muscle|Anatomy|false|false||trapeziusnull|tongue midline|Finding|true|false||Tongue midlinenull|Benign neoplasm of tongue|Disorder|true|false||Tonguenull|Procedure on tongue|Procedure|true|false||Tonguenull|Tongue|Anatomy|true|false||Tonguenull|midline cell component|Anatomy|true|false||midlinenull|Midline (qualifier value)|Modifier|true|false||midlinenull|Muscular fasciculation|Finding|true|false||fasciculationsnull|motor movement|Finding|false|false||Motornull|Motor Device|Device|false|false||Motornull|Bulk (conceptual)|Drug|false|false||bulk
null|Dietary Fiber|Drug|false|false||bulknull|Dyskinetic syndrome|Disorder|true|false||abnormal movementsnull|Abnormal movement|Finding|true|false||abnormal movementsnull|Observation Interpretation - Abnormal|Finding|true|false||abnormal
null|Abnormal|Finding|true|false||abnormalnull|Movement|Finding|true|false||movementsnull|Academic Research Enhancement Awards|Event|false|false||areanull|Geographic Locations|Entity|false|false||areanull|Area|Modifier|false|false||areanull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false||skinnull|Skin Specimen Source Code|Finding|false|false||skin
null|Skin Specimen|Finding|false|false||skinnull|Skin, Human|Anatomy|false|false||skin
null|Skin|Anatomy|false|false||skinnull|THYROID HORMONE PLASMA MEMBRANE TRANSPORT DEFECT|Disorder|false|false||defectnull|Defect|Finding|false|false||defectnull|Underlying|Finding|false|false||underlyingnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false||skinnull|Skin Specimen Source Code|Finding|false|false||skin
null|Skin Specimen|Finding|false|false||skinnull|Skin, Human|Anatomy|false|false||skin
null|Skin|Anatomy|false|false||skinnull|Different|Modifier|false|false||Differentnull|Act Relationship Subset - previous|Time|false|false||previous
null|Previous|Time|false|false||previousnull|Part|Modifier|false|false||portionnull|Piece Unit|LabModifier|false|false||piecenull|Body Substance Discharge|Finding|true|false||discharge
null|Discharge Body Fluid|Finding|true|false||discharge
null|Body Fluid Discharge|Finding|true|false||discharge
null|null|Finding|true|false||dischargenull|Patient Discharge|Procedure|true|false||dischargenull|Swelling|Finding|true|false||swelling
null|Edema|Finding|true|false||swellingnull|Benign|Modifier|false|false||benignnull|Aspect (characteristic)|Modifier|false|false||aspectnull|Aspect - Kind of quantity|LabModifier|false|false||aspectnull|physical examination (physical finding)|Finding|false|false||PHYSICAL EXAMnull|Physical Examination|Procedure|false|false||PHYSICAL EXAMnull|physical examination (physical finding)|Finding|false|false||PHYSICAL
null|Physical|Finding|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||PHYSICALnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|null|Time|false|false||PRIOR TOnull|null|Time|false|false||PRIORnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Obesity|Disorder|false|false||obesenull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Gen
null|GEN1 wt Allele|Finding|false|false||Gen
null|GEN1 gene|Finding|false|false||Gennull|Feeling comfortable|Finding|false|false||comfortablenull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|HEENT|Anatomy|false|false||HEENTnull|Extraocular|Finding|false|false||EOMsnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Passive joint movement of neck (finding)|Finding|false|false||Neck
null|Neck problem|Finding|false|false||Necknull|dendritic spine neck|Anatomy|false|false||Neck
null|Neck|Anatomy|false|false||Necknull|Supple|Finding|false|false||Supplenull|Surgical wound|Disorder|false|false||Incisionnull|Surgical incisions|Procedure|false|false||Incisionnull|Cranial incision point|Anatomy|false|false||Incisionnull|Cleaning (activity)|Event|false|false||cleannull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Erythema|Disorder|true|false||rednessnull|Redness|Finding|true|false||rednessnull|Red color|Modifier|true|false||rednessnull|Swelling|Finding|true|false||swelling
null|Edema|Finding|true|false||swellingnull|Erythema|Disorder|true|false||erythemanull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Suture Joint|Anatomy|false|false||Suturesnull|Surgical sutures|Device|false|false||Suturesnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Diagnostic Service Section ID - Hematology|Finding|false|false||Hematologynull|diagnostic service sources hematology (procedure)|Procedure|false|false||Hematology
null|Hematology procedure|Procedure|false|false||Hematology
null|Hematologic Tests|Procedure|false|false||Hematologynull|hematology (field)|Title|false|false||Hematologynull|Complete Blood Count|Procedure|false|false||COMPLETE BLOOD COUNTnull|Complete, Multiple Vitamins with Iron|Drug|false|false||COMPLETE
null|Complete, Multiple Vitamins with Iron|Drug|false|false||COMPLETE
null|Complete, Multiple Vitamins with Iron|Drug|false|false||COMPLETEnull|Completion Status for valid values - Complete|Finding|false|false||COMPLETE
null|Data operation - complete|Finding|false|false||COMPLETE
null|Finish - dosing instruction imperative|Finding|false|false||COMPLETEnull|Complete|Modifier|false|false||COMPLETEnull|Blood Cell Count|Procedure|false|false||BLOOD COUNTnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Count Dosing Unit|LabModifier|false|false||COUNT
null|Count|LabModifier|false|false||COUNTnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Base|Drug|false|false||BASICnull|Basis - conceptual entity|Finding|false|false||BASICnull|Basic (cigarettes)|Device|false|false||BASICnull|Coagulation process|Finding|false|false||COAGULATION
null|Blood coagulation|Finding|false|false||COAGULATIONnull|Observation Method - Coagulation|Procedure|false|false||COAGULATION
null|Coagulation procedure|Procedure|false|false||COAGULATION
null|Blood coagulation tests|Procedure|false|false||COAGULATIONnull|Blood coagulation pathway observation|Lab|false|false||COAGULATIONnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Primed lymphocyte test|Procedure|false|false||PLTnull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|Primed lymphocyte test|Procedure|false|false||Pltnull|diagnostic service sources chemistry (fluid analysis)|Finding|false|false||Chemistry
null|chemical aspects|Finding|false|false||Chemistry
null|Chemistry Section ID|Finding|false|false||Chemistrynull|Chemical procedure|Procedure|false|false||Chemistrynull|Science of Chemistry|Subject|false|false||Chemistrynull|Urologic Diseases|Disorder|false|false||RENALnull|Kidney|Anatomy|false|false||RENALnull|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSEnull|Glucose measurement|Procedure|false|false||GLUCOSEnull|Glucose^1.5H post dose glucagon|Lab|false|false||GLUCOSEnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Neurosurgical service|Entity|false|false||neurosurgical servicenull|ActInformationPrivacyReason - service|Finding|false|false||servicenull|Software Service|Device|false|false||servicenull|Services|Event|false|false||servicenull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|Computer Hardware Device|Device|false|false||hardware
null|Diagnostic, Therapeutic, and Research Equipment|Device|false|false||hardwarenull|Act Relationship Subset - previous|Time|false|false||previous
null|Previous|Time|false|false||previousnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Problems with head|Disorder|false|false||headnull|Procedure on head|Procedure|false|false||headnull|Structure of head of caudate nucleus|Anatomy|false|false||head
null|Head|Anatomy|false|false||headnull|Head Device|Device|false|false||headnull|removal technique|Procedure|false|false||removal
null|Excision|Procedure|false|false||removal
null|Extraction|Procedure|false|false||removalnull|Removing (action)|Event|false|false||removalnull|Computer Hardware Device|Device|false|false||hardware
null|Diagnostic, Therapeutic, and Research Equipment|Device|false|false||hardwarenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Communicable Diseases|Disorder|false|false||Infectious diseasenull|Infectious Disease Medicine|Title|false|false||Infectious diseasenull|Communicable Diseases|Disorder|false|false||Infectiousnull|infectious - Entity Risk|Modifier|false|false||Infectiousnull|Disease|Disorder|false|false||diseasenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|INJECTION FLUCONAZOLE, 200 MG ADMINISTERED|Drug|false|false||fluconazole
null|fluconazole|Drug|false|false||fluconazole
null|fluconazole|Drug|false|false||fluconazolenull|5 Days|Time|false|false||5 daysnull|day|Time|false|false||daysnull|Yeast infection|Disorder|false|false||yeast infectionnull|Yeast, Dried|Drug|false|false||yeast
null|Candida albicans allergenic extract|Drug|false|false||yeast
null|Candida albicans allergenic extract|Drug|false|false||yeast
null|Candida albicans allergenic extract|Drug|false|false||yeastnull|Saccharomyces cerevisiae|Entity|false|false||yeast
null|Yeasts|Entity|false|false||yeastnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Keflex|Drug|false|false||Keflex
null|Keflex|Drug|false|false||Keflexnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|7 days|Time|false|false||7 daysnull|day|Time|false|false||daysnull|DVT prophylaxis|Procedure|false|false||DVT prophylaxisnull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|Prophylactic treatment|Procedure|false|false||prophylaxisnull|prevention & control|Modifier|false|false||prophylaxisnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|subcutaneous heparin|Drug|false|false||subcutaneous heparin
null|subcutaneous heparin|Drug|false|false||subcutaneous heparinnull|Subcutaneous Route of Administration|Finding|false|false||subcutaneousnull|subcutaneous|Modifier|false|false||subcutaneousnull|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|SCD protein, human|Drug|false|false||SCD
null|SCD protein, human|Drug|false|false||SCDnull|Schnyder crystalline corneal dystrophy|Disorder|false|false||SCD
null|Renal carnitine transport defect|Disorder|false|false||SCD
null|Anemia, Sickle Cell|Disorder|false|false||SCDnull|SCD gene|Finding|false|false||SCD
null|Doctor of Science|Finding|false|false||SCD
null|Sudden Cardiac Death|Finding|false|false||SCD
null|SLC22A5 gene|Finding|false|false||SCDnull|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|Agreement (document)|Finding|false|false||agreement
null|Agreement|Finding|false|false||agreementnull|null|Attribute|false|false||agreementnull|Comprehension|Finding|false|false||understandingnull|Discharge plan|Finding|false|false||discharge plannull|Discharge Planning|Procedure|false|false||discharge plannull|null|Attribute|false|false||discharge plannull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Infantile Neuroaxonal Dystrophy|Disorder|false|false||plannull|Treatment Plan|Finding|false|false||plan
null|Planned|Finding|false|false||plan
null|null|Finding|false|false||plannull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Inaccurate|Modifier|false|false||inaccuratenull|Act Class - investigation|Finding|false|false||investigationnull|Evaluation procedure|Procedure|false|false||investigation
null|Evaluation|Procedure|false|false||investigationnull|alprazolam|Drug|false|false||ALPRAZolam
null|alprazolam|Drug|false|false||ALPRAZolamnull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|azathioprine|Drug|false|false||Azathioprine
null|azathioprine|Drug|false|false||Azathioprine
null|azathioprine|Drug|false|false||Azathioprinenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|dicyclomine|Drug|false|false||DiCYCLOmine
null|dicyclomine|Drug|false|false||DiCYCLOminenull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Abdominal Pain|Finding|false|false||abdominal painnull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Fluticasone-Salmeterol Diskus|Drug|false|false||Fluticasone-Salmeterol Diskus
null|Fluticasone-Salmeterol Diskus|Drug|false|false||Fluticasone-Salmeterol Diskusnull|fluticasone / salmeterol|Drug|false|false||Fluticasone-Salmeterolnull|fluticasone|Drug|false|false||Fluticasone
null|fluticasone|Drug|false|false||Fluticasonenull|salmeterol|Drug|false|false||Salmeterol
null|salmeterol|Drug|false|false||Salmeterolnull|Diskus|Device|false|false||Diskusnull|Inhalant dose form|Drug|false|false||INH
null|isoniazid|Drug|false|false||INH
null|isoniazid|Drug|false|false||INHnull|Inhalation Route of Administration|Finding|false|false||INHnull|Ingush language|Entity|false|false||INHnull|Inhalation Dosing Unit|LabModifier|false|false||INHnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|hydrocodone|Drug|false|false||Hydrocodone
null|hydrocodone|Drug|false|false||Hydrocodonenull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|Every four hours|Time|false|false||Q4Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|infliximab|Drug|false|false||Infliximab
null|infliximab|Drug|false|false||Infliximab
null|infliximab|Drug|false|false||Infliximabnull|Drug assay infliximab|Procedure|false|false||Infliximabnull|week|Time|false|false||WEEKSnull|levothyroxine sodium|Drug|false|false||Levothyroxine Sodium
null|levothyroxine sodium|Drug|false|false||Levothyroxine Sodium
null|levothyroxine sodium|Drug|false|false||Levothyroxine Sodiumnull|Synthetic Levothyroxine|Drug|false|false||Levothyroxine
null|Synthetic Levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxinenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|microgram|LabModifier|false|false||mcgnull|Daily|Time|false|false||DAILYnull|mesalamine|Drug|false|false||Mesalamine
null|mesalamine|Drug|false|false||Mesalaminenull|Four times daily|Time|false|false||QIDnull|omeprazole|Drug|false|false||Omeprazole
null|omeprazole|Drug|false|false||Omeprazolenull|Daily|Time|false|false||DAILYnull|promethazine|Drug|false|false||Promethazine
null|promethazine|Drug|false|false||Promethazinenull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Topamax|Drug|false|false||Topiramate (Topamax)
null|Topamax|Drug|false|false||Topiramate (Topamax)null|topiramate|Drug|false|false||Topiramate
null|topiramate|Drug|false|false||Topiramatenull|Topiramate measurement|Procedure|false|false||Topiramatenull|Topamax|Drug|false|false||Topamax
null|Topamax|Drug|false|false||Topamaxnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|venlafaxine|Drug|false|false||Venlafaxine
null|venlafaxine|Drug|false|false||Venlafaxinenull|Daily|Time|false|false||DAILYnull|zolpidem tartrate|Drug|false|false||Zolpidem Tartrate
null|zolpidem tartrate|Drug|false|false||Zolpidem Tartratenull|zolpidem|Drug|false|false||Zolpidem
null|zolpidem|Drug|false|false||Zolpidemnull|tartrate|Drug|false|false||Tartrate
null|Tartrates|Drug|false|false||Tartrate
null|tartrate|Drug|false|false||Tartratenull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|alprazolam|Drug|false|false||ALPRAZolam
null|alprazolam|Drug|false|false||ALPRAZolamnull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|azathioprine|Drug|false|false||Azathioprine
null|azathioprine|Drug|false|false||Azathioprine
null|azathioprine|Drug|false|false||Azathioprinenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|dicyclomine|Drug|false|false||DiCYCLOmine
null|dicyclomine|Drug|false|false||DiCYCLOminenull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Abdominal Pain|Finding|false|false||abdominal painnull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|levothyroxine sodium|Drug|false|false||Levothyroxine Sodium
null|levothyroxine sodium|Drug|false|false||Levothyroxine Sodium
null|levothyroxine sodium|Drug|false|false||Levothyroxine Sodiumnull|Synthetic Levothyroxine|Drug|false|false||Levothyroxine
null|Synthetic Levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxinenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|microgram|LabModifier|false|false||mcgnull|Daily|Time|false|false||DAILYnull|mesalamine|Drug|false|false||Mesalamine
null|mesalamine|Drug|false|false||Mesalaminenull|Four times daily|Time|false|false||QIDnull|omeprazole|Drug|false|false||Omeprazole
null|omeprazole|Drug|false|false||Omeprazolenull|Daily|Time|false|false||DAILYnull|Topamax|Drug|false|false||Topiramate (Topamax)
null|Topamax|Drug|false|false||Topiramate (Topamax)null|topiramate|Drug|false|false||Topiramate
null|topiramate|Drug|false|false||Topiramatenull|Topiramate measurement|Procedure|false|false||Topiramatenull|Topamax|Drug|false|false||Topamax
null|Topamax|Drug|false|false||Topamaxnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|venlafaxine|Drug|false|false||Venlafaxine
null|venlafaxine|Drug|false|false||Venlafaxinenull|Daily|Time|false|false||DAILYnull|zolpidem tartrate|Drug|false|false||Zolpidem Tartrate
null|zolpidem tartrate|Drug|false|false||Zolpidem Tartratenull|zolpidem|Drug|false|false||Zolpidem
null|zolpidem|Drug|false|false||Zolpidemnull|tartrate|Drug|false|false||Tartrate
null|Tartrates|Drug|false|false||Tartrate
null|tartrate|Drug|false|false||Tartratenull|hydrocodone|Drug|false|false||Hydrocodone
null|hydrocodone|Drug|false|false||Hydrocodonenull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|Every four hours|Time|false|false||Q4Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Body temperature measurement|Procedure|false|false||temperaturenull|Body Temperature|Subject|false|false||temperaturenull|Temperature|LabModifier|false|false||temperaturenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Constipation|Finding|false|false||constipationnull|docusate sodium|Drug|false|false||docusate sodium
null|docusate sodium|Drug|false|false||docusate sodiumnull|docusate|Drug|false|false||docusate
null|docusate|Drug|false|false||docusatenull|Sodium supplements|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|Sodium Drug Class|Drug|false|false||sodiumnull|Sodium metabolic function|Finding|false|false||sodiumnull|Sodium measurement|Procedure|false|false||sodiumnull|capsule (pharmacologic)|Drug|false|false||capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||capsule
null|Structure of organ capsule|Anatomy|false|false||capsulenull|Capsule Shape|Modifier|false|false||capsulenull|Capsule (unit of presentation)|LabModifier|false|false||capsule
null|Capsule Dosing Unit|LabModifier|false|false||capsulenull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Twice a day|Time|false|false||twice a daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|refill|Finding|false|false||Refillsnull|INJECTION FLUCONAZOLE, 200 MG ADMINISTERED|Drug|false|false||Fluconazole
null|fluconazole|Drug|false|false||Fluconazole
null|fluconazole|Drug|false|false||Fluconazolenull|Every twenty four hours|Time|false|false||Q24Hnull|Duration brand of oxymetazoline|Drug|false|false||Durationnull|Duration (temporal concept)|Time|false|false||Durationnull|4 Days|Time|false|false||4 Daysnull|day|Time|false|false||Daysnull|INJECTION FLUCONAZOLE, 200 MG ADMINISTERED|Drug|false|false||fluconazole
null|fluconazole|Drug|false|false||fluconazole
null|fluconazole|Drug|false|false||fluconazolenull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Daily|Time|false|false||dailynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|oxycodone|Drug|false|false||OxycoDONE
null|oxycodone|Drug|false|false||OxycoDONEnull|Oxycodone measurement|Procedure|false|false||OxycoDONEnull|Immediate Release Dosage Form|Drug|false|false||Immediate Releasenull|Query Priority - Immediate|Finding|false|false||Immediate
null|immediate - ResponseCode|Finding|false|false||Immediatenull|Immediate|Time|false|false||Immediate
null|Stat (do immediately)|Time|false|false||Immediatenull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Moderate - Severity of Illness Code|Finding|false|false||moderate
null|Moderate|Finding|false|false||moderatenull|Moderate (severity modifier)|Modifier|false|false||moderate
null|Moderate - Allergy Severity|Modifier|false|false||moderate
null|Moderation|Modifier|false|false||moderatenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|oxycodone|Drug|false|false||oxycodone
null|oxycodone|Drug|false|false||oxycodonenull|Oxycodone measurement|Procedure|false|false||oxycodonenull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Hour|Time|false|false||hoursnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|cephalexin|Drug|false|false||Cephalexin
null|cephalexin|Drug|false|false||Cephalexinnull|Every twelve hours|Time|false|false||Q12Hnull|Duration brand of oxymetazoline|Drug|false|false||Durationnull|Duration (temporal concept)|Time|false|false||Durationnull|7 days|Time|false|false||7 Daysnull|day|Time|false|false||Daysnull|cephalexin|Drug|false|false||cephalexin
null|cephalexin|Drug|false|false||cephalexinnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Twice a day|Time|false|false||twice a daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Hardware Removal|Procedure|false|false||Hardware removalnull|Computer Hardware Device|Device|false|false||Hardware
null|Diagnostic, Therapeutic, and Research Equipment|Device|false|false||Hardwarenull|removal technique|Procedure|false|false||removal
null|Excision|Procedure|false|false||removal
null|Extraction|Procedure|false|false||removalnull|Removing (action)|Event|false|false||removalnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|INJECTION FLUCONAZOLE, 200 MG ADMINISTERED|Drug|false|false||Fluconazole
null|fluconazole|Drug|false|false||Fluconazole
null|fluconazole|Drug|false|false||Fluconazolenull|Once daily|Time|false|false||once dailynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Daily|Time|false|false||dailynull|4 Days|Time|false|false||4 daysnull|day|Time|false|false||daysnull|Keflex|Drug|false|false||Keflex
null|Keflex|Drug|false|false||Keflexnull|7 days|Time|false|false||7 daysnull|day|Time|false|false||daysnull|Wound Infection|Finding|false|false||wound infectionnull|Traumatic Wound|Disorder|false|false||wound
null|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Clearance procedure|Procedure|false|false||Clearancenull|Clearance of substance|Attribute|false|false||Clearancenull|Clearance [PK]|Phenomenon|false|false||Clearancenull|Clearance|Modifier|false|false||Clearancenull|Intrinsic drive|Finding|false|false||drivenull|Work|Event|false|false||worknull|Postoperative Period|Time|false|false||post-operativenull|Office Visits|Procedure|false|false||office visitnull|Address type - Office|Finding|false|false||officenull|Office|Device|false|false||officenull|Organization unit type - Office|Entity|false|false||officenull|Visit|Finding|false|false||visitnull|Call - dosing instruction fragment|Finding|false|false||CALL
null|Call (Instruction)|Finding|false|false||CALL
null|Decision|Finding|false|false||CALL
null|CHL1 gene|Finding|false|false||CALLnull|null|Attribute|false|false||SURGEONnull|Surgeon|Subject|false|false||SURGEONnull|Stat (do immediately)|Time|false|false||IMMEDIATELYnull|Experience (Practice)|Finding|true|false||EXPERIENCE
null|Experience|Finding|true|false||EXPERIENCEnull|Following|Time|true|false||FOLLOWING
null|Status post|Time|true|false||FOLLOWINGnull|new onset|Finding|false|false||New onsetnull|Query Status Code - new|Finding|false|false||New
null|Act Status - new|Finding|false|false||Newnull|Newar Language|Entity|false|false||Newnull|New|Modifier|false|false||Newnull|Onset of (contextual qualifier)|Modifier|false|false||onset ofnull|Onset of (contextual qualifier)|Modifier|false|false||onsetnull|Age of Onset|LabModifier|false|false||onsetnull|Tremor|Finding|false|false||tremorsnull|Seizures|Finding|false|false||seizuresnull|Confusion|Disorder|true|false||confusionnull|Clouded consciousness|Finding|true|false||confusionnull|Mental status changes|Finding|true|false||change in mental statusnull|null|Attribute|true|false||change in mental statusnull|Changing|Finding|true|false||change innull|Changed status|LabModifier|true|false||change innull|Changing|Finding|true|false||changenull|Change - procedure|Procedure|true|false||changenull|Changed status|LabModifier|true|false||change
null|Delta (difference)|LabModifier|true|false||changenull|Mental state|Finding|true|false||mental statusnull|null|Attribute|true|false||mental status
null|null|Attribute|true|false||mental statusnull|Psyche structure|Finding|true|false||mentalnull|What subject filter - Status|Finding|true|false||statusnull|null|Attribute|true|false||statusnull|Social status|Modifier|true|false||status
null|Status|Modifier|true|false||statusnull|Numbness|Finding|true|false||numbness
null|Hypesthesia|Finding|true|false||numbnessnull|Paresthesia|Disorder|true|false||tinglingnull|Has tingling sensation|Finding|true|false||tinglingnull|Weakness|Finding|true|false||weakness
null|Asthenia|Finding|true|false||weaknessnull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Headache|Finding|true|false||headachenull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Pharmaceutical Preparations|Drug|true|false||medicationnull|medication - HL7 publishing domain|Finding|true|false||medication
null|Medications|Finding|true|false||medicationnull|Aspects of signs|Finding|true|false||signs
null|Physical findings|Finding|true|false||signsnull|Manufactured sign|Device|true|false||signsnull|Communicable Diseases|Disorder|true|false||infectionnull|Infection|Finding|true|false||infectionnull|Traumatic Wound|Disorder|true|false||wound
null|Wounds and Injuries|Disorder|true|false||wound
null|Traumatic injury|Disorder|true|false||woundnull|Route of Administration - Wound|Finding|true|false||wound
null|null|Finding|true|false||wound
null|Specimen Type - Wound|Finding|true|false||woundnull|null|Finding|true|false||sitenull|Anatomic Site|Anatomy|true|false||sitenull|Study Site|Modifier|true|false||site
null|Site|Modifier|true|false||sitenull|Erythema|Disorder|false|false||rednessnull|Redness|Finding|false|false||rednessnull|Red color|Modifier|false|false||rednessnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Emotional tenderness|Finding|false|false||tenderness
null|Sore to touch|Finding|false|false||tendernessnull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|Fever symptoms (finding)|Finding|false|false||Fever
null|Fever|Finding|false|false||Fevernull|Greater Than or Equal To|LabModifier|false|false||greater than or equal tonull|Greater Than or Equal To|LabModifier|false|false||greater than or equalnull|Greater Than|LabModifier|false|false||greater thannull|Greater|LabModifier|false|false||greaternull|Equal|Modifier|false|false||equal tonull|Relational Operator - Equal|Finding|false|false||equalnull|Equal|Modifier|false|false||equalnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions