CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|omeprazole|Drug|false|false||omeprazole
null|omeprazole|Drug|false|false||omeprazolenull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Chief complaint (finding)|Finding|false|false||Chief Complaintnull|Complaint (finding)|Finding|false|false||Complaintnull|null|Attribute|false|false||Complaintnull|Deglutition Disorders|Disorder|false|false||dysphagianull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Upper Surface|Modifier|false|false||Upper
null|Upper|Modifier|false|false||Uppernull|Endoscopy, Gastrointestinal|Procedure|false|false||endoscopy
null|Endoscopy (procedure)|Procedure|false|false||endoscopynull|History of present illness (finding)|Finding|false|false||History of Present Illnessnull|null|Attribute|false|false||History of Present Illnessnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Present illness|Finding|false|false||Present Illnessnull|Present|Finding|false|false||Present
null|Presentation|Finding|false|false||Presentnull|Illness (finding)|Finding|false|false||Illnessnull|Anxiety Disorders|Disorder|false|false||anxiety
null|Anxiety|Disorder|false|false||anxietynull|Anxiety symptoms|Finding|false|false||anxietynull|Several|LabModifier|false|false||severalnull|year|Time|false|false||yearsnull|Deglutition Disorders|Disorder|false|false||dysphagianull|Got Worse|Finding|false|false||worsened
null|Worse|Finding|false|false||worsenednull|Foreign body sensation (finding)|Finding|false|false|C0460148;C0444584;C4082212;C1268086;C0152338|foreign body sensation
null|Foreign body sensation in eyes|Finding|false|false|C0460148;C0444584;C4082212;C1268086;C0152338|foreign body sensationnull|Foreign Bodies|Disorder|false|false|C0460148;C0444584;C4082212;C1268086;C0152338|foreign bodynull|Foreign body (physical object)|Entity|false|false||foreign bodynull|International Aspects|Finding|false|false|C0460148;C0444584;C4082212;C1268086;C0152338|foreignnull|foreign|Modifier|false|false||foreignnull|Document Body|Finding|false|false|C0460148;C0444584;C4082212;C1268086;C0152338|bodynull|Structure of body of caudate nucleus|Anatomy|false|false|C0036658;C0542538;C0016542;C0920171;C0423602;C0376327;C1551342;C2229507|body
null|Human body structure|Anatomy|false|false|C0036658;C0542538;C0016542;C0920171;C0423602;C0376327;C1551342;C2229507|body
null|Body structure|Anatomy|false|false|C0036658;C0542538;C0016542;C0920171;C0423602;C0376327;C1551342;C2229507|body
null|Adult human body|Anatomy|false|false|C0036658;C0542538;C0016542;C0920171;C0423602;C0376327;C1551342;C2229507|body
null|Whole body|Anatomy|false|false|C0036658;C0542538;C0016542;C0920171;C0423602;C0376327;C1551342;C2229507|bodynull|Human body|Subject|false|false||bodynull|Observation of Sensation|Finding|false|false|C0460148;C0444584;C4082212;C1268086;C0152338|sensation
null|Sensory perception|Finding|false|false|C0460148;C0444584;C4082212;C1268086;C0152338|sensationnull|sensory exam|Procedure|false|false|C0460148;C0444584;C4082212;C1268086;C0152338|sensationnull|Sensation quality|Modifier|false|false||sensationnull|Food allergenic extracts|Drug|false|false||food
null|Food|Drug|false|false||food
null|Food allergenic extracts|Drug|false|false||foodnull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|neck
null|Neck problem|Finding|false|false|C0027530;C3159206|necknull|dendritic spine neck|Anatomy|false|false|C0812434;C0684335|neck
null|Neck|Anatomy|false|false|C0812434;C0684335|necknull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Last|Modifier|false|false||lastnull|10 days|Time|false|false||10 daysnull|day|Time|false|false||daysnull|Food allergenic extracts|Drug|false|false|C0230069;C3665375;C0031354|food
null|Food|Drug|false|false|C0230069;C3665375;C0031354|food
null|Food allergenic extracts|Drug|false|false|C0230069;C3665375;C0031354|foodnull|Throat Homeopathic Medication|Drug|false|false|C0230069;C3665375;C0031354|throatnull|Specimen Type - Throat|Finding|false|false|C0230069;C3665375;C0031354|throat
null|null|Finding|false|false|C0230069;C3665375;C0031354|throatnull|Throat|Anatomy|false|false|C1950455;C1550663;C1547926;C3540798;C0016452|throat
null|Anterior portion of neck|Anatomy|false|false|C1950455;C1550663;C1547926;C3540798;C0016452|throat
null|Pharyngeal structure|Anatomy|false|false|C1950455;C1550663;C1547926;C3540798;C0016452|throatnull|Nearly|Modifier|false|false||almostnull|Breath|Finding|false|false||breathnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Medical History|Finding|true|false||history ofnull|History of present illness (finding)|Finding|true|false||history
null|History of previous events|Finding|true|false||history
null|Historical aspects qualifier|Finding|true|false||history
null|Medical History|Finding|true|false||history
null|Concept History|Finding|true|false||historynull|History|Subject|false|false||historynull|Food Allergy|Disorder|true|false||food allergiesnull|Food allergenic extracts|Drug|false|false||food
null|Food|Drug|false|false||food
null|Food allergenic extracts|Drug|false|false||foodnull|Hypersensitivity|Finding|false|false||allergiesnull|null|Attribute|false|false||allergiesnull|Skin rash|Finding|false|false|C1123023;C4520765|skin rashesnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765|skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765|skinnull|Skin Specimen Source Code|Finding|false|false|C1123023;C4520765|skin
null|Skin Specimen|Finding|false|false|C1123023;C4520765|skinnull|Skin, Human|Anatomy|false|false|C1546781;C0444099;C0178298;C0496955;C5779628|skin
null|Skin|Anatomy|false|false|C1546781;C0444099;C0178298;C0496955;C5779628|skinnull|Skin rash|Finding|false|false||rashes
null|Exanthema|Finding|false|false||rashesnull|Initial (abbreviation)|Finding|false|false||initialnull|Initially|Time|false|false||initialnull|Firstly|Modifier|false|false||initialnull|Imaging problem|Finding|false|false||Imagingnull|Diagnostic Imaging|Procedure|false|false||Imaging
null|Imaging Techniques|Procedure|false|false||Imagingnull|Imaging Technology|Title|false|false||Imagingnull|Plain chest X-ray|Procedure|false|false||CXRnull|Prominent|Modifier|false|false||prominentnull|Carcinoma in situ of esophagus|Disorder|false|false|C4266613;C0014876|esophagus
null|Esophageal Diseases|Disorder|false|false|C4266613;C0014876|esophagus
null|Benign neoplasm of esophagus|Disorder|false|false|C4266613;C0014876|esophagusnull|Esophagus problem|Finding|false|false|C4266613;C0014876|esophagusnull|Procedures on the esophagus|Procedure|false|false|C4266613;C0014876|esophagusnull|Chest>Esophagus|Anatomy|false|false|C0812418;C0872395;C0014852;C0154059;C0153942|esophagus
null|Esophagus|Anatomy|false|false|C0812418;C0872395;C0014852;C0154059;C0153942|esophagusnull|Consultation|Procedure|false|false||Consultsnull|Esophagogastroduodenoscopy|Procedure|false|false|C4266613;C0014876|EGDnull|Carcinoma in situ of esophagus|Disorder|false|false|C4266613;C0014876|esophagus
null|Esophageal Diseases|Disorder|false|false|C4266613;C0014876|esophagus
null|Benign neoplasm of esophagus|Disorder|false|false|C4266613;C0014876|esophagusnull|Esophagus problem|Finding|false|false|C4266613;C0014876|esophagusnull|Procedures on the esophagus|Procedure|false|false|C4266613;C0014876|esophagusnull|Chest>Esophagus|Anatomy|false|false|C0872395;C0812418;C0079304;C0014852;C0154059;C0153942|esophagus
null|Esophagus|Anatomy|false|false|C0872395;C0812418;C0079304;C0014852;C0154059;C0153942|esophagusnull|Biopsy|Procedure|false|false||Biopsiesnull|Current (present time)|Time|false|false||Currentlynull|Anxiety Disorders|Disorder|false|false||anxiety
null|Anxiety|Disorder|false|false||anxietynull|Anxiety symptoms|Finding|false|false||anxietynull|null|Time|false|false||prior tonull|null|Time|false|false||priornull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Gastroesophageal reflux disease|Disorder|false|false||GERDnull|Hypercholesterolemia|Disorder|false|false||Hypercholesterolemianull|Hypercholesterolemia result|Finding|false|false||Hypercholesterolemianull|NEPHROLITHIASIS, CALCIUM OXALATE, 1|Disorder|false|false|C0227665;C0022646|Kidney stones
null|Nephrolithiasis|Disorder|false|false|C0227665;C0022646|Kidney stonesnull|Kidney Calculi|Finding|false|false|C0227665;C0022646|Kidney stonesnull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false|C0227665;C0022646|Kidney
null|Benign neoplasm of kidney|Disorder|false|false|C0227665;C0022646|Kidneynull|Kidney problem|Finding|false|false|C0227665;C0022646|Kidneynull|examination of kidney|Procedure|false|false|C0227665;C0022646|Kidney
null|Procedures on Kidney|Procedure|false|false|C0227665;C0022646|Kidneynull|Kidney|Anatomy|false|false|C0496927;C0496892;C0022650;C0812426;C4554465;C0869841;C0006736;C0392525;C5779632|Kidney
null|Both kidneys|Anatomy|false|false|C0496927;C0496892;C0022650;C0812426;C4554465;C0869841;C0006736;C0392525;C5779632|Kidneynull|Calculi|Finding|false|false|C0227665;C0022646|stonesnull|stones - unit|LabModifier|false|false||stonesnull|Mitral Valve Prolapse Syndrome|Disorder|false|false|C1186983;C0026264|Mitral valve prolapsenull|Mitral Valve|Anatomy|false|false|C0033377;C0026267|Mitral valvenull|mitral|Modifier|false|false||Mitralnull|Anatomical valve|Anatomy|false|false|C0026267;C0033377|valvenull|Valve (physical object)|Device|false|false||valve
null|Valve Device|Device|false|false||valve
null|medical valve|Device|false|false||valvenull|Ptosis|Disorder|false|false|C0026264;C1186983|prolapsenull|Uterine Fibroids|Disorder|false|false|C0042149|Uterine fibroidsnull|Uterus|Anatomy|false|false|C0042133;C0023267;C0042133|Uterinenull|Uterine Fibroids|Disorder|false|false|C0042149|fibroids
null|Fibroid Tumor|Disorder|false|false|C0042149|fibroidsnull|Osteoporosis|Disorder|false|false||Osteoporosisnull|Encounter due to family history of osteoporosis|Finding|false|false||Osteoporosisnull|Migraine Disorders|Disorder|false|false||Migraine headachesnull|Migraine Disorders|Disorder|false|false||Migrainenull|Headache|Finding|false|false||headachesnull|Social and personal history|Finding|false|false||Social History
null|Social History|Finding|false|false||Social Historynull|Social|Finding|false|false||Socialnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Family Medical History|Finding|false|false||Family Historynull|Entity Name Part Type - family|Finding|false|false||Family
null|Last Name|Finding|false|false||Family
null|Living Arrangement - Family|Finding|false|false||Family
null|Family (taxonomic)|Finding|false|false||Family
null|Family Collection|Finding|false|false||Familynull|Family|Subject|false|false||Familynull|History of present illness (finding)|Finding|false|true||History
null|History of previous events|Finding|false|true||History
null|Historical aspects qualifier|Finding|false|true||History
null|Medical History|Finding|false|true||History
null|Concept History|Finding|false|true||Historynull|History|Subject|false|false||Historynull|Hypertensive disease|Disorder|false|false||HTNnull|Indirect exposure mechanism - Father|Finding|false|false||father
null|Relationship - Father|Finding|false|false||father
null|Father - courtesy title|Finding|false|false||fathernull|Father (person)|Subject|false|false||fathernull|Presenile dementia|Disorder|false|false||Dementia
null|Dementia|Disorder|false|false||Dementianull|Indirect exposure mechanism - Father|Finding|false|false||father
null|Relationship - Father|Finding|false|false||father
null|Father - courtesy title|Finding|false|false||fathernull|Father (person)|Subject|false|false||fathernull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GEN
null|GEN1 wt Allele|Finding|false|false||GEN
null|GEN1 gene|Finding|false|false||GENnull|Anxiety|Disorder|false|false||anxiousnull|Woman|Subject|false|false||woman
null|Human, Female adult|Subject|false|false||womannull|BORNHOLM EYE DISEASE|Disorder|false|false||bednull|Bachelor of Education|Finding|false|false||bednull|Beds|Device|false|false||bednull|Patient Location - Bed|Modifier|false|false||bednull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|false|false||acutenull|Emotional distress|Finding|true|false||distress
null|Distress|Finding|true|false||distressnull|HEENT|Anatomy|false|false||HEENTnull|Moist|Modifier|false|false||Moistnull|Anicteric|Finding|false|false||anictericnull|Pupil equal round and reacting to light|Finding|false|false||PERRLnull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|NECK
null|Neck problem|Finding|false|false|C0027530;C3159206|NECKnull|dendritic spine neck|Anatomy|false|false|C0812434;C0684335|NECK
null|Neck|Anatomy|false|false|C0812434;C0684335|NECKnull|Supple|Finding|false|false|C0226032|Supplenull|Leukocyte adhesion deficiency type 1|Disorder|true|false|C0226032|LAD
null|Leukocyte adhesion deficiency|Disorder|true|false|C0226032|LADnull|ITGB2 wt Allele|Finding|true|false|C0226032|LAD
null|DLD gene|Finding|true|false|C0226032|LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false|C5550999;C0398738;C1414063;C1706333;C0332254|LADnull|Ladino Language|Entity|true|false||LADnull|Jugular venous engorgement|Finding|true|false||JVDnull|Pulmonary ventilator management|Procedure|false|false||PULMnull|cordycepin|Drug|false|false|C0018787|COR
null|cordycepin|Drug|false|false|C0018787|CORnull|Heart|Anatomy|false|false|C0056331|CORnull|Cornish language|Entity|false|false||CORnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false|C0449202;C0000726|ABDnull|ABD (body structure)|Anatomy|false|false|C3811055|ABD
null|Abdomen|Anatomy|false|false|C3811055|ABDnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|LRRC4B gene|Finding|true|false||HSMnull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Neurology speciality|Title|false|false||NEUROnull|Neurologic (qualifier value)|Modifier|false|false||NEUROnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Motor function (finding)|Finding|false|false||motor functionnull|Motor function (observable entity)|Phenomenon|false|false||motor functionnull|motor movement|Finding|false|false||motornull|Motor Device|Device|false|false||motornull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|Observation of Sensation|Finding|false|false||sensation
null|Sensory perception|Finding|false|false||sensationnull|sensory exam|Procedure|false|false||sensationnull|Sensation quality|Modifier|false|false||sensationnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0005768;C0229664;C0005767;C0851353|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C0014792;C1114281|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false|C1185650|ALT
null|Atypical Lipoma|Disorder|false|false|C1185650|ALTnull|null|Finding|false|false|C1185650|ALT
null|Alternative Billing Concepts|Finding|false|false|C1185650|ALT
null|GPT gene|Finding|false|false|C1185650|ALTnull|Antibiotic Lock Therapy|Procedure|false|false|C1185650|ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|ASTnull|Atypical Spitz Nevus|Disorder|false|false|C1185650|ASTnull|SLC17A5 wt Allele|Finding|false|false|C1185650|AST
null|SLC17A5 gene|Finding|false|false|C1185650|AST
null|GOT1 gene|Finding|false|false|C1185650|ASTnull|Asterion|Anatomy|false|false|C2257651;C1415274;C1140170;C0202113;C0851148;C1415181;C1420113;C5960784;C1266129;C1370889;C4522245;C0004002;C0242192;C1121182;C4553172|ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Lactate Dehydrogenase|Drug|false|false||LDH
null|Lactate Dehydrogenase|Drug|false|false||LDHnull|Lifetime Drinking History|Finding|false|false|C1185650|LDHnull|Lactate dehydrogenase measurement|Procedure|false|false|C1185650|LDHnull|Alkaline Phosphatase|Drug|false|false||AlkPhos
null|Alkaline Phosphatase|Drug|false|false||AlkPhosnull|Blood albumin|Procedure|false|false||BLOOD Albuminnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Albumin|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumin|Drug|false|false||Albuminnull|Albumin metabolic function|Finding|false|false||Albumin
null|ALB gene|Finding|false|false||Albuminnull|Albumin measurement|Procedure|false|false||Albuminnull|Imaging problem|Finding|false|false||IMAGINGnull|Diagnostic Imaging|Procedure|false|false||IMAGING
null|Imaging Techniques|Procedure|false|false||IMAGINGnull|Imaging Technology|Title|false|false||IMAGINGnull|Plain chest X-ray|Procedure|false|false||CXRnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Prominent|Modifier|false|false||Prominentnull|Carcinoma in situ of esophagus|Disorder|false|false|C4266613;C0014876|esophagus
null|Esophageal Diseases|Disorder|false|false|C4266613;C0014876|esophagus
null|Benign neoplasm of esophagus|Disorder|false|false|C4266613;C0014876|esophagusnull|Esophagus problem|Finding|false|false|C4266613;C0014876|esophagusnull|Procedures on the esophagus|Procedure|false|false|C4266613;C0014876|esophagusnull|Chest>Esophagus|Anatomy|false|false|C0872395;C0812418;C2681903;C1140091;C1866503;C0014852;C0154059;C0153942|esophagus
null|Esophagus|Anatomy|false|false|C0872395;C0812418;C2681903;C1140091;C1866503;C0014852;C0154059;C0153942|esophagusnull|Lateral|Modifier|false|false||lateralnull|View|Modifier|false|false||viewnull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false|C4266613;C0014876|air
null|AIRN gene|Finding|false|false|C4266613;C0014876|air
null|AI/RHEUM|Finding|false|false|C4266613;C0014876|airnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Radiographic|Phenomenon|false|false||radiographicnull|patient appearance regarding mental status exam|Procedure|false|false||appearancenull|null|Attribute|false|false||appearancenull|Personal appearance|Subject|false|false||appearancenull|Appearance|Modifier|false|false||appearancenull|Kind of quantity - Appearance|LabModifier|false|false||appearancenull|barium|Drug|false|false||bariumnull|Swallow - dosing instruction imperative|Finding|false|false||swallow
null|Swallow (administration method)|Finding|false|false||swallownull|Family Hirundinidae|Entity|false|false||swallownull|Neck X-ray|Procedure|false|false|C0027530;C3159206|NECK X-ray
null|Radiographic procedure on neck|Procedure|false|false|C0027530;C3159206|NECK X-raynull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|NECK
null|Neck problem|Finding|false|false|C0027530;C3159206|NECKnull|dendritic spine neck|Anatomy|false|false|C0043309;C1963529;C0202757;C0034571;C3244296;C0043299;C1962945;C1306645;C0812434;C0684335|NECK
null|Neck|Anatomy|false|false|C0043309;C1963529;C0202757;C0034571;C3244296;C0043299;C1962945;C1306645;C0812434;C0684335|NECKnull|ActClaimAttachmentCategoryCode - x-ray|Finding|false|false|C0027530;C3159206|X-ray
null|roentgenographic|Finding|false|false|C0027530;C3159206|X-raynull|Plain x-ray|Procedure|false|false|C0027530;C3159206|X-ray
null|Diagnostic radiologic examination|Procedure|false|false|C0027530;C3159206|X-ray
null|Radiographic imaging procedure|Procedure|false|false|C0027530;C3159206|X-raynull|Roentgen Rays|Phenomenon|false|false|C0027530;C3159206|X-raynull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Limitation|Finding|false|false||limitation
null|Restricted|Finding|false|false||limitationnull|Plain x-ray|Procedure|false|false||plain radiographynull|roentgenographic|Finding|false|false||radiographynull|Diagnostic radiologic examination|Procedure|false|false||radiography
null|Radiographic imaging procedure|Procedure|false|false||radiography
null|Radiographic Examination|Procedure|false|false||radiographynull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Soft tissue swelling|Disorder|false|false|C0040300;C0225317;C4532079|soft tissue swellingnull|Neck+Chest>Soft tissue|Anatomy|false|false|C1547928;C3542022;C0013604;C0038999;C0037580|soft tissue
null|soft tissue|Anatomy|false|false|C1547928;C3542022;C0013604;C0038999;C0037580|soft tissuenull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false|C0225317;C4532079|softnull|Soft|Modifier|false|false||softnull|Tissue Specimen Code|Finding|false|false|C0225317;C4532079;C0040300|tissuenull|Body tissue|Anatomy|false|false|C1547928;C0037580;C0013604;C0038999|tissuenull|Swelling|Finding|false|false|C0040300;C0225317;C4532079|swelling
null|Edema|Finding|false|false|C0040300;C0225317;C4532079|swellingnull|Soft tissue mass|Disorder|false|false|C0040300;C0225317;C4532079|soft tissue massnull|Neck+Chest>Soft tissue|Anatomy|false|false|C3542022;C4283905;C1546709;C2700045;C0577573;C0577559;C1414542;C0457193;C1547928|soft tissue
null|soft tissue|Anatomy|false|false|C3542022;C4283905;C1546709;C2700045;C0577573;C0577559;C1414542;C0457193;C1547928|soft tissuenull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false|C0225317;C4532079;C0040300|softnull|Soft|Modifier|false|false||softnull|Tissue Specimen Code|Finding|false|false|C0040300;C0225317;C4532079|tissuenull|Body tissue|Anatomy|false|false|C0457193;C3542022;C1547928;C4283905;C1546709;C2700045;C0577573;C0577559;C1414542|tissuenull|Mass of body structure|Finding|false|false|C0225317;C4532079;C0040300|mass
null|Morphology, Attenuation, Size, and Structure Criteria|Finding|false|false|C0225317;C4532079;C0040300|mass
null|null|Finding|false|false|C0225317;C4532079;C0040300|mass
null|FBN1 wt Allele|Finding|false|false|C0225317;C4532079;C0040300|mass
null|FBN1 gene|Finding|false|false|C0225317;C4532079;C0040300|mass
null|Mass of body region|Finding|false|false|C0225317;C4532079;C0040300|massnull|Mass, a measure of quantity of matter|LabModifier|false|false||mass
null|Molecular Mass|LabModifier|false|false||massnull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|neck
null|Neck problem|Finding|false|false|C0027530;C3159206|necknull|dendritic spine neck|Anatomy|false|false|C0812434;C0684335|neck
null|Neck|Anatomy|false|false|C0812434;C0684335|necknull|Esophagogastroduodenoscopy|Procedure|false|false||EGDnull|impression (attitude)|Finding|false|false||Impression
null|EKG impression|Finding|false|false||Impressionnull|Hiatal Hernia|Disorder|false|false||Hiatal hernianull|Hernia|Disorder|false|false||hernianull|Angiectasis|Disorder|false|false|C3714551;C0038351;C4266636|Angioectasianull|Carcinoma in situ of stomach|Disorder|false|false|C3714551;C0038351;C4266636|stomach
null|Stomach Diseases|Disorder|false|false|C3714551;C0038351;C4266636|stomach
null|Benign neoplasm of stomach|Disorder|false|false|C3714551;C0038351;C4266636|stomach
null|Neoplasm of uncertain or unknown behavior of stomach|Disorder|false|false|C3714551;C0038351;C4266636|stomachnull|Stomach problem|Finding|false|false|C3714551;C0038351;C4266636|stomachnull|Procedure on stomach|Procedure|false|false|C3714551;C0038351;C4266636|stomachnull|Stomach structure|Anatomy|false|false|C0002959;C0038354;C0496905;C0153943;C0154060;C0872393;C0577027|stomach
null|Abdomen>Stomach|Anatomy|false|false|C0002959;C0038354;C0496905;C0153943;C0154060;C0872393;C0577027|stomach
null|Stomach|Anatomy|false|false|C0002959;C0038354;C0496905;C0153943;C0154060;C0872393;C0577027|stomachnull|Angiectasis|Disorder|false|false|C0013303|Angioectasianull|Malignant neoplasm of duodenum|Disorder|false|false|C0013303|duodenum
null|Benign neoplasm of duodenum|Disorder|false|false|C0013303|duodenumnull|Duodenum|Anatomy|false|false|C0496869;C0153426;C0002959|duodenumnull|biopsy characteristics|Finding|false|false||biopsy
null|null|Finding|false|false||biopsynull|Biopsy Procedures on the Pharynx, Adenoids, and Tonsils|Procedure|false|false||biopsy
null|Biopsy|Procedure|false|false||biopsy
null|Consent Type - biopsy|Procedure|false|false||biopsynull|biopsy characteristics|Finding|false|false||biopsy
null|null|Finding|false|false||biopsynull|Biopsy Procedures on the Pharynx, Adenoids, and Tonsils|Procedure|false|false||biopsy
null|Biopsy|Procedure|false|false||biopsy
null|Consent Type - biopsy|Procedure|false|false||biopsynull|Esophagogastroduodenoscopy|Procedure|false|false|C0013303|EGDnull|III (suffix)|Modifier|false|false||thirdnull|Third|LabModifier|false|false||thirdnull|part of|Modifier|false|false||part ofnull|Role Class - part|Finding|false|false|C0013303|partnull|Part|Modifier|false|false||partnull|Part Dosing Unit|LabModifier|false|false||partnull|Malignant neoplasm of duodenum|Disorder|false|false|C0013303|duodenum
null|Benign neoplasm of duodenum|Disorder|false|false|C0013303|duodenumnull|Duodenum|Anatomy|false|false|C0496869;C0153426;C1552020;C0079304|duodenumnull|Recommendation|Finding|false|false||Recommendationsnull|Obvious|Modifier|false|false||obviousnull|anatomic|Modifier|false|false||anatomicnull|Science of Etiology|Finding|false|false||cause
null|Etiology aspects|Finding|false|false||causenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Follow-up status|Finding|false|false||follow-upnull|follow-up|Procedure|false|false||follow-upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|biopsy characteristics|Finding|false|false||biopsy
null|null|Finding|false|false||biopsynull|Biopsy Procedures on the Pharynx, Adenoids, and Tonsils|Procedure|false|false||biopsy
null|Biopsy|Procedure|false|false||biopsy
null|Consent Type - biopsy|Procedure|false|false||biopsynull|Eosinophilic esophagitis|Disorder|false|false||eosinophilic esophagitisnull|Eosinophilic infiltration of the esophagus|Finding|false|false||eosinophilic esophagitisnull|eosinophilic|Finding|false|false||eosinophilicnull|Esophagitis|Disorder|false|false||esophagitisnull|Follow-up status|Finding|false|false||follow-upnull|follow-up|Procedure|false|false||follow-upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|Biopsy|Procedure|false|false||biopsiesnull|eosinophilic|Finding|false|false||eosinophilicnull|Esophagitis|Disorder|false|false||esophagitisnull|BRIEF Health Literacy Screening Tool|Finding|false|false||Brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||Briefnull|Brief|Time|false|false||Briefnull|Shortened|Modifier|false|false||Briefnull|Hospital course|Finding|false|false||Hospital Coursenull|null|Attribute|false|false||Hospital Coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||Coursenull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Gastroesophageal reflux disease|Disorder|false|false||GERDnull|Subacute|Time|false|false||subacutenull|Patient Outcome - Worsening|Finding|false|false||worseningnull|Worsening (qualifier value)|Modifier|false|false||worseningnull|Deglutition Disorders|Disorder|false|false||dysphagianull|Foreign body sensation (finding)|Finding|false|false|C0460148;C0444584;C4082212;C1268086;C0152338|foreign body sensation
null|Foreign body sensation in eyes|Finding|false|false|C0460148;C0444584;C4082212;C1268086;C0152338|foreign body sensationnull|Foreign Bodies|Disorder|false|false|C0460148;C0444584;C4082212;C1268086;C0152338|foreign bodynull|Foreign body (physical object)|Entity|false|false||foreign bodynull|International Aspects|Finding|false|false||foreignnull|foreign|Modifier|false|false||foreignnull|Document Body|Finding|false|false|C0460148;C0444584;C4082212;C1268086;C0152338|bodynull|Structure of body of caudate nucleus|Anatomy|false|false|C1551342;C0036658;C0542538;C2229507;C0920171;C0423602;C0016542|body
null|Human body structure|Anatomy|false|false|C1551342;C0036658;C0542538;C2229507;C0920171;C0423602;C0016542|body
null|Body structure|Anatomy|false|false|C1551342;C0036658;C0542538;C2229507;C0920171;C0423602;C0016542|body
null|Adult human body|Anatomy|false|false|C1551342;C0036658;C0542538;C2229507;C0920171;C0423602;C0016542|body
null|Whole body|Anatomy|false|false|C1551342;C0036658;C0542538;C2229507;C0920171;C0423602;C0016542|bodynull|Human body|Subject|false|false||bodynull|Observation of Sensation|Finding|false|false|C0460148;C0444584;C4082212;C1268086;C0152338|sensation
null|Sensory perception|Finding|false|false|C0460148;C0444584;C4082212;C1268086;C0152338|sensationnull|sensory exam|Procedure|false|false|C0460148;C0444584;C4082212;C1268086;C0152338|sensationnull|Sensation quality|Modifier|false|false||sensationnull|Point|Modifier|false|false||pointnull|point - UnitsOfMeasure|LabModifier|false|false||pointnull|Pureed|Modifier|false|false||pureednull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Last|Modifier|false|false||lastnull|10 days|Time|false|false||10 daysnull|day|Time|false|false||daysnull|Plain chest X-ray|Procedure|false|false||CXRnull|Prominent|Modifier|false|false||prominentnull|Carcinoma in situ of esophagus|Disorder|false|false|C4266613;C0014876|esophagus
null|Esophageal Diseases|Disorder|false|false|C4266613;C0014876|esophagus
null|Benign neoplasm of esophagus|Disorder|false|false|C4266613;C0014876|esophagusnull|Esophagus problem|Finding|false|false|C4266613;C0014876|esophagusnull|Procedures on the esophagus|Procedure|false|false|C4266613;C0014876|esophagusnull|Chest>Esophagus|Anatomy|false|false|C0014852;C0154059;C0153942;C0872395;C0812418|esophagus
null|Esophagus|Anatomy|false|false|C0014852;C0154059;C0153942;C0872395;C0812418|esophagusnull|Gastrointestinal studies and measurements|Finding|false|false||Gastroenterologynull|gastroenterology (field)|Title|false|false||Gastroenterologynull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Endoscopy, Gastrointestinal|Procedure|false|false||endoscopy
null|Endoscopy (procedure)|Procedure|false|false||endoscopynull|Carcinoma in situ of esophagus|Disorder|false|false|C4266613;C0014876|esophagus
null|Esophageal Diseases|Disorder|false|false|C4266613;C0014876|esophagus
null|Benign neoplasm of esophagus|Disorder|false|false|C4266613;C0014876|esophagusnull|Esophagus problem|Finding|false|false|C4266613;C0014876|esophagusnull|Procedures on the esophagus|Procedure|false|false|C4266613;C0014876|esophagusnull|Chest>Esophagus|Anatomy|false|false|C0014852;C0154059;C0153942;C0812418;C0872395|esophagus
null|Esophagus|Anatomy|false|false|C0014852;C0154059;C0153942;C0812418;C0872395|esophagusnull|Biopsy|Procedure|false|false||Biopsiesnull|Marketing basis - Transitional|Finding|false|false||TRANSITIONALnull|Transitional cell morphology|Modifier|false|false||TRANSITIONALnull|Biopsy|Procedure|false|false||biopsiesnull|Esophagogastroduodenoscopy|Procedure|false|false||EGDnull|Eosinophilic esophagitis|Disorder|false|false||eosinophilic esophagitisnull|Eosinophilic infiltration of the esophagus|Finding|false|false||eosinophilic esophagitisnull|eosinophilic|Finding|false|false||eosinophilicnull|Esophagitis|Disorder|false|false||esophagitisnull|Disease Management|Procedure|false|false||managementnull|Management Occupations|Subject|false|false||managementnull|Management procedure|Event|false|false||management
null|Administration occupational activities|Event|false|false||managementnull|Barium swallow|Procedure|false|false||barium swallownull|barium|Drug|false|false||bariumnull|Swallow - dosing instruction imperative|Finding|false|false||swallow
null|Swallow (administration method)|Finding|false|false||swallownull|Family Hirundinidae|Entity|false|false||swallownull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Further|Modifier|false|false||furthernull|Deglutition Disorders|Disorder|false|false||dysphagianull|ENT problem|Finding|false|false|C0150934;C0175196|ENT
null|NT5E gene|Finding|false|false|C0150934;C0175196|ENT
null|NT5E wt Allele|Finding|false|false|C0150934;C0175196|ENTnull|Structure of entorhinal cortex|Anatomy|false|false|C0262471;C3889152;C1417861|ENT
null|Ear, nose and throat|Anatomy|false|false|C0262471;C3889152;C1417861|ENTnull|Otolaryngology specialty|Title|false|false||ENTnull|MDF Attribute Type - Code|Finding|false|false||Code
null|A Codes|Finding|false|false||Code
null|Code|Finding|false|false||Codenull|Coding|Event|false|false||Codenull|Full|Modifier|false|false||Fullnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Accurate (qualifier value)|Modifier|false|false||accuratenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|omeprazole|Drug|false|false||Omeprazole
null|omeprazole|Drug|false|false||Omeprazolenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|omeprazole|Drug|false|false||Omeprazole
null|omeprazole|Drug|false|false||Omeprazolenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|null|Attribute|false|false||PRIMARY DIAGNOSISnull|Principal diagnosis|Modifier|false|false||PRIMARY DIAGNOSISnull|True primary (qualifier value)|Time|false|false||PRIMARYnull|Primary|Modifier|false|false||PRIMARYnull|Diagnosis Classification - Diagnosis|Finding|false|false||DIAGNOSIS
null|diagnosis aspects|Finding|false|false||DIAGNOSISnull|Diagnosis|Procedure|false|false||DIAGNOSISnull|null|Attribute|false|false||DIAGNOSISnull|Deglutition Disorders|Disorder|false|false||dysphagianull|Foreign body sensation (finding)|Finding|false|false|C0460148;C0444584;C4082212;C1268086;C0152338|foreign body sensation
null|Foreign body sensation in eyes|Finding|false|false|C0460148;C0444584;C4082212;C1268086;C0152338|foreign body sensationnull|Foreign Bodies|Disorder|false|false|C0460148;C0444584;C4082212;C1268086;C0152338|foreign bodynull|Foreign body (physical object)|Entity|false|false||foreign bodynull|International Aspects|Finding|false|false|C0460148;C0444584;C4082212;C1268086;C0152338|foreignnull|foreign|Modifier|false|false||foreignnull|Document Body|Finding|false|false|C0460148;C0444584;C4082212;C1268086;C0152338|bodynull|Structure of body of caudate nucleus|Anatomy|false|false|C0376327;C0016542;C0920171;C0423602;C1551342;C2229507|body
null|Human body structure|Anatomy|false|false|C0376327;C0016542;C0920171;C0423602;C1551342;C2229507|body
null|Body structure|Anatomy|false|false|C0376327;C0016542;C0920171;C0423602;C1551342;C2229507|body
null|Adult human body|Anatomy|false|false|C0376327;C0016542;C0920171;C0423602;C1551342;C2229507|body
null|Whole body|Anatomy|false|false|C0376327;C0016542;C0920171;C0423602;C1551342;C2229507|bodynull|Human body|Subject|false|false||bodynull|Observation of Sensation|Finding|false|false||sensation
null|Sensory perception|Finding|false|false||sensationnull|sensory exam|Procedure|false|false|C0460148;C0444584;C4082212;C1268086;C0152338|sensationnull|Sensation quality|Modifier|false|false||sensationnull|Secondary diagnosis|Finding|false|false||SECONDARY DIAGNOSISnull|null|Attribute|false|false||SECONDARY DIAGNOSISnull|Neoplasm Metastasis|Disorder|false|false||SECONDARYnull|metastatic qualifier|Finding|false|false||SECONDARYnull|Secondary to|Modifier|false|false||SECONDARYnull|second (number)|LabModifier|false|false||SECONDARYnull|Diagnosis Classification - Diagnosis|Finding|false|false||DIAGNOSIS
null|diagnosis aspects|Finding|false|false||DIAGNOSISnull|Diagnosis|Procedure|false|false||DIAGNOSISnull|null|Attribute|false|false||DIAGNOSISnull|Gastroesophageal reflux disease|Disorder|false|false||GERDnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Disease|Disorder|false|false||Conditionnull|Logical Condition|Finding|false|false||Conditionnull|null|Attribute|false|false||Conditionnull|Condition|Modifier|false|false||Conditionnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|Discharge instructions|Finding|false|false||Discharge Instructionsnull|hospital discharge instructions (treatment)|Procedure|false|false||Discharge Instructionsnull|null|Attribute|false|false||Discharge Instructionsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|FBXW7-AS1 gene|Finding|false|false||Dearnull|Has difficulty doing (qualifier value)|Finding|false|false||difficultynull|Endoscopy, Gastrointestinal|Procedure|false|false||endoscopy
null|Endoscopy (procedure)|Procedure|false|false||endoscopynull|Congenital Abnormality|Disorder|false|false|C4266613;C0014876|abnormalitiesnull|teratologic|Finding|false|false|C4266613;C0014876|abnormalitiesnull|Carcinoma in situ of esophagus|Disorder|false|false|C4266613;C0014876|esophagus
null|Esophageal Diseases|Disorder|false|false|C4266613;C0014876|esophagus
null|Benign neoplasm of esophagus|Disorder|false|false|C4266613;C0014876|esophagusnull|Esophagus problem|Finding|false|false|C4266613;C0014876|esophagusnull|Procedures on the esophagus|Procedure|false|false|C4266613;C0014876|esophagusnull|Chest>Esophagus|Anatomy|false|false|C0872395;C0812418;C0014852;C0154059;C0153942;C0000768;C0000769|esophagus
null|Esophagus|Anatomy|false|false|C0872395;C0812418;C0014852;C0154059;C0153942;C0000768;C0000769|esophagusnull|Biopsy|Procedure|false|false||biopsiesnull|Tests (qualifier value)|Finding|false|false|C4318744|test
null|Testing|Finding|false|false|C4318744|testnull|Laboratory Procedures|Procedure|false|false|C4318744|testnull|Test - temporal region|Anatomy|false|false|C0022885;C0004749;C0203065;C0456984;C4521686;C1706486;C0039593;C0392366|testnull|Test Result|Lab|false|false|C4318744|testnull|Test Dosing Unit|LabModifier|false|false||testnull|Barium swallow|Procedure|false|false|C4318744|barium swallownull|barium|Drug|false|false|C4318744|bariumnull|Swallow - dosing instruction imperative|Finding|false|false|C4318744|swallow
null|Swallow (administration method)|Finding|false|false|C4318744|swallownull|Family Hirundinidae|Entity|false|false||swallownull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Vitelliform Macular Dystrophy|Disorder|false|false||bestnull|BEST1 wt Allele|Finding|false|false||best
null|BEST1 gene|Finding|false|false||bestnull|best (quality)|Modifier|false|false||bestnull|Team|Subject|false|false||Teamnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions