﻿Numbered||(?:^[\t ]*[\d]{1,2}(?::|\.)[\t ]+(?:(?!^[ ]*[\d]{1,2}(?::|\.)[\t ]+)(?:[^\t\r\n]+\r?\n))+){2,}||^[\t ]*[\d]{1,2}(?::|\.)[\t ]+(?:(?!^[\t ]*[\d]{1,2}(?::|\.)[\t ]+)(?:[^\t\r\n]+\r?\n))+
Alpha Sentence||(?:^[\t ]*[A-Z](?::|\.)+\)?[\t ]+(?:[^\t\n\.]+(?:\.|\n))+\r?\n){2,}||^[\t ]*[A-Z](?::|\.)+\)?[\t ]+(?:[^\t\n\.]+(?:\.|\n))+\r?\n
// Name Value||(?:^[^\t\r\n]{2,50}:[\t ]+(?:[^\t\r\n:]+\r?\n)+){3,}||^[^\t\r\n]{2,50}:[\t ]+(?:[^\t\r\n:]+\r?\n)+
Name Value||(?:^[^\r\n:]{2,}:[\s]+[^\r\n]+\r?\n){2,}||^[^\r\n:]{2,80}:[\s]+[^\r\n]+\r?\n
// Multi Column||(?:^(?:[^\s:]+(?: [^\s:]+)*(?:\t+| {3,}))+(?:[^\s]+(?: [^\s]+)*)[\t ]*\r?\n){3,}||\r?\n
// Mixed Column||(?:^(?:[^\s:]+(?: [^\s:]+)*(?:\t+| {3,}))+(?:[^\s]+(?: [^\s]+)*)[\t ]*\r?\n[\t ]*(?:[^\s]+(?: [^\s]+)*)[\t ]*\r?\n){3,}||[\r\n][\t ]*(?:[^\s]+(?: [^\s]+)*)[\t ]*\r?\n
// Header||(?:^[^\t\r\n\.]+\.{3,}[^\t\r\n\.]+\r?\n){3,}||\r?\n
Dash||(?:^[\t ]*-{1,3}[\t ]+(?:(?:[^\t\r\n-]+-?)+\r?\n){1,3}){2,}||^[\t ]*-{1,3}[\t ]+(?:(?:[^\t\r\n-]+-?)+\r?\n)+
// Document Header||(?:^[^\t\r\n\.]+\.{3,}[^\t\r\n\.]+\r?\n){3,}||\r?\n
Checkbox||(?:^(?:[^\r\n:]{2,80}:\r?\n)?(?:[\t ]*\[[XYN _]*\][^\r\n]+\r?\n)+)+||^(?:[^\r\n:]{2,80}:\r?\n)?(?:[\t ]*\[[XYN _]*\][^\r\n]+\r?\n)+
// Name Colon Value||(?:^[\t ]*[^\t\r\n:]+:[^\t\r\n:]+\r?\n){2,}||^[\t ]*[^\t\r\n:]+:[^\t\r\n:]+\r?\n
