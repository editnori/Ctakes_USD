 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|48,57|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|48,57|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|48,62|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|82,91|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|82,91|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|82,91|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|82,91|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|82,91|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|82,96|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|114,119|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|114,119|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|114,119|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|138,141|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|138,141|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|138,141|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|138,141|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|138,141|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|149,156|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|149,156|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|SIMPLE_SEGMENT|158,170|true|false|false|||NEUROSURGERY
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|158,170|true|false|false|C0524850|Neurosurgical Procedures|NEUROSURGERY
Attribute|Clinical Attribute|Allergies|194,203|true|false|false|C1717415||Allergies
Event|Event|Allergies|194,203|true|false|false|||Allergies
Finding|Pathologic Function|Allergies|194,203|true|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|Allergies|206,228|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|Allergies|214,218|true|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|Allergies|214,218|true|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|Allergies|214,228|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Event|Event|Allergies|219,228|true|false|false|||Reactions
Event|Event|Allergies|231,240|false|false|false|||Attending
Finding|Functional Concept|Allergies|231,240|false|false|false|C1999232|Attending (action)|Attending
Event|Event|Chief Complaint|266,275|false|false|false|||Headaches
Finding|Sign or Symptom|Chief Complaint|266,275|false|false|false|C0018681|Headache|Headaches
Finding|Classification|Chief Complaint|278,283|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|284,292|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|284,292|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|296,314|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|305,314|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|305,314|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|305,314|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|305,314|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|305,314|false|false|false|C0184661|Interventional procedure|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|322,345|false|false|false|C2066670|suboccipital craniotomy|Suboccipital craniotomy
Event|Event|Chief Complaint|335,345|false|false|false|||craniotomy
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|335,345|false|false|false|C0010280|Craniotomy|craniotomy
Event|Event|Chief Complaint|350,359|false|false|false|||resection
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|350,359|false|false|false|C0015252;C0728940|Excision;removal technique|resection
Anatomy|Body Part, Organ, or Organ Component|Chief Complaint|363,373|false|false|false|C0007765|Cerebellum|cerebellar
Event|Event|Chief Complaint|375,381|false|false|false|||lesion
Finding|Finding|Chief Complaint|375,381|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|Chief Complaint|375,381|false|false|false|C0221198;C1546698|Lesion|lesion
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|441,449|false|false|false|C0006104;C0228174|Brain;Cerebral hemisphere structure (body structure)|cerebral
Disorder|Disease or Syndrome|History of Present Illness|441,458|false|false|false|C0917996|Cerebral Aneurysm|cerebral aneurysm
Event|Event|History of Present Illness|450,458|false|false|false|||aneurysm
Finding|Pathologic Function|History of Present Illness|450,458|false|false|false|C0002940|Aneurysm|aneurysm
Event|Event|History of Present Illness|460,468|false|false|false|||clipping
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|460,468|false|false|false|C0185010|Closure by clip (procedure)|clipping
Event|Event|History of Present Illness|480,488|false|false|false|||presents
Event|Event|History of Present Illness|494,497|false|false|false|||OSH
Finding|Functional Concept|History of Present Illness|503,507|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|508,518|false|false|false|C0007765|Cerebellum|cerebellar
Event|Event|History of Present Illness|520,531|false|false|false|||hypodensity
Event|Event|History of Present Illness|558,564|false|false|false|||lesion
Finding|Finding|History of Present Illness|558,564|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|History of Present Illness|558,564|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Body Substance|History of Present Illness|566,573|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|566,573|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|566,573|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|566,581|false|false|false|C0747307|Patient-Reported|Patient reports
Event|Event|History of Present Illness|574,581|false|false|false|||reports
Finding|Intellectual Product|History of Present Illness|574,581|false|false|false|C0684224|Report (document)|reports
Procedure|Health Care Activity|History of Present Illness|574,581|false|false|false|C0700287|Reporting|reports
Finding|Gene or Genome|History of Present Illness|600,603|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|History of Present Illness|608,615|false|false|false|||started
Event|Event|History of Present Illness|623,632|false|false|false|||headaches
Finding|Sign or Symptom|History of Present Illness|623,632|false|false|false|C0018681|Headache|headaches
Event|Event|History of Present Illness|644,652|false|false|false|||abnormal
Finding|Finding|History of Present Illness|644,652|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Finding|Idea or Concept|History of Present Illness|644,652|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Event|Event|History of Present Illness|666,675|false|false|false|||describes
Event|Event|History of Present Illness|680,689|false|false|false|||headaches
Finding|Sign or Symptom|History of Present Illness|680,689|false|false|false|C0018681|Headache|headaches
Event|Event|History of Present Illness|708,715|false|false|false|||resolve
Drug|Organic Chemical|History of Present Illness|721,728|false|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|History of Present Illness|721,728|false|false|false|C0699142|Tylenol|Tylenol
Event|Event|History of Present Illness|769,776|false|false|false|||reports
Event|Event|History of Present Illness|784,794|false|false|false|||difficulty
Finding|Finding|History of Present Illness|784,794|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Finding|Finding|History of Present Illness|784,802|false|false|false|C0311394|Difficulty walking|difficulty walking
Event|Event|History of Present Illness|795,802|false|false|false|||walking
Finding|Daily or Recreational Activity|History of Present Illness|795,802|false|false|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Finding|Finding|History of Present Illness|795,802|false|false|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Finding|Sign or Symptom|History of Present Illness|795,802|false|false|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Event|Event|History of Present Illness|815,822|false|false|false|||started
Finding|Gene or Genome|History of Present Illness|842,845|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|History of Present Illness|851,860|false|false|false|||describes
Event|Event|History of Present Illness|865,872|false|false|false|||walking
Finding|Daily or Recreational Activity|History of Present Illness|865,872|false|false|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Finding|Finding|History of Present Illness|865,872|false|false|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Finding|Sign or Symptom|History of Present Illness|865,872|false|false|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Disorder|Disease or Syndrome|History of Present Illness|877,887|false|false|false|C0344191|Cerebellar decompression injury|staggering
Finding|Sign or Symptom|History of Present Illness|877,887|false|false|false|C0701824|Staggering gait|staggering
Finding|Finding|History of Present Illness|894,901|false|false|false|C0516750|side to side|to side
Event|Event|History of Present Illness|908,914|true|false|false|||denies
Attribute|Clinical Attribute|History of Present Illness|919,925|true|false|false|C2707266||vision
Finding|Organism Function|History of Present Illness|919,925|true|false|false|C0042789|Vision|vision
Event|Event|History of Present Illness|926,933|true|false|false|||changes
Finding|Functional Concept|History of Present Illness|926,933|true|false|false|C0392747|Changing|changes
Attribute|Clinical Attribute|History of Present Illness|935,941|true|false|false|C4255480||nausea
Event|Event|History of Present Illness|935,941|true|false|false|||nausea
Finding|Sign or Symptom|History of Present Illness|935,941|true|false|false|C0027497|Nausea|nausea
Event|Event|History of Present Illness|943,951|true|false|false|||vomiting
Finding|Sign or Symptom|History of Present Illness|943,951|true|false|false|C0042963|Vomiting|vomiting
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|954,963|false|false|false|C0009676|Confusion|confusion
Event|Event|History of Present Illness|954,963|false|false|false|||confusion
Finding|Finding|History of Present Illness|954,963|false|false|false|C0683369|Clouded consciousness|confusion
Finding|Idea or Concept|History of Present Illness|968,972|false|false|false|C1705313|Term (lexical)|word
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|968,991|false|false|false|C0454643|Word finding difficulty (disorder)|word finding difficulty
Finding|Finding|History of Present Illness|973,980|false|false|false|C0037088;C0243095;C2825141|Experimental Finding;Finding;Signs and Symptoms|finding
Finding|Sign or Symptom|History of Present Illness|973,980|false|false|false|C0037088;C0243095;C2825141|Experimental Finding;Finding;Signs and Symptoms|finding
Event|Event|History of Present Illness|981,991|false|false|false|||difficulty
Finding|Finding|History of Present Illness|981,991|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Event|Event|History of Present Illness|997,1000|false|false|false|||saw
Anatomy|Body Location or Region|History of Present Illness|1005,1008|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1005,1008|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Disorder|Disease or Syndrome|History of Present Illness|1005,1008|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Disorder|Neoplastic Process|History of Present Illness|1005,1008|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Finding|Body Substance|History of Present Illness|1005,1008|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Finding|History of Present Illness|1005,1008|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Intellectual Product|History of Present Illness|1005,1008|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Event|Event|History of Present Illness|1009,1015|false|false|false|||doctor
Finding|Intellectual Product|History of Present Illness|1009,1015|false|false|false|C2348314|Doctor - Title|doctor
Finding|Idea or Concept|History of Present Illness|1034,1041|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|routine
Finding|Intellectual Product|History of Present Illness|1034,1041|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|routine
Procedure|Laboratory Procedure|History of Present Illness|1034,1041|false|false|false|C1979801|Routine coag|routine
Event|Event|History of Present Illness|1042,1047|false|false|false|||visit
Finding|Social Behavior|History of Present Illness|1042,1047|false|false|false|C0545082|Visit|visit
Event|Event|History of Present Illness|1053,1061|false|false|false|||referred
Event|Event|History of Present Illness|1081,1091|false|false|false|||evaluation
Finding|Idea or Concept|History of Present Illness|1081,1091|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|History of Present Illness|1081,1091|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Event|Event|History of Present Illness|1101,1109|false|false|false|||symptoms
Finding|Functional Concept|History of Present Illness|1101,1109|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|History of Present Illness|1101,1109|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|History of Present Illness|1118,1124|false|false|false|||showed
Event|Event|History of Present Illness|1128,1132|false|false|false|||area
Event|Governmental or Regulatory Activity|History of Present Illness|1128,1132|false|false|false|C1510751|Academic Research Enhancement Awards|area
Event|Event|History of Present Illness|1137,1148|false|false|false|||hypodensity
Finding|Functional Concept|History of Present Illness|1156,1160|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1161,1171|false|false|false|C0007765|Cerebellum|cerebellum
Disorder|Neoplastic Process|History of Present Illness|1161,1171|false|false|false|C0153640|Malignant neoplasm of cerebellum|cerebellum
Event|Event|History of Present Illness|1188,1198|false|false|false|||underlying
Finding|Finding|History of Present Illness|1188,1198|false|false|false|C4722602|Underlying|underlying
Event|Event|History of Present Illness|1200,1206|false|false|false|||lesion
Finding|Finding|History of Present Illness|1200,1206|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|History of Present Illness|1200,1206|false|false|false|C0221198;C1546698|Lesion|lesion
Event|Event|History of Present Illness|1229,1240|false|false|false|||transferred
Finding|Body Substance|History of Present Illness|1260,1267|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1260,1267|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1260,1267|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|1268,1275|true|false|false|||reports
Finding|Pathologic Function|History of Present Illness|1280,1288|true|false|false|C0002940|Aneurysm|aneurysm
Event|Event|History of Present Illness|1289,1293|true|false|false|||clip
Finding|Gene or Genome|History of Present Illness|1289,1293|true|false|false|C1337111;C1413237;C1561603;C1704793;C1824746;C1824747;C2827463|CD74 gene;CLIP - Codes for radiology reports;CLIP1 gene;CLIP1 wt Allele;CLIP2 gene;POMC gene;POMC wt Allele|clip
Finding|Intellectual Product|History of Present Illness|1289,1293|true|false|false|C1337111;C1413237;C1561603;C1704793;C1824746;C1824747;C2827463|CD74 gene;CLIP - Codes for radiology reports;CLIP1 gene;CLIP1 wt Allele;CLIP2 gene;POMC gene;POMC wt Allele|clip
Procedure|Health Care Activity|History of Present Illness|1289,1293|true|false|false|C5552742|Comprehensive Lifestyle Intervention Program|clip
Event|Event|History of Present Illness|1301,1304|true|false|false|||MRI
Finding|Gene or Genome|History of Present Illness|1301,1304|true|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|History of Present Illness|1301,1304|true|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|History of Present Illness|1301,1304|true|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Event|Event|History of Present Illness|1306,1316|true|false|false|||compatible
Finding|Idea or Concept|History of Present Illness|1306,1316|true|false|false|C0332290|Consistent with|compatible
Disorder|Disease or Syndrome|Past Medical History|1352,1364|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|Past Medical History|1352,1364|false|false|false|||Hypertension
Finding|Pathologic Function|Past Medical History|1372,1380|false|false|false|C0002940|Aneurysm|aneurysm
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1372,1389|false|false|false|C0189711|Clipping arterial aneurysm|aneurysm clipping
Event|Event|Past Medical History|1381,1389|false|false|false|||clipping
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1381,1389|false|false|false|C0185010|Closure by clip (procedure)|clipping
Event|Event|Family Medical History|1459,1466|true|false|false|||history
Finding|Conceptual Entity|Family Medical History|1459,1466|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|1459,1466|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Family Medical History|1459,1466|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|1459,1469|true|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|Family Medical History|1470,1476|true|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|Family Medical History|1470,1476|true|false|false|||stroke
Finding|Finding|Family Medical History|1470,1476|true|false|false|C5977286|Stroke (heart beat)|stroke
Disorder|Neoplastic Process|Family Medical History|1478,1484|true|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Family Medical History|1478,1484|true|false|false|||cancer
Event|Event|Family Medical History|1486,1494|false|false|false|||aneurysm
Finding|Pathologic Function|Family Medical History|1486,1494|true|false|false|C0002940|Aneurysm|aneurysm
Procedure|Health Care Activity|General Exam|1518,1527|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|General Exam|1588,1591|false|false|false|||Gen
Finding|Classification|General Exam|1588,1591|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Finding|Gene or Genome|General Exam|1588,1591|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Event|Event|General Exam|1600,1611|false|false|false|||comfortable
Finding|Finding|General Exam|1600,1611|false|false|false|C5546696|Feeling comfortable|comfortable
Disorder|Disease or Syndrome|General Exam|1613,1616|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|1613,1616|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|1613,1616|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|1613,1616|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|1613,1616|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|General Exam|1613,1616|false|false|false|||NAD
Finding|Finding|General Exam|1613,1616|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|General Exam|1618,1623|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|General Exam|1625,1631|false|false|false|C0034121|Pupil|Pupils
Finding|Functional Concept|General Exam|1653,1657|false|false|false|C0241886|Extraocular|EOMs
Anatomy|Body Location or Region|General Exam|1663,1667|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|General Exam|1663,1667|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|General Exam|1663,1667|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|General Exam|1669,1675|false|false|false|||Supple
Finding|Functional Concept|General Exam|1669,1675|false|false|false|C0332254|Supple|Supple
Event|Event|General Exam|1685,1689|false|false|false|||Warm
Finding|Finding|General Exam|1685,1689|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|1685,1689|false|false|false|C0687712|warming process|Warm
Finding|Finding|General Exam|1694,1698|false|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|1699,1707|false|false|false|||perfused
Finding|Mental Process|General Exam|1717,1723|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|General Exam|1717,1730|false|false|false|C0488568;C0488569||Mental status
Finding|Finding|General Exam|1717,1730|false|false|false|C0278060|Mental state|Mental status
Attribute|Clinical Attribute|General Exam|1724,1730|false|false|false|C5889824||status
Event|Event|General Exam|1724,1730|false|false|false|||status
Finding|Idea or Concept|General Exam|1724,1730|false|false|false|C1546481|What subject filter - Status|status
Event|Event|General Exam|1732,1737|false|false|false|||Awake
Attribute|Clinical Attribute|General Exam|1742,1747|false|false|false|C5890168||alert
Drug|Organic Chemical|General Exam|1742,1747|false|false|false|C0718338|Alert brand of caffeine|alert
Drug|Pharmacologic Substance|General Exam|1742,1747|false|false|false|C0718338|Alert brand of caffeine|alert
Event|Event|General Exam|1742,1747|false|false|false|||alert
Finding|Finding|General Exam|1742,1747|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Functional Concept|General Exam|1742,1747|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Intellectual Product|General Exam|1742,1747|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Event|Event|General Exam|1749,1760|false|false|false|||cooperative
Event|Event|General Exam|1766,1770|false|false|false|||exam
Finding|Functional Concept|General Exam|1766,1770|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|General Exam|1766,1770|false|false|false|C0582103|Medical Examination|exam
Event|Event|General Exam|1772,1778|false|false|false|||normal
Event|Event|General Exam|1779,1785|false|false|false|||affect
Finding|Mental Process|General Exam|1779,1785|false|false|false|C0001721|Affect (mental function)|affect
Procedure|Health Care Activity|General Exam|1779,1785|false|false|false|C2237113|assessment of affect|affect
Event|Event|General Exam|1787,1798|false|false|false|||Orientation
Finding|Mental Process|General Exam|1787,1798|false|false|false|C0029266|Mental Orientation|Orientation
Event|Event|General Exam|1800,1808|false|false|false|||Oriented
Finding|Finding|General Exam|1800,1808|false|false|false|C1961028|Oriented to place|Oriented
Finding|Finding|General Exam|1800,1818|false|false|false|C1961030|Oriented to person|Oriented to person
Attribute|Clinical Attribute|General Exam|1812,1818|false|false|false|C5890614||person
Event|Event|General Exam|1812,1818|false|false|false|||person
Finding|Intellectual Product|General Exam|1812,1818|false|false|false|C1522390|Person Info|person
Event|Activity|General Exam|1820,1825|false|false|false|C1882509|put - instruction imperative|place
Event|Event|General Exam|1820,1825|false|false|false|||place
Finding|Functional Concept|General Exam|1820,1825|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|General Exam|1820,1825|false|false|false|C1533810||place
Attribute|Clinical Attribute|General Exam|1837,1845|false|false|false|C2706915||Language
Event|Event|General Exam|1837,1845|false|false|false|||Language
Finding|Intellectual Product|General Exam|1837,1845|false|false|false|C0033348|Programming Languages|Language
Event|Event|General Exam|1847,1853|false|false|false|||Speech
Finding|Organism Function|General Exam|1847,1853|false|false|false|C0037817|Speech|Speech
Procedure|Diagnostic Procedure|General Exam|1847,1853|false|false|false|C0846595|Speech assessment|Speech
Finding|Idea or Concept|General Exam|1866,1870|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Event|Event|General Exam|1871,1884|false|false|false|||comprehension
Finding|Mental Process|General Exam|1871,1884|false|false|false|C0162340|Comprehension|comprehension
Event|Event|General Exam|1889,1899|false|false|false|||repetition
Finding|Finding|General Exam|1889,1899|false|false|false|C0205341;C2018025|Repeat;speech fluency repetition (physical finding)|repetition
Finding|Functional Concept|General Exam|1889,1899|false|false|false|C0205341;C2018025|Repeat;speech fluency repetition (physical finding)|repetition
Event|Event|General Exam|1901,1907|false|false|false|||Naming
Finding|Mental Process|General Exam|1901,1907|false|false|false|C0233735|Naming (function)|Naming
Event|Event|General Exam|1908,1914|false|false|false|||intact
Finding|Finding|General Exam|1908,1914|false|false|false|C1554187|Gender Status - Intact|intact
Disorder|Mental or Behavioral Dysfunction|General Exam|1919,1929|true|false|false|C0013362|Dysarthria|dysarthria
Event|Event|General Exam|1919,1929|true|false|false|||dysarthria
Event|Event|General Exam|1944,1950|true|false|false|||errors
Anatomy|Body Part, Organ, or Organ Component|General Exam|1953,1960|false|false|false|C0037303|Bone structure of cranium|Cranial
Anatomy|Body Part, Organ, or Organ Component|General Exam|1953,1967|false|false|false|C0010268|Cranial Nerves|Cranial Nerves
Disorder|Neoplastic Process|General Exam|1953,1967|false|false|false|C0004992;C0496937|Benign neoplasm of cranial nerves;Neoplasm of uncertain or unknown behavior of cranial nerves|Cranial Nerves
Anatomy|Body Part, Organ, or Organ Component|General Exam|1961,1967|false|false|false|C0027740|Nerve|Nerves
Event|Event|General Exam|1976,1982|true|false|false|||tested
Finding|Functional Concept|General Exam|1987,1991|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|General Exam|1987,1997|false|false|false|C0229187|Structure of pupil of left eye|Left pupil
Anatomy|Body Part, Organ, or Organ Component|General Exam|1992,1997|false|false|false|C0034121;C1305618|Pupil|pupil
Finding|Functional Concept|General Exam|2005,2010|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Event|Event|General Exam|2031,2039|false|false|false|||reactive
Procedure|Therapeutic or Preventive Procedure|General Exam|2031,2039|false|false|false|C4722408|Reactive Therapy|reactive
Drug|Amino Acid, Peptide, or Protein|General Exam|2043,2048|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|General Exam|2043,2048|false|false|false|C1570446|TNFSF14 protein, human|light
Event|Event|General Exam|2043,2048|false|false|false|||light
Finding|Finding|General Exam|2043,2048|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|General Exam|2043,2048|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|General Exam|2043,2048|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|General Exam|2043,2048|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|General Exam|2043,2048|false|false|false|C0031765|Phototherapy|light
Finding|Functional Concept|General Exam|2064,2075|true|false|false|C0241886|Extraocular|Extraocular
Procedure|Diagnostic Procedure|General Exam|2064,2085|true|false|false|C2228439|examination of extraocular movements|Extraocular movements
Event|Event|General Exam|2076,2085|true|false|false|||movements
Finding|Organism Function|General Exam|2076,2085|true|false|false|C0026649|Movement|movements
Event|Event|General Exam|2086,2092|true|false|false|||intact
Finding|Finding|General Exam|2086,2092|true|false|false|C1554187|Gender Status - Intact|intact
Disorder|Disease or Syndrome|General Exam|2113,2122|true|false|false|C0028738|Nystagmus|nystagmus
Event|Event|General Exam|2113,2122|true|false|false|||nystagmus
Anatomy|Body Part, Organ, or Organ Component|General Exam|2127,2130|false|false|false|C2338708;C3496273;C3496274|Lamina VII of gray matter of spinal cord;layer VII (Cajal);lobule VII|VII
Finding|Intellectual Product|General Exam|2127,2130|false|false|false|C0445385|Roman numeral VII|VII
Anatomy|Body Location or Region|General Exam|2132,2138|false|false|false|C0015450|Face|Facial
Event|Event|General Exam|2139,2147|false|false|false|||strength
Finding|Idea or Concept|General Exam|2139,2147|false|false|false|C0808080|Strength (attribute)|strength
Event|Event|General Exam|2152,2161|false|false|false|||sensation
Finding|Finding|General Exam|2152,2161|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|General Exam|2152,2161|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|General Exam|2152,2161|false|false|false|C2229507|sensory exam|sensation
Event|Event|General Exam|2162,2168|false|false|false|||intact
Finding|Finding|General Exam|2162,2168|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|General Exam|2173,2182|false|false|false|||symmetric
Finding|Conceptual Entity|General Exam|2173,2182|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|General Exam|2173,2182|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Anatomy|Body Part, Organ, or Organ Component|General Exam|2188,2207|false|false|false|C0224153|Structure of sternocleidomastoid muscle|Sternocleidomastoid
Anatomy|Body Part, Organ, or Organ Component|General Exam|2212,2221|false|false|false|C0224361|Structure of trapezius muscle|trapezius
Event|Event|General Exam|2222,2228|false|false|false|||normal
Anatomy|Body Part, Organ, or Organ Component|General Exam|2247,2253|true|false|false|C0040408|Tongue|Tongue
Disorder|Neoplastic Process|General Exam|2247,2253|true|false|false|C0153933|Benign neoplasm of tongue|Tongue
Procedure|Health Care Activity|General Exam|2247,2253|true|false|false|C0872394|Procedure on tongue|Tongue
Finding|Finding|General Exam|2247,2261|true|false|false|C3693372|tongue midline|Tongue midline
Anatomy|Cell Component|General Exam|2254,2261|true|false|false|C1660780|midline cell component|midline
Event|Event|General Exam|2270,2284|true|false|false|||fasciculations
Finding|Sign or Symptom|General Exam|2270,2284|true|false|false|C0015644|Muscular fasciculation|fasciculations
Event|Event|General Exam|2287,2292|false|false|false|||Motor
Finding|Functional Concept|General Exam|2287,2292|false|false|false|C1513492|motor movement|Motor
Drug|Biomedical or Dental Material|General Exam|2301,2305|false|false|false|C0012173;C1337615|Bulk (conceptual);Dietary Fiber|bulk
Drug|Food|General Exam|2301,2305|false|false|false|C0012173;C1337615|Bulk (conceptual);Dietary Fiber|bulk
Event|Event|General Exam|2301,2305|false|false|false|||bulk
Event|Event|General Exam|2310,2314|false|false|false|||tone
Finding|Finding|General Exam|2331,2339|true|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Finding|Idea or Concept|General Exam|2331,2339|true|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Disorder|Disease or Syndrome|General Exam|2331,2349|true|false|false|C0013384|Dyskinetic syndrome|abnormal movements
Finding|Finding|General Exam|2331,2349|true|false|false|C0558189|Abnormal movement|abnormal movements
Event|Event|General Exam|2340,2349|true|false|false|||movements
Finding|Organism Function|General Exam|2340,2349|true|false|false|C0026649|Movement|movements
Event|Event|General Exam|2351,2358|true|false|false|||tremors
Finding|Sign or Symptom|General Exam|2351,2358|true|false|false|C0040822|Tremor|tremors
Finding|Idea or Concept|General Exam|2360,2368|false|false|false|C0808080|Strength (attribute)|Strength
Finding|Social Behavior|General Exam|2374,2379|false|false|false|C0032863|Power (Psychology)|power
Finding|Finding|General Exam|2396,2402|false|false|false|C5202796|Intensity and Distress 1|Slight
Finding|Functional Concept|General Exam|2403,2407|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Event|Event|General Exam|2423,2432|false|false|false|||Sensation
Finding|Finding|General Exam|2423,2432|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Finding|Organ or Tissue Function|General Exam|2423,2432|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Procedure|Health Care Activity|General Exam|2423,2432|false|false|false|C2229507|sensory exam|Sensation
Event|Event|General Exam|2434,2440|false|false|false|||Intact
Finding|Finding|General Exam|2434,2440|false|false|false|C1554187|Gender Status - Intact|Intact
Drug|Amino Acid, Peptide, or Protein|General Exam|2444,2449|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|General Exam|2444,2449|false|false|false|C1570446|TNFSF14 protein, human|light
Event|Event|General Exam|2444,2449|false|false|false|||light
Finding|Finding|General Exam|2444,2449|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|General Exam|2444,2449|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|General Exam|2444,2449|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|General Exam|2444,2449|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|General Exam|2444,2449|false|false|false|C0031765|Phototherapy|light
Finding|Physiologic Function|General Exam|2444,2455|false|false|false|C0423553|Light touch|light touch
Event|Event|General Exam|2450,2455|false|false|false|||touch
Finding|Mental Process|General Exam|2450,2455|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Finding|Organ or Tissue Function|General Exam|2450,2455|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Procedure|Therapeutic or Preventive Procedure|General Exam|2450,2455|false|false|false|C0152054|Therapeutic Touch|touch
Event|Event|General Exam|2457,2469|false|false|false|||Coordination
Finding|Functional Concept|General Exam|2457,2469|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Finding|Idea or Concept|General Exam|2457,2469|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Finding|Physiologic Function|General Exam|2457,2469|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Event|Event|General Exam|2471,2477|false|false|false|||normal
Anatomy|Body Part, Organ, or Organ Component|General Exam|2481,2487|false|false|false|C0016129;C0851278;C4299059|Fingers;Fingers not including thumb;Upper extremity>Finger|finger
Anatomy|Body Part, Organ, or Organ Component|General Exam|2493,2499|false|false|false|C0016129;C0851278;C4299059|Fingers;Fingers not including thumb;Upper extremity>Finger|finger
Anatomy|Body Part, Organ, or Organ Component|General Exam|2504,2508|false|false|false|C0018870|Heel|heel
Anatomy|Body Location or Region|General Exam|2512,2516|false|false|false|C0230444|Shin|shin
Finding|Body Substance|General Exam|2577,2586|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|2577,2586|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|2577,2586|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|2577,2586|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|General Exam|2589,2593|false|false|false|||Exam
Finding|Functional Concept|General Exam|2589,2593|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|General Exam|2589,2593|false|false|false|C0582103|Medical Examination|Exam
Anatomy|Body Part, Organ, or Organ Component|General Exam|2602,2606|false|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|General Exam|2602,2606|false|false|false|C5848506||eyes
Event|Event|General Exam|2611,2622|false|false|false|||Spontaneous
Event|Event|General Exam|2650,2661|false|false|false|||Orientation
Finding|Mental Process|General Exam|2650,2661|false|false|false|C0029266|Mental Orientation|Orientation
Attribute|Clinical Attribute|General Exam|2666,2672|false|false|false|C5890614||Person
Finding|Intellectual Product|General Exam|2666,2672|false|false|false|C1522390|Person Info|Person
Event|Activity|General Exam|2676,2681|false|false|false|C1882509|put - instruction imperative|Place
Event|Event|General Exam|2676,2681|false|false|false|||Place
Finding|Functional Concept|General Exam|2676,2681|false|false|false|C1704765|Place - dosing instruction imperative|Place
Procedure|Health Care Activity|General Exam|2676,2681|false|false|false|C1533810||Place
Finding|Finding|General Exam|2685,2689|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Finding|Idea or Concept|General Exam|2685,2689|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Finding|Intellectual Product|General Exam|2685,2689|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Event|Event|General Exam|2699,2707|false|false|false|||commands
Finding|Gene or Genome|General Exam|2712,2718|true|false|false|C1424587|LITAF gene|Simple
Drug|Chemical Viewed Structurally|General Exam|2722,2729|true|false|false|C1704241|complex (molecular entity)|Complex
Anatomy|Body Part, Organ, or Organ Component|General Exam|2739,2745|true|false|false|C0034121|Pupil|Pupils
Finding|Functional Concept|General Exam|2748,2753|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Finding|Functional Concept|General Exam|2766,2770|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Event|Event|General Exam|2779,2786|false|false|false|||chronic
Finding|Intellectual Product|General Exam|2779,2786|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|General Exam|2779,2786|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Anatomy|Body Part, Organ, or Organ Component|General Exam|2788,2791|false|false|false|C0028863|Muscle of orbit|EOM
Finding|Functional Concept|General Exam|2788,2791|false|false|false|C0241886|Extraocular|EOM
Event|Event|General Exam|2817,2824|false|false|false|||chronic
Finding|Intellectual Product|General Exam|2817,2824|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|General Exam|2817,2824|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Finding|Functional Concept|General Exam|2841,2845|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|General Exam|2856,2860|false|false|false|C0015450;C4266571|Face;Head>Face|Face
Disorder|Disease or Syndrome|General Exam|2856,2860|false|false|false|C3160739|FANCONI ANEMIA, COMPLEMENTATION GROUP E|Face
Event|Event|General Exam|2856,2860|false|false|false|||Face
Finding|Gene or Genome|General Exam|2856,2860|false|false|false|C1414531;C1423759;C2828055|ELOVL6 gene;FANCE gene;FANCE wt Allele|Face
Finding|Conceptual Entity|General Exam|2861,2870|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|Symmetric
Finding|Finding|General Exam|2861,2870|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|Symmetric
Finding|Finding|General Exam|2875,2878|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Gene or Genome|General Exam|2875,2878|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Idea or Concept|General Exam|2875,2878|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Intellectual Product|General Exam|2875,2878|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Anatomy|Cell Component|General Exam|2891,2898|false|false|false|C1660780|midline cell component|Midline
Finding|Finding|General Exam|2903,2906|true|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Gene or Genome|General Exam|2903,2906|true|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Idea or Concept|General Exam|2903,2906|true|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Intellectual Product|General Exam|2903,2906|true|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Pathologic Function|General Exam|2914,2928|true|false|false|C1504476|Pronator drift|Pronator Drift
Event|Event|General Exam|2923,2928|true|false|false|||Drift
Finding|Finding|General Exam|2933,2936|true|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Gene or Genome|General Exam|2933,2936|true|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Idea or Concept|General Exam|2933,2936|true|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Intellectual Product|General Exam|2933,2936|true|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Event|Event|General Exam|2946,2952|true|false|false|||Speech
Finding|Organism Function|General Exam|2946,2952|true|false|false|C0037817|Speech|Speech
Procedure|Diagnostic Procedure|General Exam|2946,2952|true|false|false|C0846595|Speech assessment|Speech
Finding|Finding|General Exam|2964,2967|true|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Gene or Genome|General Exam|2964,2967|true|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Idea or Concept|General Exam|2964,2967|true|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Intellectual Product|General Exam|2964,2967|true|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Mental Process|General Exam|2975,2988|true|false|false|C0162340|Comprehension|Comprehension
Event|Event|General Exam|2989,2995|true|false|false|||Intact
Finding|Finding|General Exam|2989,2995|true|false|false|C1554187|Gender Status - Intact|Intact
Finding|Finding|General Exam|3000,3003|true|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Gene or Genome|General Exam|3000,3003|true|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Idea or Concept|General Exam|3000,3003|true|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Intellectual Product|General Exam|3000,3003|true|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Event|Event|General Exam|3011,3016|true|false|false|||Motor
Finding|Functional Concept|General Exam|3011,3016|true|false|false|C1513492|motor movement|Motor
Finding|Functional Concept|General Exam|3047,3052|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Finding|Functional Concept|General Exam|3088,3092|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Event|Event|General Exam|3249,3258|false|false|false|||Sensation
Finding|Finding|General Exam|3249,3258|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Finding|Organ or Tissue Function|General Exam|3249,3258|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Procedure|Health Care Activity|General Exam|3249,3258|false|false|false|C2229507|sensory exam|Sensation
Event|Event|General Exam|3259,3265|false|false|false|||intact
Finding|Finding|General Exam|3259,3265|false|false|false|C1554187|Gender Status - Intact|intact
Drug|Amino Acid, Peptide, or Protein|General Exam|3269,3274|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|General Exam|3269,3274|false|false|false|C1570446|TNFSF14 protein, human|light
Finding|Finding|General Exam|3269,3274|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|General Exam|3269,3274|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|General Exam|3269,3274|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|General Exam|3269,3274|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|General Exam|3269,3274|false|false|false|C0031765|Phototherapy|light
Finding|Physiologic Function|General Exam|3269,3280|false|false|false|C0423553|Light touch|light touch
Event|Event|General Exam|3275,3280|false|false|false|||touch
Finding|Mental Process|General Exam|3275,3280|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Finding|Organ or Tissue Function|General Exam|3275,3280|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Procedure|Therapeutic or Preventive Procedure|General Exam|3275,3280|false|false|false|C0152054|Therapeutic Touch|touch
Event|Event|General Exam|3310,3313|false|false|false|||see
Event|Event|General Exam|3314,3317|false|false|false|||OMR
Finding|Gene or Genome|General Exam|3314,3317|false|false|false|C1412647|ATP5F1A gene|OMR
Event|Event|General Exam|3332,3335|false|false|false|||lab
Finding|Gene or Genome|General Exam|3332,3335|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|lab
Finding|Intellectual Product|General Exam|3332,3335|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|lab
Finding|Finding|General Exam|3340,3347|false|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|General Exam|3340,3347|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Event|Event|General Exam|3348,3355|false|false|false|||results
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|3383,3388|false|false|false|C0006104;C4266577|Brain;Head>Brain|Brain
Disorder|Disease or Syndrome|Hospital Course|3383,3388|false|false|false|C0006111|Brain Diseases|Brain
Finding|Finding|Hospital Course|3383,3395|false|false|false|C0221505|Lesion of brain|Brain lesion
Event|Event|Hospital Course|3389,3395|false|false|false|||lesion
Finding|Finding|Hospital Course|3389,3395|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|Hospital Course|3389,3395|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Body Substance|Hospital Course|3396,3403|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|3396,3403|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|3396,3403|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|3408,3413|false|false|false|||found
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|3422,3432|false|false|false|C0007765|Cerebellum|cerebellar
Event|Event|Hospital Course|3433,3444|false|false|false|||hypodensity
Event|Event|Hospital Course|3460,3463|false|false|false|||OSH
Event|Event|Hospital Course|3465,3467|false|false|false|||CT
Drug|Indicator, Reagent, or Diagnostic Aid|Hospital Course|3473,3481|false|false|false|C0009924|Contrast Media|contrast
Event|Event|Hospital Course|3473,3481|false|false|false|||contrast
Event|Event|Hospital Course|3486,3494|false|false|false|||obtained
Event|Event|Hospital Course|3529,3539|false|false|false|||concerning
Event|Event|Hospital Course|3544,3554|false|false|false|||underlying
Finding|Finding|Hospital Course|3555,3559|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|Hospital Course|3555,3559|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Hospital Course|3555,3559|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Disorder|Neoplastic Process|Hospital Course|3555,3566|false|false|false|C0746408|mass lesion|mass lesion
Event|Event|Hospital Course|3560,3566|false|false|false|||lesion
Finding|Finding|Hospital Course|3560,3566|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|Hospital Course|3560,3566|false|false|false|C0221198;C1546698|Lesion|lesion
Disorder|Disease or Syndrome|Hospital Course|3572,3585|false|false|false|C0020255|Hydrocephalus|hydrocephalus
Event|Event|Hospital Course|3572,3585|false|false|false|||hydrocephalus
Event|Event|Hospital Course|3605,3611|false|false|false|||unable
Finding|Finding|Hospital Course|3605,3611|false|false|false|C1299582|Unable|unable
Event|Event|Hospital Course|3619,3622|false|false|false|||MRI
Finding|Gene or Genome|Hospital Course|3619,3622|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|Hospital Course|3619,3622|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|Hospital Course|3619,3622|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Finding|Pathologic Function|Hospital Course|3666,3674|false|false|false|C0002940|Aneurysm|aneurysm
Event|Event|Hospital Course|3675,3679|false|false|false|||clip
Finding|Gene or Genome|Hospital Course|3675,3679|false|false|false|C1337111;C1413237;C1561603;C1704793;C1824746;C1824747;C2827463|CD74 gene;CLIP - Codes for radiology reports;CLIP1 gene;CLIP1 wt Allele;CLIP2 gene;POMC gene;POMC wt Allele|clip
Finding|Intellectual Product|Hospital Course|3675,3679|false|false|false|C1337111;C1413237;C1561603;C1704793;C1824746;C1824747;C2827463|CD74 gene;CLIP - Codes for radiology reports;CLIP1 gene;CLIP1 wt Allele;CLIP2 gene;POMC gene;POMC wt Allele|clip
Procedure|Health Care Activity|Hospital Course|3675,3679|false|false|false|C5552742|Comprehensive Lifestyle Intervention Program|clip
Event|Event|Hospital Course|3689,3695|false|false|false|||placed
Finding|Body Substance|Hospital Course|3712,3719|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|3712,3719|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|3712,3719|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|3724,3732|false|false|false|||admitted
Event|Event|Hospital Course|3748,3753|false|false|false|||close
Finding|Finding|Hospital Course|3748,3753|false|false|false|C0587267;C3810854|Close;Closed|close
Finding|Functional Concept|Hospital Course|3748,3753|false|false|false|C0587267;C3810854|Close;Closed|close
Event|Activity|Hospital Course|3755,3765|false|false|false|C1283169||monitoring
Event|Event|Hospital Course|3755,3765|false|false|false|||monitoring
Procedure|Health Care Activity|Hospital Course|3755,3765|false|false|false|C0150369|Preventive monitoring|monitoring
Procedure|Health Care Activity|Hospital Course|3770,3778|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3770,3778|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Event|Event|Hospital Course|3779,3787|false|false|false|||planning
Finding|Functional Concept|Hospital Course|3779,3787|false|false|false|C0032074;C1301732|Planned|planning
Finding|Mental Process|Hospital Course|3779,3787|false|false|false|C0032074;C1301732|Planned|planning
Event|Event|Hospital Course|3797,3804|false|false|false|||started
Drug|Organic Chemical|Hospital Course|3809,3822|false|false|false|C0011777|dexamethasone|dexamethasone
Drug|Pharmacologic Substance|Hospital Course|3809,3822|false|false|false|C0011777|dexamethasone|dexamethasone
Finding|Finding|Hospital Course|3836,3840|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|Hospital Course|3836,3840|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Hospital Course|3836,3840|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Finding|Hospital Course|3836,3847|false|false|false|C4086564|Mass Effect|mass effect
Event|Event|Hospital Course|3841,3847|false|false|false|||effect
Anatomy|Body Location or Region|Hospital Course|3852,3857|false|false|false|C0460005|Trunk structure|torso
Event|Event|Hospital Course|3862,3870|false|false|false|||obtained
Event|Event|Hospital Course|3878,3884|false|false|false|||showed
Anatomy|Body Location or Region|Hospital Course|3889,3893|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|3889,3893|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Hospital Course|3889,3893|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Hospital Course|3889,3893|false|false|false|C0740941|Lung Problem|lung
Finding|Finding|Hospital Course|3889,3901|false|false|false|C0034079||lung nodules
Event|Event|Hospital Course|3894,3901|false|false|false|||nodules
Event|Event|Hospital Course|3903,3906|false|false|false|||see
Event|Event|Hospital Course|3922,3933|false|false|false|||information
Finding|Idea or Concept|Hospital Course|3922,3933|false|false|false|C0870705;C1533716;C1561527;C1561528|Acknowledgement Detail Type - Information;Error severity - Information;Information;control act - information|information
Finding|Intellectual Product|Hospital Course|3922,3933|false|false|false|C0870705;C1533716;C1561527;C1561528|Acknowledgement Detail Type - Information;Error severity - Information;Information;control act - information|information
Phenomenon|Natural Phenomenon or Process|Hospital Course|3946,3955|false|false|false|C0034519;C0851346|Electromagnetic Radiation;Radiation|radiation
Procedure|Research Activity|Hospital Course|3946,3955|false|false|false|C1522449;C1524020;C1524021|Radiation Ionizing Radiotherapy;Radiation therapy (procedure);Radiotherapy Research|radiation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3946,3955|false|false|false|C1522449;C1524020;C1524021|Radiation Ionizing Radiotherapy;Radiation therapy (procedure);Radiotherapy Research|radiation
Procedure|Laboratory Procedure|Hospital Course|3946,3964|false|false|false|C2183259|diagnostic service sources radiology labs radiation oncology|radiation oncology
Disorder|Neoplastic Process|Hospital Course|3956,3964|false|false|false|C0027651|Neoplasms|oncology
Event|Event|Hospital Course|3956,3964|false|false|false|||oncology
Procedure|Health Care Activity|Hospital Course|3956,3964|false|false|false|C1555459|oncology services|oncology
Event|Event|Hospital Course|3970,3979|false|false|false|||consulted
Disorder|Disease or Syndrome|Hospital Course|3981,3985|false|false|false|C0270724|Infantile Neuroaxonal Dystrophy|Plan
Event|Event|Hospital Course|3981,3985|false|false|false|||Plan
Finding|Functional Concept|Hospital Course|3981,3985|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|Plan
Finding|Intellectual Product|Hospital Course|3981,3985|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|Plan
Finding|Mental Process|Hospital Course|3981,3985|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|Plan
Procedure|Health Care Activity|Hospital Course|4000,4008|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4000,4008|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4000,4018|false|false|false|C0015252;C0728940|Excision;removal technique|surgical resection
Event|Event|Hospital Course|4009,4018|false|false|false|||resection
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4009,4018|false|false|false|C0015252;C0728940|Excision;removal technique|resection
Event|Event|Hospital Course|4026,4032|false|false|false|||lesion
Finding|Finding|Hospital Course|4026,4032|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|Hospital Course|4026,4032|false|false|false|C0221198;C1546698|Lesion|lesion
Event|Event|Hospital Course|4049,4059|false|false|false|||determined
Finding|Pathologic Function|Hospital Course|4070,4078|false|false|false|C0002940|Aneurysm|aneurysm
Event|Event|Hospital Course|4079,4083|false|false|false|||clip
Finding|Gene or Genome|Hospital Course|4079,4083|false|false|false|C1337111;C1413237;C1561603;C1704793;C1824746;C1824747;C2827463|CD74 gene;CLIP - Codes for radiology reports;CLIP1 gene;CLIP1 wt Allele;CLIP2 gene;POMC gene;POMC wt Allele|clip
Finding|Intellectual Product|Hospital Course|4079,4083|false|false|false|C1337111;C1413237;C1561603;C1704793;C1824746;C1824747;C2827463|CD74 gene;CLIP - Codes for radiology reports;CLIP1 gene;CLIP1 wt Allele;CLIP2 gene;POMC gene;POMC wt Allele|clip
Procedure|Health Care Activity|Hospital Course|4079,4083|false|false|false|C5552742|Comprehensive Lifestyle Intervention Program|clip
Event|Event|Hospital Course|4088,4091|false|false|false|||MRI
Finding|Gene or Genome|Hospital Course|4088,4091|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|Hospital Course|4088,4091|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|Hospital Course|4088,4091|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Event|Event|Hospital Course|4092,4102|false|false|false|||compatible
Finding|Idea or Concept|Hospital Course|4092,4102|false|false|false|C0332290|Consistent with|compatible
Event|Event|Hospital Course|4115,4119|false|false|false|||able
Finding|Finding|Hospital Course|4115,4119|false|false|false|C1299581|Able (qualifier value)|able
Event|Event|Hospital Course|4131,4134|false|false|false|||MRI
Finding|Gene or Genome|Hospital Course|4131,4134|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|Hospital Course|4131,4134|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|Hospital Course|4131,4134|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Diagnostic Procedure|Hospital Course|4131,4140|false|false|false|C4028269|Nuclear magnetic resonance imaging brain|MRI Brain
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4135,4140|false|false|false|C0006104;C4266577|Brain;Head>Brain|Brain
Disorder|Disease or Syndrome|Hospital Course|4135,4140|false|false|false|C0006111|Brain Diseases|Brain
Event|Event|Hospital Course|4135,4140|false|false|false|||Brain
Procedure|Health Care Activity|Hospital Course|4145,4153|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4145,4153|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Event|Event|Hospital Course|4154,4162|false|false|false|||planning
Finding|Functional Concept|Hospital Course|4154,4162|false|false|false|C0032074;C1301732|Planned|planning
Finding|Mental Process|Hospital Course|4154,4162|false|false|false|C0032074;C1301732|Planned|planning
Event|Event|Hospital Course|4168,4172|false|false|false|||went
Event|Event|Hospital Course|4188,4195|false|false|false|||evening
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4209,4232|false|false|false|C2066670|suboccipital craniotomy|suboccipital craniotomy
Event|Event|Hospital Course|4222,4232|false|false|false|||craniotomy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4222,4232|false|false|false|C0010280|Craniotomy|craniotomy
Event|Event|Hospital Course|4237,4246|false|false|false|||resection
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4237,4246|false|false|false|C0015252;C0728940|Excision;removal technique|resection
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4255,4265|false|false|false|C0007765|Cerebellum|cerebellar
Disorder|Disease or Syndrome|Hospital Course|4255,4272|false|false|false|C0742035||cerebellar lesion
Event|Event|Hospital Course|4266,4272|false|false|false|||lesion
Finding|Finding|Hospital Course|4266,4272|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|Hospital Course|4266,4272|false|false|false|C0221198;C1546698|Lesion|lesion
Event|Event|Hospital Course|4298,4307|false|false|false|||monitored
Anatomy|Body Space or Junction|Hospital Course|4318,4321|false|false|false|C0228479|Structure of intraculminate fissure|ICU
Event|Event|Hospital Course|4318,4321|false|false|false|||ICU
Finding|Intellectual Product|Hospital Course|4318,4321|false|false|false|C4554035|Inventory of Callous-Unemotional Traits|ICU
Event|Event|Hospital Course|4333,4341|false|false|false|||remained
Event|Event|Hospital Course|4378,4384|false|false|false|||stable
Finding|Intellectual Product|Hospital Course|4378,4384|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|Hospital Course|4394,4405|false|false|false|||transferred
Anatomy|Anatomical Structure|Hospital Course|4435,4440|false|false|false|C3714591|Floor (anatomic)|floor
Attribute|Clinical Attribute|Hospital Course|4442,4448|false|false|false|C5889824||status
Event|Event|Hospital Course|4442,4448|false|false|false|||status
Finding|Idea or Concept|Hospital Course|4442,4448|false|false|false|C1546481|What subject filter - Status|status
Drug|Organic Chemical|Hospital Course|4454,4467|false|false|false|C0011777|dexamethasone|Dexamethasone
Drug|Pharmacologic Substance|Hospital Course|4454,4467|false|false|false|C0011777|dexamethasone|Dexamethasone
Event|Event|Hospital Course|4454,4467|false|false|false|||Dexamethasone
Event|Event|Hospital Course|4472,4479|false|false|false|||ordered
Event|Event|Hospital Course|4483,4488|false|false|false|||taper
Event|Activity|Hospital Course|4500,4511|false|false|false|C0024501|Maintenance|maintenance
Event|Event|Hospital Course|4512,4516|false|false|false|||dose
Disorder|Mental or Behavioral Dysfunction|Hospital Course|4524,4527|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4524,4527|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|4524,4527|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|4524,4527|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|4524,4527|false|false|false|C1332410|BID gene|BID
Finding|Intellectual Product|Hospital Course|4551,4555|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|Hospital Course|4562,4571|false|false|false|||pathology
Finding|Functional Concept|Hospital Course|4562,4571|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Finding|Pathologic Function|Hospital Course|4562,4571|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Procedure|Laboratory Procedure|Hospital Course|4562,4571|false|false|false|C0919386|Pathology procedure|pathology
Event|Event|Hospital Course|4572,4581|false|false|false|||finalized
Disorder|Neoplastic Process|Hospital Course|4585,4610|false|false|false|C0149925|Small cell carcinoma of lung|small cell lung carcinoma
Anatomy|Cell|Hospital Course|4591,4595|false|false|false|C0007634|Cells|cell
Finding|Gene or Genome|Hospital Course|4591,4595|false|false|false|C1413336;C1413337|CEL gene;CELP gene|cell
Anatomy|Body Location or Region|Hospital Course|4596,4600|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4596,4600|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Hospital Course|4596,4600|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Hospital Course|4596,4600|false|false|false|C0740941|Lung Problem|lung
Disorder|Neoplastic Process|Hospital Course|4596,4610|false|false|false|C0684249|Carcinoma of lung|lung carcinoma
Disorder|Neoplastic Process|Hospital Course|4601,4610|false|false|false|C0007097|Carcinoma|carcinoma
Event|Event|Hospital Course|4601,4610|false|false|false|||carcinoma
Anatomy|Body Location or Region|Hospital Course|4615,4619|false|false|false|C0024109;C4037972|Chest>Lung;Lung|Lung
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4615,4619|false|false|false|C0024109;C4037972|Chest>Lung;Lung|Lung
Disorder|Disease or Syndrome|Hospital Course|4615,4619|false|false|false|C0024115|Lung diseases|Lung
Finding|Finding|Hospital Course|4615,4619|false|false|false|C0740941|Lung Problem|Lung
Event|Event|Hospital Course|4620,4627|false|false|false|||lesions
Finding|Finding|Hospital Course|4620,4627|false|false|false|C0221198|Lesion|lesions
Anatomy|Body Location or Region|Hospital Course|4631,4636|false|false|false|C0460005|Trunk structure|torso
Event|Event|Hospital Course|4641,4649|false|false|false|||obtained
Event|Event|Hospital Course|4656,4662|false|false|false|||showed
Anatomy|Body Location or Region|Hospital Course|4667,4671|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4667,4671|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Hospital Course|4667,4671|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Hospital Course|4667,4671|false|false|false|C0740941|Lung Problem|lung
Finding|Finding|Hospital Course|4667,4679|false|false|false|C0034079||lung nodules
Event|Event|Hospital Course|4672,4679|false|false|false|||nodules
Finding|Functional Concept|Hospital Course|4693,4697|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4722,4728|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4722,4733|false|false|false|C0003489;C4037976|Aortic arch structure;Chest>Aortic arch|aortic arch
Disorder|Anatomical Abnormality|Hospital Course|4722,4733|false|false|false|C4759703|Aortic arch malformation|aortic arch
Anatomy|Body Location or Region|Hospital Course|4729,4733|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4729,4733|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Anatomy|Body Space or Junction|Hospital Course|4729,4733|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Finding|Finding|Hospital Course|4729,4733|false|false|false|C1538146;C4722404|Age-Related Clonal Hematopoiesis;ZBTB8OS gene|arch
Finding|Gene or Genome|Hospital Course|4729,4733|false|false|false|C1538146;C4722404|Age-Related Clonal Hematopoiesis;ZBTB8OS gene|arch
Finding|Functional Concept|Hospital Course|4756,4761|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4756,4772|false|false|false|C1261074|Structure of right upper lobe of lung|right upper lobe
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4762,4772|false|false|false|C0225756|Structure of upper lobe of lung|upper lobe
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4768,4772|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|Hospital Course|4768,4772|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4774,4783|true|false|false|C0024109|Lung|Pulmonary
Attribute|Clinical Attribute|Hospital Course|4774,4783|true|false|false|C2707265||Pulmonary
Finding|Finding|Hospital Course|4774,4783|true|false|false|C4522268|Pulmonary (intended site)|Pulmonary
Event|Event|Hospital Course|4788,4797|true|false|false|||consulted
Event|Event|Hospital Course|4802,4808|true|false|false|||stated
Event|Event|Hospital Course|4826,4838|true|false|false|||intervention
Procedure|Health Care Activity|Hospital Course|4826,4838|true|false|false|C0184661;C0886296;C1273869|Intervention regimes;Interventional procedure;Nursing interventions|intervention
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4826,4838|true|false|false|C0184661;C0886296;C1273869|Intervention regimes;Interventional procedure;Nursing interventions|intervention
Event|Event|Hospital Course|4843,4852|true|false|false|||indicated
Finding|Idea or Concept|Hospital Course|4859,4864|true|false|false|C1546485|Diagnosis Type - Final|final
Event|Event|Hospital Course|4865,4874|false|false|false|||pathology
Finding|Functional Concept|Hospital Course|4865,4874|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Finding|Pathologic Function|Hospital Course|4865,4874|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Procedure|Laboratory Procedure|Hospital Course|4865,4874|false|false|false|C0919386|Pathology procedure|pathology
Event|Event|Hospital Course|4880,4884|false|false|false|||back
Drug|Biologically Active Substance|Hospital Course|4886,4890|false|false|false|C0018966|Heme|Heme
Drug|Organic Chemical|Hospital Course|4886,4890|false|false|false|C0018966|Heme|Heme
Event|Event|Hospital Course|4904,4913|true|false|false|||consulted
Event|Event|Hospital Course|4924,4939|true|false|false|||recommendations
Finding|Idea or Concept|Hospital Course|4924,4939|true|false|false|C0034866|Recommendation|recommendations
Anatomy|Body Location or Region|Hospital Course|4957,4961|true|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4957,4961|true|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Hospital Course|4957,4961|true|false|false|C0024115|Lung diseases|lung
Finding|Finding|Hospital Course|4957,4961|true|false|false|C0740941|Lung Problem|lung
Procedure|Diagnostic Procedure|Hospital Course|4957,4969|true|false|false|C0203683|Radioisotope scan of lung|lung imaging
Event|Event|Hospital Course|4962,4969|true|false|false|||imaging
Finding|Finding|Hospital Course|4962,4969|true|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|Hospital Course|4962,4969|true|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Anatomy|Body Location or Region|Hospital Course|4982,4986|true|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4982,4986|true|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Hospital Course|4982,4986|true|false|false|C0024115|Lung diseases|lung
Finding|Finding|Hospital Course|4982,4986|true|false|false|C0740941|Lung Problem|lung
Procedure|Diagnostic Procedure|Hospital Course|4982,4993|true|false|false|C0189485|Biopsy of lung|lung biopsy
Event|Event|Hospital Course|4987,4993|true|false|false|||biopsy
Finding|Finding|Hospital Course|4987,4993|true|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Finding|Intellectual Product|Hospital Course|4987,4993|true|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Procedure|Diagnostic Procedure|Hospital Course|4987,4993|true|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Procedure|Health Care Activity|Hospital Course|4987,4993|true|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Event|Event|Hospital Course|4998,5004|false|false|false|||needed
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5012,5021|false|false|false|C0024109|Lung|Pulmonary
Attribute|Clinical Attribute|Hospital Course|5012,5021|false|false|false|C2707265||Pulmonary
Finding|Finding|Hospital Course|5012,5021|false|false|false|C4522268|Pulmonary (intended site)|Pulmonary
Drug|Biologically Active Substance|Hospital Course|5026,5030|false|false|false|C0018966|Heme|Heme
Drug|Organic Chemical|Hospital Course|5026,5030|false|false|false|C0018966|Heme|Heme
Event|Event|Hospital Course|5035,5041|false|false|false|||stated
Event|Event|Hospital Course|5047,5054|false|false|false|||staging
Finding|Functional Concept|Hospital Course|5047,5054|false|false|false|C0332305|With staging|staging
Event|Event|Hospital Course|5059,5068|false|false|false|||treatment
Finding|Conceptual Entity|Hospital Course|5059,5068|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Hospital Course|5059,5068|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Hospital Course|5059,5068|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5059,5068|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Event|Event|Hospital Course|5079,5089|false|false|false|||determined
Anatomy|Tissue|Hospital Course|5103,5109|false|false|false|C0040300|Body tissue|tissue
Finding|Intellectual Product|Hospital Course|5103,5109|false|false|false|C1547928|Tissue Specimen Code|tissue
Event|Event|Hospital Course|5110,5119|false|false|false|||pathology
Finding|Functional Concept|Hospital Course|5110,5119|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Finding|Pathologic Function|Hospital Course|5110,5119|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Procedure|Laboratory Procedure|Hospital Course|5110,5119|false|false|false|C0919386|Pathology procedure|pathology
Event|Event|Hospital Course|5125,5134|false|false|false|||resection
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5125,5134|false|false|false|C0015252;C0728940|Excision;removal technique|resection
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5143,5148|false|false|false|C0006104;C4266577|Brain;Head>Brain|brain
Disorder|Disease or Syndrome|Hospital Course|5143,5148|false|false|false|C0006111|Brain Diseases|brain
Finding|Finding|Hospital Course|5143,5155|false|false|false|C0221505|Lesion of brain|brain lesion
Event|Event|Hospital Course|5149,5155|false|false|false|||lesion
Finding|Finding|Hospital Course|5149,5155|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|Hospital Course|5149,5155|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Idea or Concept|Hospital Course|5161,5166|false|false|false|C1546485|Diagnosis Type - Final|final
Event|Event|Hospital Course|5167,5176|false|false|false|||pathology
Finding|Functional Concept|Hospital Course|5167,5176|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Finding|Pathologic Function|Hospital Course|5167,5176|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Procedure|Laboratory Procedure|Hospital Course|5167,5176|false|false|false|C0919386|Pathology procedure|pathology
Event|Event|Hospital Course|5177,5181|false|false|false|||came
Anatomy|Cell|Hospital Course|5196,5200|false|false|false|C0007634|Cells|cell
Finding|Gene or Genome|Hospital Course|5196,5200|false|false|false|C1413336;C1413337|CEL gene;CELP gene|cell
Anatomy|Body Location or Region|Hospital Course|5202,5206|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5202,5206|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Hospital Course|5202,5206|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Hospital Course|5202,5206|false|false|false|C0740941|Lung Problem|lung
Disorder|Neoplastic Process|Hospital Course|5202,5216|false|false|false|C0684249|Carcinoma of lung|lung carcinoma
Disorder|Neoplastic Process|Hospital Course|5207,5216|false|false|false|C0007097|Carcinoma|carcinoma
Event|Event|Hospital Course|5207,5216|false|false|false|||carcinoma
Event|Event|Hospital Course|5227,5233|false|false|false|||follow
Anatomy|Body Location or Region|Hospital Course|5246,5254|false|false|false|C0817096|Chest|thoracic
Disorder|Disease or Syndrome|Hospital Course|5246,5254|false|false|false|C5779551|Dissecting Thoracic Aortic Aneurysm|thoracic
Drug|Organic Chemical|Hospital Course|5278,5285|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|Steroid
Drug|Pharmacologic Substance|Hospital Course|5278,5285|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|Steroid
Disorder|Disease or Syndrome|Hospital Course|5278,5307|false|false|false|C0745098|Hyperglycemia steroid-induced|Steroid-induced hyperglycemia
Disorder|Disease or Syndrome|Hospital Course|5294,5307|false|false|false|C0020456|Hyperglycemia|hyperglycemia
Event|Event|Hospital Course|5294,5307|false|false|false|||hyperglycemia
Finding|Finding|Hospital Course|5294,5307|false|false|false|C2919432|Glucose in blood specimen above reference range|hyperglycemia
Event|Event|Hospital Course|5323,5332|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|5323,5332|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Body Substance|Hospital Course|5338,5345|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|5338,5345|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|5338,5345|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|5361,5369|false|false|false|||required
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5379,5384|false|false|false|C0222045|Integumentary scale|scale
Event|Activity|Hospital Course|5379,5384|false|false|false|C1947916|Scaling|scale
Finding|Conceptual Entity|Hospital Course|5379,5384|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Finding|Intellectual Product|Hospital Course|5379,5384|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5385,5392|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Hormone|Hospital Course|5385,5392|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Pharmacologic Substance|Hospital Course|5385,5392|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Event|Event|Hospital Course|5385,5392|false|false|false|||Insulin
Finding|Gene or Genome|Hospital Course|5385,5392|false|false|false|C1337112|INS gene|Insulin
Procedure|Laboratory Procedure|Hospital Course|5385,5392|false|false|false|C0202098|Insulin measurement|Insulin
Disorder|Disease or Syndrome|Hospital Course|5406,5411|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Hospital Course|5406,5411|false|false|false|||blood
Finding|Body Substance|Hospital Course|5406,5411|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Organic Chemical|Hospital Course|5406,5418|false|false|false|C0005802|Blood Glucose|blood sugars
Drug|Organic Chemical|Hospital Course|5412,5418|false|false|false|C0242209|Sugars|sugars
Drug|Pharmacologic Substance|Hospital Course|5412,5418|false|false|false|C0242209|Sugars|sugars
Event|Event|Hospital Course|5412,5418|false|false|false|||sugars
Procedure|Laboratory Procedure|Hospital Course|5412,5418|false|false|false|C2239291|sugars (lab test)|sugars
Drug|Organic Chemical|Hospital Course|5429,5442|false|false|false|C0011777|dexamethasone|Dexamethasone
Drug|Pharmacologic Substance|Hospital Course|5429,5442|false|false|false|C0011777|dexamethasone|Dexamethasone
Event|Event|Hospital Course|5429,5442|false|false|false|||Dexamethasone
Event|Event|Hospital Course|5452,5461|false|false|false|||evaluated
Event|Event|Hospital Course|5473,5482|false|false|false|||inpatient
Finding|Idea or Concept|Hospital Course|5473,5482|false|false|false|C1548438;C1549404|Patient Class - Inpatient;Referral category - Inpatient|inpatient
Procedure|Health Care Activity|Hospital Course|5473,5482|false|false|false|C1555324|inpatient encounter|inpatient
Event|Event|Hospital Course|5501,5508|false|false|false|||decided
Event|Event|Hospital Course|5526,5530|true|false|false|||need
Event|Event|Hospital Course|5537,5541|true|false|false|||home
Finding|Idea or Concept|Hospital Course|5537,5541|true|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|5537,5541|true|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|5537,5541|true|false|false|C1553498|home health encounter|home
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5545,5552|true|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Hormone|Hospital Course|5545,5552|true|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Pharmacologic Substance|Hospital Course|5545,5552|true|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Event|Event|Hospital Course|5545,5552|true|false|false|||Insulin
Finding|Gene or Genome|Hospital Course|5545,5552|true|false|false|C1337112|INS gene|Insulin
Procedure|Laboratory Procedure|Hospital Course|5545,5552|true|false|false|C0202098|Insulin measurement|Insulin
Event|Event|Hospital Course|5560,5571|false|false|false|||recommended
Event|Event|Hospital Course|5572,5583|false|false|false|||discharging
Event|Event|Hospital Course|5595,5605|false|false|false|||glucometer
Event|Event|Hospital Course|5625,5630|false|false|false|||check
Disorder|Disease or Syndrome|Hospital Course|5635,5640|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Hospital Course|5635,5640|false|false|false|||blood
Finding|Body Substance|Hospital Course|5635,5640|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Organic Chemical|Hospital Course|5635,5647|false|false|false|C0005802|Blood Glucose|blood sugars
Drug|Organic Chemical|Hospital Course|5641,5647|false|false|false|C0242209|Sugars|sugars
Drug|Pharmacologic Substance|Hospital Course|5641,5647|false|false|false|C0242209|Sugars|sugars
Event|Event|Hospital Course|5641,5647|false|false|false|||sugars
Procedure|Laboratory Procedure|Hospital Course|5641,5647|false|false|false|C2239291|sugars (lab test)|sugars
Finding|Idea or Concept|Hospital Course|5661,5665|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Finding|Intellectual Product|Hospital Course|5661,5665|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Disorder|Disease or Syndrome|Hospital Course|5666,5671|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Hospital Course|5666,5671|false|false|false|||blood
Finding|Body Substance|Hospital Course|5666,5671|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Organic Chemical|Hospital Course|5666,5677|false|false|false|C0005802|Blood Glucose|blood sugar
Procedure|Laboratory Procedure|Hospital Course|5666,5677|false|false|false|C0392201|Blood glucose measurement|blood sugar
Drug|Biomedical or Dental Material|Hospital Course|5672,5677|false|false|false|C0007004;C0242209;C3665462|Carbohydrates;Sugars;raw sugar|sugar
Drug|Organic Chemical|Hospital Course|5672,5677|false|false|false|C0007004;C0242209;C3665462|Carbohydrates;Sugars;raw sugar|sugar
Drug|Pharmacologic Substance|Hospital Course|5672,5677|false|false|false|C0007004;C0242209;C3665462|Carbohydrates;Sugars;raw sugar|sugar
Event|Event|Hospital Course|5678,5682|false|false|false|||less
Event|Event|Hospital Course|5702,5709|false|false|false|||advised
Event|Event|Hospital Course|5713,5719|false|false|false|||record
Event|Event|Hospital Course|5724,5732|false|false|false|||readings
Event|Event|Hospital Course|5737,5743|false|false|false|||follow
Disorder|Disease or Syndrome|Hospital Course|5757,5760|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|Hospital Course|5757,5760|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|Hospital Course|5757,5760|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5757,5760|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|Hospital Course|5757,5760|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|Hospital Course|5757,5760|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|Hospital Course|5757,5760|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|Hospital Course|5757,5760|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|Hospital Course|5757,5760|false|false|false|||PCP
Finding|Gene or Genome|Hospital Course|5757,5760|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|Hospital Course|5757,5760|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|Hospital Course|5773,5784|false|false|false|||Bradycardia
Finding|Finding|Hospital Course|5773,5784|false|false|false|C0428977;C3812171|Bradycardia;Bradycardia by ECG Finding|Bradycardia
Event|Event|Hospital Course|5800,5808|false|false|false|||transfer
Finding|Functional Concept|Hospital Course|5800,5808|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|Hospital Course|5800,5808|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|Hospital Course|5800,5808|false|false|false|C4706767|Transfer (immobility management)|transfer
Finding|Gene or Genome|Hospital Course|5827,5831|false|false|false|C1420638;C1539127;C1710283|CORO7 gene;TCF21 gene;TCF21 wt Allele|POD1
Event|Event|Hospital Course|5846,5850|false|false|false|||kept
Anatomy|Body Space or Junction|Hospital Course|5858,5861|false|false|false|C0228479|Structure of intraculminate fissure|ICU
Finding|Intellectual Product|Hospital Course|5858,5861|false|false|false|C4554035|Inventory of Callous-Unemotional Traits|ICU
Finding|Finding|Hospital Course|5866,5878|false|false|false|C0231221;C0332151|Asymptomatic (finding);Asymptomatic diagnosis of|asymptomatic
Disorder|Disease or Syndrome|Hospital Course|5866,5890|false|false|false|C0741624|Asymptomatic bradycardia|asymptomatic bradycardia
Event|Event|Hospital Course|5879,5890|false|false|false|||bradycardia
Finding|Finding|Hospital Course|5879,5890|false|false|false|C0428977;C3812171|Bradycardia;Bradycardia by ECG Finding|bradycardia
Event|Event|Hospital Course|5908,5916|false|false|false|||remained
Event|Event|Hospital Course|5917,5929|false|false|false|||asymptomatic
Finding|Finding|Hospital Course|5917,5929|false|false|false|C0231221;C0332151|Asymptomatic (finding);Asymptomatic diagnosis of|asymptomatic
Event|Event|Hospital Course|5939,5948|false|false|false|||heartrate
Event|Event|Hospital Course|5949,5957|false|false|false|||improved
Drug|Substance|Hospital Course|5963,5969|false|false|false|C0302908|Liquid substance|fluids
Event|Event|Hospital Course|5963,5969|false|false|false|||fluids
Finding|Body Substance|Hospital Course|5963,5969|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5963,5969|false|false|false|C0016286|Fluid Therapy|fluids
Event|Event|Hospital Course|5976,5990|false|false|false|||administration
Event|Occupational Activity|Hospital Course|5976,5990|false|false|false|C0001554|Administration occupational activities|administration
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5976,5990|false|false|false|C1533734|Administration (procedure)|administration
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5998,6011|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Hormone|Hospital Course|5998,6011|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Organic Chemical|Hospital Course|5998,6011|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Pharmacologic Substance|Hospital Course|5998,6011|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Event|Event|Hospital Course|5998,6011|false|false|false|||levothyroxine
Event|Event|Hospital Course|6033,6039|false|false|false|||dipped
Event|Event|Hospital Course|6060,6068|false|false|false|||remained
Event|Event|Hospital Course|6069,6081|false|false|false|||asymptomatic
Finding|Finding|Hospital Course|6069,6081|false|false|false|C0231221;C0332151|Asymptomatic (finding);Asymptomatic diagnosis of|asymptomatic
Disorder|Disease or Syndrome|Hospital Course|6085,6097|false|false|false|C0015469;C0376175|Bell Palsy;Facial paralysis|Bell's palsy
Event|Event|Hospital Course|6092,6097|false|false|false|||palsy
Finding|Finding|Hospital Course|6092,6097|false|false|false|C0522224;C3887651|Palsy;Paralysed|palsy
Finding|Body Substance|Hospital Course|6102,6109|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|6102,6109|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|6102,6109|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|6114,6121|false|false|false|||resumed
Finding|Idea or Concept|Hospital Course|6129,6133|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|6129,6133|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|6129,6133|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|6134,6146|false|false|false|C0249458|valacyclovir|Valacyclovir
Drug|Pharmacologic Substance|Hospital Course|6134,6146|false|false|false|C0249458|valacyclovir|Valacyclovir
Event|Event|Hospital Course|6134,6146|false|false|false|||Valacyclovir
Event|Event|Hospital Course|6151,6162|false|false|false|||Prenisolone
Event|Event|Hospital Course|6164,6168|false|false|false|||gtts
Procedure|Laboratory Procedure|Hospital Course|6164,6168|false|false|false|C0017741|Glucose tolerance test|gtts
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6173,6180|false|false|false|C0042027|Urinary tract|Urinary
Finding|Sign or Symptom|Hospital Course|6173,6188|false|false|false|C0085606|Urgency of micturition|Urinary urgency
Event|Event|Hospital Course|6181,6188|false|false|false|||urgency
Finding|Body Substance|Hospital Course|6203,6210|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|6203,6210|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|6203,6210|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|6211,6221|false|false|false|||complained
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6225,6232|false|false|false|C0042027|Urinary tract|urinary
Finding|Sign or Symptom|Hospital Course|6225,6240|false|false|false|C0085606|Urgency of micturition|urinary urgency
Event|Event|Hospital Course|6246,6255|false|false|false|||increased
Event|Event|Hospital Course|6256,6265|false|false|false|||frequency
Finding|Intellectual Product|Hospital Course|6256,6265|false|false|false|C3898838;C4321352|Frequency;How Often|frequency
Event|Event|Hospital Course|6275,6283|false|false|false|||negative
Finding|Classification|Hospital Course|6275,6283|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|6275,6283|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|6275,6283|false|false|false|C5237010|Expression Negative|negative
Drug|Biomedical or Dental Material|Hospital Course|6288,6295|false|false|false|C1706355|Culture Dose Form|culture
Event|Event|Hospital Course|6288,6295|false|false|false|||culture
Finding|Functional Concept|Hospital Course|6288,6295|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Finding|Idea or Concept|Hospital Course|6288,6295|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Procedure|Laboratory Procedure|Hospital Course|6288,6295|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|culture
Event|Event|Hospital Course|6300,6308|false|false|false|||negative
Finding|Classification|Hospital Course|6300,6308|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|6300,6308|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|6300,6308|false|false|false|C5237010|Expression Negative|negative
Event|Event|Hospital Course|6315,6323|false|false|false|||symptoms
Finding|Functional Concept|Hospital Course|6315,6323|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Hospital Course|6315,6323|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|Hospital Course|6328,6336|false|false|false|||resolved
Finding|Finding|Hospital Course|6344,6348|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Hospital Course|6344,6348|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Hospital Course|6344,6348|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|Hospital Course|6352,6361|false|false|false|||discharge
Finding|Body Substance|Hospital Course|6352,6361|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|6352,6361|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|6352,6361|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|6352,6361|false|false|false|C0030685|Patient Discharge|discharge
Finding|Body Substance|Hospital Course|6376,6383|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|6376,6383|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|6376,6383|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|6388,6397|false|false|false|||evaluated
Event|Event|Hospital Course|6416,6423|false|false|false|||cleared
Event|Event|Hospital Course|6432,6436|false|false|false|||home
Finding|Idea or Concept|Hospital Course|6432,6436|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|6432,6436|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|6432,6436|false|false|false|C1553498|home health encounter|home
Event|Event|Hospital Course|6443,6451|false|false|false|||services
Event|Occupational Activity|Hospital Course|6443,6451|false|false|false|C0557854|Services|services
Procedure|Health Care Activity|Hospital Course|6443,6451|false|false|false|C1704289|Clinical Service|services
Event|Event|Hospital Course|6461,6471|false|false|false|||discharged
Finding|Intellectual Product|Hospital Course|6482,6488|false|false|false|C1547311|Patient Condition Code - Stable|stable
Attribute|Clinical Attribute|Hospital Course|6489,6498|false|false|false|C3864998||condition
Disorder|Disease or Syndrome|Hospital Course|6489,6498|false|false|false|C0012634|Disease|condition
Event|Event|Hospital Course|6489,6498|false|false|false|||condition
Finding|Conceptual Entity|Hospital Course|6489,6498|false|false|false|C1705253|Logical Condition|condition
Event|Event|Hospital Course|6510,6516|false|false|false|||follow
Attribute|Clinical Attribute|Hospital Course|6538,6549|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|6538,6549|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|6538,6549|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|6538,6549|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|6538,6562|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|6553,6562|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|6553,6562|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6566,6569|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Enzyme|Hospital Course|6566,6569|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Organic Chemical|Hospital Course|6566,6569|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Pharmacologic Substance|Hospital Course|6566,6569|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Event|Event|Hospital Course|6566,6569|false|false|false|||ASA
Finding|Gene or Genome|Hospital Course|6566,6569|false|false|false|C1412553|ARSA gene|ASA
Drug|Organic Chemical|Hospital Course|6577,6588|false|false|false|C0102118|alendronate|Alendronate
Drug|Pharmacologic Substance|Hospital Course|6577,6588|false|false|false|C0102118|alendronate|Alendronate
Drug|Organic Chemical|Hospital Course|6603,6610|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|6603,6610|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|6603,6610|false|false|false|C0042890|Vitamins|Vitamin
Drug|Organic Chemical|Hospital Course|6603,6613|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|Vitamin D3
Drug|Pharmacologic Substance|Hospital Course|6603,6613|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|Vitamin D3
Drug|Vitamin|Hospital Course|6603,6613|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|Vitamin D3
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6632,6645|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Hormone|Hospital Course|6632,6645|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Organic Chemical|Hospital Course|6632,6645|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Pharmacologic Substance|Hospital Course|6632,6645|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6660,6670|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|Hospital Course|6660,6670|false|false|false|C0065374|lisinopril|Lisinopril
Event|Event|Hospital Course|6685,6694|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|6685,6694|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|6685,6694|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|6685,6694|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|6685,6694|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|6685,6706|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|6695,6706|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|6695,6706|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|6695,6706|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|6695,6706|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|6712,6725|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|6712,6725|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Hospital Course|6712,6725|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|6712,6725|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|Hospital Course|6740,6743|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|6744,6748|false|false|false|C2598155||Pain
Event|Event|Hospital Course|6744,6748|false|false|false|||Pain
Finding|Functional Concept|Hospital Course|6744,6748|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Hospital Course|6744,6748|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Intellectual Product|Hospital Course|6751,6755|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Finding|Finding|Hospital Course|6756,6761|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Finding|Sign or Symptom|Hospital Course|6756,6761|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Drug|Organic Chemical|Hospital Course|6768,6777|false|false|false|C0005632|bisacodyl|Bisacodyl
Drug|Pharmacologic Substance|Hospital Course|6768,6777|false|false|false|C0005632|bisacodyl|Bisacodyl
Drug|Organic Chemical|Hospital Course|6802,6815|false|false|false|C0011777|dexamethasone|Dexamethasone
Drug|Pharmacologic Substance|Hospital Course|6802,6815|false|false|false|C0011777|dexamethasone|Dexamethasone
Event|Event|Hospital Course|6802,6815|false|false|false|||Dexamethasone
Drug|Pharmacologic Substance|Hospital Course|6828,6836|false|false|false|C0720099|Duration brand of oxymetazoline|Duration
Event|Event|Hospital Course|6828,6836|false|false|false|||Duration
Event|Event|Hospital Course|6847,6852|false|false|false|||start
Event|Event|Hospital Course|6873,6883|false|false|false|||2tabsq8hrs
Event|Event|Hospital Course|6888,6899|false|false|false|||2tabsq12hrs
Event|Activity|Hospital Course|6901,6912|false|false|false|C0024501|Maintenance|maintenance
Event|Event|Hospital Course|6913,6917|false|false|false|||dose
Attribute|Clinical Attribute|Hospital Course|6929,6935|false|false|false|C1114758||dose #
Event|Event|Hospital Course|6951,6956|false|false|false|||doses
Event|Event|Hospital Course|6957,6959|false|false|false|||RX
Drug|Organic Chemical|Hospital Course|6961,6974|false|false|false|C0011777|dexamethasone|dexamethasone
Drug|Pharmacologic Substance|Hospital Course|6961,6974|false|false|false|C0011777|dexamethasone|dexamethasone
Event|Event|Hospital Course|6961,6974|false|false|false|||dexamethasone
Drug|Biomedical or Dental Material|Hospital Course|6982,6988|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|6992,7000|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|6995,7000|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|6995,7000|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Biomedical or Dental Material|Hospital Course|7035,7041|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|7042,7049|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|7042,7049|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|7058,7066|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|7058,7066|false|false|false|C1692318|docusate|Docusate
Event|Event|Hospital Course|7058,7066|false|false|false|||Docusate
Drug|Organic Chemical|Hospital Course|7058,7073|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|Hospital Course|7058,7073|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|Hospital Course|7067,7073|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|7067,7073|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|7067,7073|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|7067,7073|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|7067,7073|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|7067,7073|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|Hospital Course|7084,7087|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7084,7087|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|7084,7087|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|7084,7087|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|7084,7087|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|7094,7104|false|false|false|C0015620|famotidine|Famotidine
Drug|Pharmacologic Substance|Hospital Course|7094,7104|false|false|false|C0015620|famotidine|Famotidine
Drug|Organic Chemical|Hospital Course|7124,7134|false|false|false|C0015620|famotidine|famotidine
Drug|Pharmacologic Substance|Hospital Course|7124,7134|false|false|false|C0015620|famotidine|famotidine
Event|Event|Hospital Course|7124,7134|false|false|false|||famotidine
Drug|Biomedical or Dental Material|Hospital Course|7143,7149|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|7153,7161|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|7156,7161|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|7156,7161|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|Hospital Course|7170,7173|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|7170,7173|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biomedical or Dental Material|Hospital Course|7185,7191|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|7192,7199|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|7192,7199|false|false|false|C0807726|refill|Refills
Drug|Biomedical or Dental Material|Hospital Course|7208,7220|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Drug|Organic Chemical|Hospital Course|7208,7220|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Event|Event|Hospital Course|7208,7220|false|false|false|||Polyethylene
Drug|Organic Chemical|Hospital Course|7208,7227|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Pharmacologic Substance|Hospital Course|7208,7227|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Hazardous or Poisonous Substance|Hospital Course|7221,7227|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Drug|Organic Chemical|Hospital Course|7221,7227|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Event|Event|Hospital Course|7221,7227|false|false|false|||Glycol
Finding|Gene or Genome|Hospital Course|7242,7245|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|7246,7258|false|false|false|||Constipation
Finding|Sign or Symptom|Hospital Course|7246,7258|false|false|false|C0009806|Constipation|Constipation
Drug|Biologically Active Substance|Hospital Course|7268,7272|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Hospital Course|7268,7272|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Drug|Substance|Hospital Course|7268,7272|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Finding|Intellectual Product|Hospital Course|7268,7272|false|false|false|C1546701|line source specimen code|Line
Drug|Organic Chemical|Hospital Course|7279,7284|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|Hospital Course|7279,7284|false|false|false|C3489575|sennosides, USP|Senna
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7305,7318|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Hormone|Hospital Course|7305,7318|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Organic Chemical|Hospital Course|7305,7318|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Pharmacologic Substance|Hospital Course|7305,7318|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7305,7325|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Hormone|Hospital Course|7305,7325|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Pharmacologic Substance|Hospital Course|7305,7325|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Biologically Active Substance|Hospital Course|7319,7325|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|7319,7325|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|7319,7325|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|7319,7325|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|7319,7325|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|7319,7325|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7348,7358|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|Hospital Course|7348,7358|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Organic Chemical|Hospital Course|7381,7393|false|false|false|C0032950|prednisolone|PrednisoLONE
Drug|Pharmacologic Substance|Hospital Course|7381,7393|false|false|false|C0032950|prednisolone|PrednisoLONE
Drug|Organic Chemical|Hospital Course|7381,7401|false|false|false|C0071839|prednisolone acetate|PrednisoLONE Acetate
Drug|Pharmacologic Substance|Hospital Course|7381,7401|false|false|false|C0071839|prednisolone acetate|PrednisoLONE Acetate
Drug|Organic Chemical|Hospital Course|7394,7401|false|false|false|C0000975|acetate|Acetate
Drug|Pharmacologic Substance|Hospital Course|7394,7401|false|false|false|C0000975|acetate|Acetate
Finding|Functional Concept|Hospital Course|7405,7410|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|Hospital Course|7420,7424|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|Hospital Course|7420,7424|false|false|false|C1705648|Dropping|DROP
Event|Event|Hospital Course|7425,7429|false|false|false|||LEFT
Finding|Functional Concept|Hospital Course|7425,7429|false|false|false|C1552822|Table Cell Horizontal Align - left|LEFT
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7425,7433|false|false|false|C0229090|Left eye structure|LEFT EYE
Procedure|Diagnostic Procedure|Hospital Course|7425,7433|false|false|false|C2141124|examination of left eye|LEFT EYE
Anatomy|Body Location or Region|Hospital Course|7430,7433|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|EYE
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7430,7433|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|EYE
Disorder|Disease or Syndrome|Hospital Course|7430,7433|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|EYE
Disorder|Neoplastic Process|Hospital Course|7430,7433|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|EYE
Event|Event|Hospital Course|7430,7433|false|false|false|||EYE
Finding|Body Substance|Hospital Course|7430,7433|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Finding|Finding|Hospital Course|7430,7433|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Finding|Intellectual Product|Hospital Course|7430,7433|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Drug|Organic Chemical|Hospital Course|7445,7457|false|false|false|C0249458|valacyclovir|ValACYclovir
Drug|Pharmacologic Substance|Hospital Course|7445,7457|false|false|false|C0249458|valacyclovir|ValACYclovir
Drug|Organic Chemical|Hospital Course|7480,7487|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|7480,7487|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|7480,7487|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|Hospital Course|7480,7489|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|Hospital Course|7480,7489|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|Hospital Course|7480,7489|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|Hospital Course|7480,7489|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|Hospital Course|7480,7489|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|Hospital Course|7488,7489|false|false|false|||D
Event|Event|Hospital Course|7494,7498|false|false|false|||UNIT
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7514,7518|false|false|false|C0675390|ARID1A protein, human|HELD
Drug|Biologically Active Substance|Hospital Course|7514,7518|false|false|false|C0675390|ARID1A protein, human|HELD
Event|Event|Hospital Course|7514,7518|false|false|false|||HELD
Finding|Gene or Genome|Hospital Course|7514,7518|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|HELD
Finding|Idea or Concept|Hospital Course|7514,7518|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|HELD
Drug|Organic Chemical|Hospital Course|7520,7531|false|false|false|C0102118|alendronate|Alendronate
Drug|Pharmacologic Substance|Hospital Course|7520,7531|false|false|false|C0102118|alendronate|Alendronate
Drug|Organic Chemical|Hospital Course|7520,7538|false|false|false|C0700482|alendronate sodium|Alendronate Sodium
Drug|Pharmacologic Substance|Hospital Course|7520,7538|false|false|false|C0700482|alendronate sodium|Alendronate Sodium
Drug|Biologically Active Substance|Hospital Course|7532,7538|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|7532,7538|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|7532,7538|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|7532,7538|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|7532,7538|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|7532,7538|false|false|false|C0337443|Sodium measurement|Sodium
Finding|Intellectual Product|Hospital Course|7551,7555|false|false|false|C1561540|Transaction counts and value totals - week|WEEK
Drug|Pharmacologic Substance|Hospital Course|7569,7579|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Hospital Course|7569,7579|false|false|false|||medication
Finding|Intellectual Product|Hospital Course|7569,7579|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Hospital Course|7584,7588|false|false|false|||held
Event|Event|Hospital Course|7597,7604|true|false|false|||restart
Drug|Organic Chemical|Hospital Course|7605,7616|true|false|false|C0102118|alendronate|Alendronate
Drug|Pharmacologic Substance|Hospital Course|7605,7616|true|false|false|C0102118|alendronate|Alendronate
Drug|Organic Chemical|Hospital Course|7605,7623|true|false|false|C0700482|alendronate sodium|Alendronate Sodium
Drug|Pharmacologic Substance|Hospital Course|7605,7623|true|false|false|C0700482|alendronate sodium|Alendronate Sodium
Drug|Biologically Active Substance|Hospital Course|7617,7623|true|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|7617,7623|true|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|7617,7623|true|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|7617,7623|true|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|7617,7623|true|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|7617,7623|true|false|false|C0337443|Sodium measurement|Sodium
Event|Event|Hospital Course|7630,7633|true|false|false|||POD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7649,7653|false|false|false|C0675390|ARID1A protein, human|HELD
Drug|Biologically Active Substance|Hospital Course|7649,7653|false|false|false|C0675390|ARID1A protein, human|HELD
Event|Event|Hospital Course|7649,7653|false|false|false|||HELD
Finding|Gene or Genome|Hospital Course|7649,7653|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|HELD
Finding|Idea or Concept|Hospital Course|7649,7653|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|HELD
Drug|Organic Chemical|Hospital Course|7655,7662|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Hospital Course|7655,7662|false|false|false|C0004057|aspirin|Aspirin
Event|Event|Hospital Course|7655,7662|false|false|false|||Aspirin
Drug|Pharmacologic Substance|Hospital Course|7684,7694|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Hospital Course|7684,7694|false|false|false|||medication
Finding|Intellectual Product|Hospital Course|7684,7694|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Hospital Course|7699,7703|false|false|false|||held
Event|Event|Hospital Course|7713,7720|true|false|false|||restart
Drug|Organic Chemical|Hospital Course|7721,7728|true|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Hospital Course|7721,7728|true|false|false|C0004057|aspirin|Aspirin
Event|Event|Hospital Course|7721,7728|true|false|false|||Aspirin
Event|Event|Hospital Course|7735,7738|true|false|false|||POD
Event|Event|Hospital Course|7752,7762|false|false|false|||glucometer
Event|Event|Hospital Course|7789,7794|false|false|false|||Check
Disorder|Disease or Syndrome|Hospital Course|7795,7800|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Hospital Course|7795,7800|false|false|false|||blood
Finding|Body Substance|Hospital Course|7795,7800|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Organic Chemical|Hospital Course|7795,7807|false|false|false|C0005802|Blood Glucose|blood sugars
Drug|Organic Chemical|Hospital Course|7801,7807|false|false|false|C0242209|Sugars|sugars
Drug|Pharmacologic Substance|Hospital Course|7801,7807|false|false|false|C0242209|Sugars|sugars
Event|Event|Hospital Course|7801,7807|false|false|false|||sugars
Procedure|Laboratory Procedure|Hospital Course|7801,7807|false|false|false|C2239291|sugars (lab test)|sugars
Event|Event|Hospital Course|7809,7810|false|false|false|||_
Event|Event|Hospital Course|7835,7839|false|false|false|||meal
Finding|Daily or Recreational Activity|Hospital Course|7835,7839|false|false|false|C1998602|Meal (occasion for eating)|meal
Finding|Intellectual Product|Hospital Course|7841,7847|false|false|false|C0034869|Records|Record
Event|Event|Hospital Course|7860,7864|false|false|false|||show
Event|Event|Hospital Course|7873,7883|false|false|false|||Oncologist
Anatomy|Body Location or Region|Hospital Course|7890,7894|false|false|false|C4318744|Test - temporal region|test
Finding|Functional Concept|Hospital Course|7890,7894|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|Hospital Course|7890,7894|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|Hospital Course|7890,7894|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|Hospital Course|7890,7894|false|false|false|C0022885|Laboratory Procedures|test
Event|Event|Hospital Course|7895,7901|false|false|false|||strips
Event|Event|Hospital Course|7907,7912|false|false|false|||Check
Disorder|Disease or Syndrome|Hospital Course|7913,7918|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Hospital Course|7913,7918|false|false|false|||blood
Finding|Body Substance|Hospital Course|7913,7918|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Organic Chemical|Hospital Course|7913,7925|false|false|false|C0005802|Blood Glucose|blood sugars
Drug|Organic Chemical|Hospital Course|7919,7925|false|false|false|C0242209|Sugars|sugars
Drug|Pharmacologic Substance|Hospital Course|7919,7925|false|false|false|C0242209|Sugars|sugars
Event|Event|Hospital Course|7919,7925|false|false|false|||sugars
Procedure|Laboratory Procedure|Hospital Course|7919,7925|false|false|false|C2239291|sugars (lab test)|sugars
Event|Event|Hospital Course|7932,7939|false|false|false|||refills
Finding|Idea or Concept|Hospital Course|7932,7939|false|false|false|C0807726|refill|refills
Event|Event|Hospital Course|7960,7965|false|false|false|||Check
Disorder|Disease or Syndrome|Hospital Course|7966,7971|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Hospital Course|7966,7971|false|false|false|||blood
Finding|Body Substance|Hospital Course|7966,7971|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Organic Chemical|Hospital Course|7966,7978|false|false|false|C0005802|Blood Glucose|blood sugars
Drug|Organic Chemical|Hospital Course|7972,7978|false|false|false|C0242209|Sugars|sugars
Drug|Pharmacologic Substance|Hospital Course|7972,7978|false|false|false|C0242209|Sugars|sugars
Event|Event|Hospital Course|7972,7978|false|false|false|||sugars
Procedure|Laboratory Procedure|Hospital Course|7972,7978|false|false|false|C2239291|sugars (lab test)|sugars
Event|Event|Hospital Course|7985,7992|false|false|false|||refills
Finding|Idea or Concept|Hospital Course|7985,7992|false|false|false|C0807726|refill|refills
Event|Event|Hospital Course|7998,8007|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|7998,8007|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|7998,8007|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|7998,8007|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|7998,8007|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|7998,8019|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|7998,8019|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|8008,8019|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|8008,8019|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|8008,8019|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|Hospital Course|8021,8025|false|false|false|||Home
Finding|Idea or Concept|Hospital Course|8021,8025|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|8021,8025|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|8021,8025|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|Hospital Course|8031,8038|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|Hospital Course|8031,8038|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|Hospital Course|8041,8049|false|false|false|||Facility
Finding|Intellectual Product|Hospital Course|8041,8049|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|Hospital Course|8057,8066|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|8057,8066|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|8057,8066|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|8057,8066|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|8057,8066|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|8057,8076|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|8067,8076|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|8067,8076|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|8067,8076|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|8067,8076|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|8067,8076|false|false|false|C0011900|Diagnosis|Diagnosis
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8078,8083|false|false|false|C0006104;C4266577|Brain;Head>Brain|Brain
Disorder|Disease or Syndrome|Hospital Course|8078,8083|false|false|false|C0006111|Brain Diseases|Brain
Disorder|Neoplastic Process|Hospital Course|8078,8089|false|false|false|C0006118|Brain Neoplasms|Brain tumor
Disorder|Neoplastic Process|Hospital Course|8084,8089|false|false|false|C0027651|Neoplasms|tumor
Event|Event|Hospital Course|8084,8089|false|false|false|||tumor
Finding|Finding|Hospital Course|8084,8089|false|false|false|C1578706;C3273930|Tumor Mass|tumor
Finding|Intellectual Product|Hospital Course|8084,8089|false|false|false|C1578706;C3273930|Tumor Mass|tumor
Finding|Mental Process|Discharge Condition|8114,8120|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|8114,8127|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|8114,8127|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|8121,8127|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|8121,8127|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|8129,8134|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|8129,8134|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|8139,8147|false|false|false|||coherent
Finding|Finding|Discharge Condition|8139,8147|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|8149,8154|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|8149,8171|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|8149,8171|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|8158,8171|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|8158,8171|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|8158,8171|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|8173,8178|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|8173,8178|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|8173,8178|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|8173,8178|false|false|false|||Alert
Finding|Finding|Discharge Condition|8173,8178|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|8173,8178|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|8173,8178|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|8183,8194|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|8183,8194|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|8196,8204|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|8196,8204|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|8196,8204|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|8205,8211|false|false|false|C5889824||Status
Event|Event|Discharge Condition|8205,8211|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|8205,8211|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|Discharge Condition|8213,8223|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|8213,8223|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|8213,8223|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|8213,8223|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|8226,8234|false|false|false|||requires
Event|Event|Discharge Condition|8235,8245|false|false|false|||assistance
Finding|Social Behavior|Discharge Condition|8235,8245|false|false|false|C0018896|Helping Behavior|assistance
Drug|Amino Acid, Peptide, or Protein|Discharge Condition|8249,8252|false|false|false|C1454018|AICDA protein, human|aid
Drug|Enzyme|Discharge Condition|8249,8252|false|false|false|C1454018|AICDA protein, human|aid
Event|Event|Discharge Condition|8249,8252|false|false|false|||aid
Finding|Gene or Genome|Discharge Condition|8249,8252|false|false|false|C1421876;C3540469|AICDA gene;AICDA wt Allele|aid
Procedure|Therapeutic or Preventive Procedure|Discharge Condition|8249,8252|false|false|false|C0021588;C0280108|AID - Artificial insemination by donor;dacarbazine/doxorubicin/ifosfamide protocol|aid
Finding|Finding|Discharge Instructions|8281,8288|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Finding|Functional Concept|Discharge Instructions|8281,8288|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Finding|Idea or Concept|Discharge Instructions|8281,8288|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|8281,8288|false|false|false|C0543467|Operative Surgical Procedures|Surgery
Event|Event|Discharge Instructions|8307,8314|false|false|false|||surgery
Finding|Finding|Discharge Instructions|8307,8314|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Discharge Instructions|8307,8314|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Discharge Instructions|8307,8314|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|8307,8314|false|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Event|Discharge Instructions|8318,8324|false|false|false|||remove
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|8327,8332|false|false|false|C0006104;C4266577|Brain;Head>Brain|brain
Disorder|Disease or Syndrome|Discharge Instructions|8327,8332|false|false|false|C0006111|Brain Diseases|brain
Finding|Finding|Discharge Instructions|8327,8339|false|false|false|C0221505|Lesion of brain|brain lesion
Event|Event|Discharge Instructions|8333,8339|false|false|false|||lesion
Finding|Finding|Discharge Instructions|8333,8339|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|Discharge Instructions|8333,8339|false|false|false|C0221198;C1546698|Lesion|lesion
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|8351,8356|false|false|false|C0006104;C4266577|Brain;Head>Brain|brain
Disorder|Disease or Syndrome|Discharge Instructions|8351,8356|false|false|false|C0006111|Brain Diseases|brain
Event|Event|Discharge Instructions|8351,8356|false|false|false|||brain
Drug|Substance|Discharge Instructions|8364,8370|false|false|false|C0370003|Specimen|sample
Event|Event|Discharge Instructions|8364,8370|false|false|false|||sample
Finding|Body Substance|Discharge Instructions|8364,8370|false|false|false|C2347026;C5551027|Biospecimen;Nucleotide Sequence Sample Name|sample
Finding|Intellectual Product|Discharge Instructions|8364,8370|false|false|false|C2347026;C5551027|Biospecimen;Nucleotide Sequence Sample Name|sample
Anatomy|Tissue|Discharge Instructions|8374,8380|false|false|false|C0040300|Body tissue|tissue
Finding|Intellectual Product|Discharge Instructions|8374,8380|false|false|false|C1547928|Tissue Specimen Code|tissue
Event|Event|Discharge Instructions|8390,8396|false|false|false|||lesion
Finding|Finding|Discharge Instructions|8390,8396|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|Discharge Instructions|8390,8396|false|false|false|C0221198;C1546698|Lesion|lesion
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|8405,8410|false|false|false|C0006104;C4266577|Brain;Head>Brain|brain
Disorder|Disease or Syndrome|Discharge Instructions|8405,8410|false|false|false|C0006111|Brain Diseases|brain
Event|Event|Discharge Instructions|8415,8419|false|false|false|||sent
Event|Event|Discharge Instructions|8424,8433|false|false|false|||pathology
Finding|Functional Concept|Discharge Instructions|8424,8433|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Finding|Pathologic Function|Discharge Instructions|8424,8433|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Procedure|Laboratory Procedure|Discharge Instructions|8424,8433|false|false|false|C0919386|Pathology procedure|pathology
Event|Event|Discharge Instructions|8438,8445|false|false|false|||testing
Finding|Functional Concept|Discharge Instructions|8438,8445|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|testing
Finding|Intellectual Product|Discharge Instructions|8438,8445|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|testing
Event|Event|Discharge Instructions|8458,8462|false|false|false|||keep
Anatomy|Body Location or Region|Discharge Instructions|8468,8476|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Discharge Instructions|8468,8476|false|false|false|C0332803|Surgical wound|incision
Event|Event|Discharge Instructions|8468,8476|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|8468,8476|false|false|false|C0184898|Surgical incisions|incision
Anatomy|Body Space or Junction|Discharge Instructions|8492,8499|false|false|false|C0502420|Suture Joint|sutures
Event|Event|Discharge Instructions|8492,8499|false|false|false|||sutures
Event|Event|Discharge Instructions|8504,8511|false|false|false|||removed
Event|Event|Discharge Instructions|8525,8531|false|false|false|||shower
Finding|Finding|Discharge Instructions|8540,8544|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Discharge Instructions|8540,8544|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Discharge Instructions|8540,8544|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Anatomy|Body Location or Region|Discharge Instructions|8559,8567|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Discharge Instructions|8559,8567|false|false|false|C0332803|Surgical wound|incision
Event|Event|Discharge Instructions|8559,8567|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|8559,8567|false|false|false|C0184898|Surgical incisions|incision
Disorder|Disease or Syndrome|Discharge Instructions|8582,8586|false|false|false|C0339510|Vitelliform Macular Dystrophy|best
Event|Event|Discharge Instructions|8582,8586|false|false|false|||best
Finding|Gene or Genome|Discharge Instructions|8582,8586|false|false|false|C1826421;C5781213|BEST1 gene;BEST1 wt Allele|best
Event|Event|Discharge Instructions|8590,8594|false|false|false|||keep
Anatomy|Body Location or Region|Discharge Instructions|8600,8608|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Discharge Instructions|8600,8608|false|false|false|C0332803|Surgical wound|incision
Event|Event|Discharge Instructions|8600,8608|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|8600,8608|false|false|false|C0184898|Surgical incisions|incision
Event|Event|Discharge Instructions|8609,8613|false|false|false|||open
Drug|Inorganic Chemical|Discharge Instructions|8617,8620|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|Discharge Instructions|8617,8620|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|Discharge Instructions|8617,8620|false|false|false|C0001861;C3536832|Air (substance);air|air
Event|Event|Discharge Instructions|8617,8620|false|false|false|||air
Finding|Finding|Discharge Instructions|8617,8620|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|Discharge Instructions|8617,8620|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|Discharge Instructions|8617,8620|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Event|Event|Discharge Instructions|8638,8643|false|false|false|||cover
Event|Event|Discharge Instructions|8665,8669|false|false|false|||Call
Finding|Functional Concept|Discharge Instructions|8665,8669|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|Call
Finding|Gene or Genome|Discharge Instructions|8665,8669|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|Call
Finding|Intellectual Product|Discharge Instructions|8665,8669|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|Call
Finding|Mental Process|Discharge Instructions|8665,8669|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|Call
Attribute|Clinical Attribute|Discharge Instructions|8675,8682|false|false|false|C5444295||surgeon
Event|Event|Discharge Instructions|8700,8705|true|false|false|||signs
Finding|Finding|Discharge Instructions|8700,8705|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Discharge Instructions|8700,8705|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Disorder|Disease or Syndrome|Discharge Instructions|8709,8718|true|false|false|C0009450|Communicable Diseases|infection
Event|Event|Discharge Instructions|8709,8718|true|false|false|||infection
Finding|Pathologic Function|Discharge Instructions|8709,8718|true|false|false|C3714514|Infection|infection
Disorder|Disease or Syndrome|Discharge Instructions|8725,8732|true|false|false|C0041834|Erythema|redness
Event|Event|Discharge Instructions|8725,8732|true|false|false|||redness
Finding|Finding|Discharge Instructions|8725,8732|true|false|false|C0332575|Redness|redness
Event|Event|Discharge Instructions|8734,8739|false|false|false|||fever
Finding|Finding|Discharge Instructions|8734,8739|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|Discharge Instructions|8734,8739|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|Discharge Instructions|8744,8752|false|false|false|||drainage
Finding|Body Substance|Discharge Instructions|8744,8752|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|Discharge Instructions|8744,8752|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|8744,8752|false|false|false|C0013103|Drainage procedure|drainage
Event|Activity|Discharge Instructions|8756,8764|false|false|false|C0441655|Activities|Activity
Event|Event|Discharge Instructions|8756,8764|false|false|false|||Activity
Finding|Daily or Recreational Activity|Discharge Instructions|8756,8764|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Instructions|8756,8764|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Event|Event|Discharge Instructions|8772,8781|false|false|false|||recommend
Event|Event|Discharge Instructions|8791,8796|false|false|false|||avoid
Event|Activity|Discharge Instructions|8803,8810|false|false|false|C0206244|Lifting|lifting
Event|Event|Discharge Instructions|8803,8810|false|false|false|||lifting
Event|Event|Discharge Instructions|8812,8819|false|false|false|||running
Finding|Daily or Recreational Activity|Discharge Instructions|8812,8819|false|false|false|C0035953;C2346414;C4722187|Go Jogging or Running Question;Running (physical activity);running (history)|running
Finding|Finding|Discharge Instructions|8812,8819|false|false|false|C0035953;C2346414;C4722187|Go Jogging or Running Question;Running (physical activity);running (history)|running
Finding|Intellectual Product|Discharge Instructions|8812,8819|false|false|false|C0035953;C2346414;C4722187|Go Jogging or Running Question;Running (physical activity);running (history)|running
Event|Event|Discharge Instructions|8821,8829|false|false|false|||climbing
Finding|Finding|Discharge Instructions|8821,8829|false|false|false|C0561942;C2362653;C2584300|Climbing;Does climb;climbing (history)|climbing
Finding|Individual Behavior|Discharge Instructions|8821,8829|false|false|false|C0561942;C2362653;C2584300|Climbing;Does climb;climbing (history)|climbing
Finding|Daily or Recreational Activity|Discharge Instructions|8841,8859|false|false|false|C1514989|Strenuous Exercise|strenuous exercise
Event|Event|Discharge Instructions|8851,8859|false|false|false|||exercise
Finding|Daily or Recreational Activity|Discharge Instructions|8851,8859|false|false|false|C0015259|Exercise|exercise
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|8851,8859|false|false|false|C1522704|Exercise Pain Management|exercise
Event|Event|Discharge Instructions|8871,8877|false|false|false|||follow
Finding|Functional Concept|Discharge Instructions|8871,8877|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|Discharge Instructions|8871,8877|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|Discharge Instructions|8871,8880|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|Discharge Instructions|8871,8880|false|false|false|C1522577|follow-up|follow-up
Event|Activity|Discharge Instructions|8881,8892|false|false|false|C0003629|Appointments|appointment
Event|Event|Discharge Instructions|8881,8892|false|false|false|||appointment
Event|Event|Discharge Instructions|8921,8926|false|false|false|||walks
Finding|Finding|Discharge Instructions|8921,8926|false|false|false|C0600108|Does walk|walks
Event|Event|Discharge Instructions|8938,8946|false|false|false|||increase
Event|Activity|Discharge Instructions|8953,8961|false|false|false|C0441655|Activities|activity
Event|Event|Discharge Instructions|8953,8961|false|false|false|||activity
Finding|Daily or Recreational Activity|Discharge Instructions|8953,8961|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Finding|Finding|Discharge Instructions|8953,8961|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Finding|Finding|Discharge Instructions|8970,8973|false|false|false|C5939094|Own|own
Drug|Amino Acid, Peptide, or Protein|Discharge Instructions|8974,8978|false|false|false|C0281567;C1310542;C4048252|FURIN protein, human;cisplatin/cyclophosphamide/doxorubicin/etoposide;cyclophosphamide/doxorubicin/etoposide/prednisone|pace
Drug|Enzyme|Discharge Instructions|8974,8978|false|false|false|C0281567;C1310542;C4048252|FURIN protein, human;cisplatin/cyclophosphamide/doxorubicin/etoposide;cyclophosphamide/doxorubicin/etoposide/prednisone|pace
Drug|Pharmacologic Substance|Discharge Instructions|8974,8978|false|false|false|C0281567;C1310542;C4048252|FURIN protein, human;cisplatin/cyclophosphamide/doxorubicin/etoposide;cyclophosphamide/doxorubicin/etoposide/prednisone|pace
Event|Event|Discharge Instructions|8974,8978|false|false|false|||pace
Finding|Gene or Genome|Discharge Instructions|8974,8978|false|false|false|C0919550;C1150256;C5444037|FURIN gene;Patient Assessment of Cancer Communication Experiences;furin activity|pace
Finding|Intellectual Product|Discharge Instructions|8974,8978|false|false|false|C0919550;C1150256;C5444037|FURIN gene;Patient Assessment of Cancer Communication Experiences;furin activity|pace
Finding|Molecular Function|Discharge Instructions|8974,8978|false|false|false|C0919550;C1150256;C5444037|FURIN gene;Patient Assessment of Cancer Communication Experiences;furin activity|pace
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|8974,8978|false|false|false|C0280022|cisplatin/cyclophosphamide/doxorubicin/vindesine protocol|pace
Attribute|Clinical Attribute|Discharge Instructions|8992,8999|false|false|false|C3854129||symptom
Event|Event|Discharge Instructions|8992,8999|false|false|false|||symptom
Finding|Sign or Symptom|Discharge Instructions|8992,8999|false|false|false|C1457887|Symptoms|symptom
Event|Event|Discharge Instructions|9000,9004|false|false|false|||free
Finding|Functional Concept|Discharge Instructions|9000,9004|false|false|false|C0332296|Free of (attribute)|free
Finding|Functional Concept|Discharge Instructions|9005,9012|false|false|false|C0443144|At rest (qualifier value)|at rest
Drug|Amino Acid, Peptide, or Protein|Discharge Instructions|9008,9012|false|false|false|C1742913|REST protein, human|rest
Drug|Biologically Active Substance|Discharge Instructions|9008,9012|false|false|false|C1742913|REST protein, human|rest
Event|Event|Discharge Instructions|9008,9012|false|false|false|||rest
Finding|Daily or Recreational Activity|Discharge Instructions|9008,9012|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Gene or Genome|Discharge Instructions|9008,9012|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Molecular Function|Discharge Instructions|9008,9012|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Finding|Discharge Instructions|9029,9037|false|false|false|C3843660|Too much|too much
Finding|Finding|Discharge Instructions|9033,9037|false|false|false|C4281574|Much|much
Finding|Intellectual Product|Discharge Instructions|9045,9049|false|false|false|C1720092|Once - dosing instruction fragment|once
Event|Event|Discharge Instructions|9057,9064|true|false|false|||driving
Finding|Daily or Recreational Activity|Discharge Instructions|9057,9064|true|false|false|C0004379|Automobile Driving|driving
Event|Event|Discharge Instructions|9071,9077|true|false|false|||taking
Drug|Hazardous or Poisonous Substance|Discharge Instructions|9082,9090|true|false|false|C0027415|Narcotics|narcotic
Drug|Pharmacologic Substance|Discharge Instructions|9082,9090|true|false|false|C0027415|Narcotics|narcotic
Event|Event|Discharge Instructions|9082,9090|true|false|false|||narcotic
Event|Event|Discharge Instructions|9094,9102|true|false|false|||sedating
Drug|Pharmacologic Substance|Discharge Instructions|9103,9113|true|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Discharge Instructions|9103,9113|true|false|false|||medication
Finding|Intellectual Product|Discharge Instructions|9103,9113|true|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Discharge Instructions|9140,9147|false|false|false|||seizure
Finding|Sign or Symptom|Discharge Instructions|9140,9147|false|false|false|C0036572|Seizures|seizure
Event|Event|Discharge Instructions|9154,9162|true|false|false|||admitted
Event|Event|Discharge Instructions|9177,9184|true|false|false|||allowed
Event|Event|Discharge Instructions|9188,9193|true|false|false|||drive
Finding|Intellectual Product|Discharge Instructions|9197,9200|true|false|false|C1947938|Law (document)|law
Event|Activity|Discharge Instructions|9209,9216|true|false|false|C3812666|Personal Contact|contact
Finding|Functional Concept|Discharge Instructions|9209,9216|true|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|contact
Finding|Idea or Concept|Discharge Instructions|9209,9216|true|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|contact
Finding|Intellectual Product|Discharge Instructions|9209,9216|true|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|contact
Phenomenon|Phenomenon or Process|Discharge Instructions|9209,9216|true|false|false|C0392367|Physical contact|contact
Event|Event|Discharge Instructions|9217,9223|true|false|false|||sports
Finding|Daily or Recreational Activity|Discharge Instructions|9217,9223|true|false|false|C0038039|Sports|sports
Event|Event|Discharge Instructions|9230,9237|true|false|false|||cleared
Event|Event|Discharge Instructions|9246,9258|true|false|false|||neurosurgeon
Event|Activity|Discharge Instructions|9278,9285|false|false|false|C3812666|Personal Contact|contact
Event|Event|Discharge Instructions|9278,9285|false|false|false|||contact
Finding|Functional Concept|Discharge Instructions|9278,9285|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|contact
Finding|Idea or Concept|Discharge Instructions|9278,9285|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|contact
Finding|Intellectual Product|Discharge Instructions|9278,9285|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|contact
Phenomenon|Phenomenon or Process|Discharge Instructions|9278,9285|false|false|false|C0392367|Physical contact|contact
Event|Event|Discharge Instructions|9286,9292|false|false|false|||sports
Finding|Daily or Recreational Activity|Discharge Instructions|9286,9292|false|false|false|C0038039|Sports|sports
Event|Event|Medications|9339,9343|true|false|false|||take
Disorder|Disease or Syndrome|Medications|9348,9353|true|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Medications|9348,9353|true|false|false|||blood
Finding|Body Substance|Medications|9348,9353|true|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Sign or Symptom|Medications|9354,9362|true|false|false|C0851184|Thinning Weight Loss|thinning
Drug|Pharmacologic Substance|Medications|9363,9373|true|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Medications|9363,9373|true|false|false|||medication
Finding|Intellectual Product|Medications|9363,9373|true|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Drug|Organic Chemical|Medications|9375,9382|true|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Medications|9375,9382|true|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|Medications|9385,9394|false|false|false|C0020740|ibuprofen|Ibuprofen
Drug|Pharmacologic Substance|Medications|9385,9394|false|false|false|C0020740|ibuprofen|Ibuprofen
Event|Event|Medications|9385,9394|false|false|false|||Ibuprofen
Drug|Organic Chemical|Medications|9396,9402|false|false|false|C0633084|Plavix|Plavix
Drug|Pharmacologic Substance|Medications|9396,9402|false|false|false|C0633084|Plavix|Plavix
Event|Event|Medications|9396,9402|false|false|false|||Plavix
Drug|Organic Chemical|Medications|9404,9412|false|false|false|C0699129|Coumadin|Coumadin
Drug|Pharmacologic Substance|Medications|9404,9412|false|false|false|C0699129|Coumadin|Coumadin
Event|Event|Medications|9404,9412|false|false|false|||Coumadin
Event|Event|Medications|9420,9427|false|false|false|||cleared
Event|Event|Medications|9453,9457|false|false|false|||held
Drug|Organic Chemical|Medications|9463,9470|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Medications|9463,9470|false|false|false|C0004057|aspirin|Aspirin
Event|Event|Medications|9491,9498|false|false|false|||cleared
Event|Event|Medications|9502,9508|false|false|false|||resume
Drug|Pharmacologic Substance|Medications|9515,9525|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Medications|9515,9525|false|false|false|||medication
Finding|Intellectual Product|Medications|9515,9525|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Medications|9529,9532|false|false|false|||POD
Event|Event|Medications|9550,9554|false|false|false|||held
Finding|Idea or Concept|Medications|9560,9564|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Medications|9560,9564|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Medications|9560,9564|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Medications|9565,9576|false|false|false|C0102118|alendronate|Alendronate
Drug|Pharmacologic Substance|Medications|9565,9576|false|false|false|C0102118|alendronate|Alendronate
Event|Event|Medications|9565,9576|false|false|false|||Alendronate
Event|Event|Medications|9589,9598|false|false|false|||admission
Procedure|Health Care Activity|Medications|9589,9598|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|Medications|9609,9616|false|false|false|||cleared
Event|Event|Medications|9620,9626|false|false|false|||resume
Drug|Pharmacologic Substance|Medications|9632,9642|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Medications|9632,9642|false|false|false|||medication
Finding|Intellectual Product|Medications|9632,9642|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Medications|9646,9649|false|false|false|||POD
Event|Event|Medications|9672,9675|false|false|false|||use
Drug|Organic Chemical|Medications|9676,9689|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Medications|9676,9689|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Medications|9676,9689|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Medications|9676,9689|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Organic Chemical|Medications|9691,9698|false|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|Medications|9691,9698|false|false|false|C0699142|Tylenol|Tylenol
Disorder|Disease or Syndrome|Medications|9704,9709|false|false|false|C1446899|minor (disease)|minor
Event|Event|Medications|9704,9709|false|false|false|||minor
Finding|Gene or Genome|Medications|9704,9709|false|false|false|C1417837;C3272493|NR4A3 gene;NR4A3 wt Allele|minor
Event|Event|Medications|9710,9720|false|false|false|||discomfort
Finding|Sign or Symptom|Medications|9710,9720|false|false|false|C2364135|Discomfort|discomfort
Event|Event|Medications|9747,9757|true|false|false|||restricted
Event|Event|Medications|9763,9769|true|false|false|||taking
Drug|Pharmacologic Substance|Medications|9775,9785|true|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Medications|9775,9785|true|false|false|||medication
Finding|Intellectual Product|Medications|9775,9785|true|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Medications|9799,9806|false|false|false|||started
Drug|Organic Chemical|Medications|9810,9823|false|false|false|C0011777|dexamethasone|Dexamethasone
Drug|Pharmacologic Substance|Medications|9810,9823|false|false|false|C0011777|dexamethasone|Dexamethasone
Event|Event|Medications|9810,9823|false|false|false|||Dexamethasone
Drug|Organic Chemical|Medications|9827,9834|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Drug|Pharmacologic Substance|Medications|9827,9834|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Event|Event|Medications|9827,9834|false|false|false|||steroid
Event|Event|Medications|9840,9846|false|false|false|||treats
Finding|Functional Concept|Medications|9840,9846|false|false|false|C1292734;C5966192|Intent To Treat;Treats (attribute)|treats
Anatomy|Body Location or Region|Medications|9848,9860|false|false|false|C0524466|Intracranial|intracranial
Finding|Functional Concept|Medications|9848,9860|false|false|false|C1522213|Intracranial Route of Administration|intracranial
Finding|Pathologic Function|Medications|9848,9869|false|false|false|C1527311|Brain Edema|intracranial swelling
Event|Event|Medications|9861,9869|false|false|false|||swelling
Finding|Finding|Medications|9861,9869|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|Medications|9861,9869|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Drug|Organic Chemical|Medications|9876,9889|false|false|false|C0011777|dexamethasone|Dexamethasone
Drug|Pharmacologic Substance|Medications|9876,9889|false|false|false|C0011777|dexamethasone|Dexamethasone
Event|Event|Medications|9876,9889|false|false|false|||Dexamethasone
Event|Event|Medications|9899,9906|false|false|false|||tapered
Event|Activity|Medications|9918,9929|false|false|false|C0024501|Maintenance|maintenance
Event|Event|Medications|9930,9934|false|false|false|||dose
Disorder|Mental or Behavioral Dysfunction|Medications|9942,9945|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Medications|9942,9945|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Medications|9942,9945|false|false|false|C1530795|BID protein, human|BID
Event|Event|Medications|9942,9945|false|false|false|||BID
Finding|Gene or Genome|Medications|9942,9945|false|false|false|C1332410|BID gene|BID
Event|Event|Medications|9954,9958|false|false|false|||take
Drug|Pharmacologic Substance|Medications|9964,9974|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Medications|9964,9974|false|false|false|||medication
Finding|Intellectual Product|Medications|9964,9974|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Medications|9979,9989|false|false|false|||prescribed
Event|Event|Medications|10000,10008|false|false|false|||admitted
Disorder|Disease or Syndrome|Medications|10018,10040|false|false|false|C0020456|Hyperglycemia|elevated blood glucose
Finding|Finding|Medications|10018,10040|false|false|false|C0595877;C2703060|Blood glucose increased;elevated random blood glucose level|elevated blood glucose
Disorder|Disease or Syndrome|Medications|10027,10032|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Medications|10027,10032|false|false|false|||blood
Finding|Body Substance|Medications|10027,10032|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Organic Chemical|Medications|10027,10040|false|false|false|C0005802|Blood Glucose|blood glucose
Lab|Laboratory or Test Result|Medications|10027,10040|false|false|false|C0428554|Finding of blood glucose level|blood glucose
Procedure|Laboratory Procedure|Medications|10027,10040|false|false|false|C0392201|Blood glucose measurement|blood glucose
Lab|Laboratory or Test Result|Medications|10027,10047|false|false|false|C0428554|Finding of blood glucose level|blood glucose levels
Drug|Biologically Active Substance|Medications|10033,10040|false|false|false|C0017725|glucose|glucose
Drug|Organic Chemical|Medications|10033,10040|false|false|false|C0017725|glucose|glucose
Drug|Pharmacologic Substance|Medications|10033,10040|false|false|false|C0017725|glucose|glucose
Event|Event|Medications|10033,10040|false|false|false|||glucose
Lab|Laboratory or Test Result|Medications|10033,10040|false|false|false|C5781949|Glucose^1.5H post dose glucagon|glucose
Procedure|Laboratory Procedure|Medications|10033,10040|false|false|false|C0337438|Glucose measurement|glucose
Lab|Laboratory or Test Result|Medications|10033,10047|false|false|false|C0428548||glucose levels
Event|Event|Medications|10041,10047|false|false|false|||levels
Event|Event|Medications|10054,10060|false|false|false|||needed
Event|Event|Medications|10067,10074|false|false|false|||treated
Drug|Amino Acid, Peptide, or Protein|Medications|10078,10085|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Hormone|Medications|10078,10085|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Pharmacologic Substance|Medications|10078,10085|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Event|Event|Medications|10078,10085|false|false|false|||Insulin
Finding|Gene or Genome|Medications|10078,10085|false|false|false|C1337112|INS gene|Insulin
Procedure|Laboratory Procedure|Medications|10078,10085|false|false|false|C0202098|Insulin measurement|Insulin
Event|Event|Medications|10098,10106|false|false|false|||continue
Event|Activity|Medications|10110,10115|false|false|false|C1283174||check
Event|Event|Medications|10110,10115|false|false|false|||check
Finding|Functional Concept|Medications|10110,10115|false|false|false|C4321547|Check|check
Disorder|Disease or Syndrome|Medications|10122,10127|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Medications|10122,10127|false|false|false|||blood
Finding|Body Substance|Medications|10122,10127|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Organic Chemical|Medications|10122,10134|false|false|false|C0005802|Blood Glucose|blood sugars
Drug|Organic Chemical|Medications|10128,10134|false|false|false|C0242209|Sugars|sugars
Drug|Pharmacologic Substance|Medications|10128,10134|false|false|false|C0242209|Sugars|sugars
Event|Event|Medications|10128,10134|false|false|false|||sugars
Procedure|Laboratory Procedure|Medications|10128,10134|false|false|false|C2239291|sugars (lab test)|sugars
Finding|Finding|Medications|10141,10148|false|false|false|C4534363|At home|at home
Event|Event|Medications|10144,10148|false|false|false|||home
Finding|Idea or Concept|Medications|10144,10148|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Medications|10144,10148|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Medications|10144,10148|false|false|false|C1553498|home health encounter|home
Event|Event|Medications|10169,10179|false|false|false|||glucometer
Event|Event|Medications|10208,10213|false|false|false|||teach
Event|Event|Medications|10225,10228|false|false|false|||use
Event|Event|Medications|10234,10240|false|false|false|||device
Finding|Functional Concept|Medications|10234,10240|false|false|false|C1550509|Participation Type - device|device
Event|Event|Medications|10245,10249|false|false|false|||home
Finding|Idea or Concept|Medications|10245,10249|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Medications|10245,10249|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Medications|10245,10249|false|false|false|C1553498|home health encounter|home
Event|Event|Medications|10258,10264|false|false|false|||record
Disorder|Disease or Syndrome|Medications|10270,10275|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Medications|10270,10275|false|false|false|||blood
Finding|Body Substance|Medications|10270,10275|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Organic Chemical|Medications|10270,10282|false|false|false|C0005802|Blood Glucose|blood sugars
Drug|Organic Chemical|Medications|10276,10282|false|false|false|C0242209|Sugars|sugars
Drug|Pharmacologic Substance|Medications|10276,10282|false|false|false|C0242209|Sugars|sugars
Event|Event|Medications|10276,10282|false|false|false|||sugars
Procedure|Laboratory Procedure|Medications|10276,10282|false|false|false|C2239291|sugars (lab test)|sugars
Event|Event|Medications|10287,10293|false|false|false|||follow
Disorder|Disease or Syndrome|Medications|10308,10311|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|Medications|10308,10311|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|Medications|10308,10311|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|Medications|10308,10311|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|Medications|10308,10311|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|Medications|10308,10311|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|Medications|10308,10311|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|Medications|10308,10311|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|Medications|10308,10311|false|false|false|||PCP
Finding|Gene or Genome|Medications|10308,10311|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|Medications|10308,10311|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|Medications|10348,10352|false|false|false|||goal
Finding|Idea or Concept|Medications|10348,10352|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Finding|Intellectual Product|Medications|10348,10352|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Disorder|Disease or Syndrome|Medications|10353,10358|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Medications|10353,10358|false|false|false|||blood
Finding|Body Substance|Medications|10353,10358|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Organic Chemical|Medications|10353,10364|false|false|false|C0005802|Blood Glucose|blood sugar
Procedure|Laboratory Procedure|Medications|10353,10364|false|false|false|C0392201|Blood glucose measurement|blood sugar
Drug|Biomedical or Dental Material|Medications|10359,10364|false|false|false|C0007004;C0242209;C3665462|Carbohydrates;Sugars;raw sugar|sugar
Drug|Organic Chemical|Medications|10359,10364|false|false|false|C0007004;C0242209;C3665462|Carbohydrates;Sugars;raw sugar|sugar
Drug|Pharmacologic Substance|Medications|10359,10364|false|false|false|C0007004;C0242209;C3665462|Carbohydrates;Sugars;raw sugar|sugar
Event|Event|Medications|10359,10364|false|false|false|||sugar
Finding|Mental Process|Medications|10399,10409|false|false|false|C0237607;C0596545|Experience;Experience (Practice)|Experience
Event|Event|Medications|10433,10442|false|false|false|||headaches
Finding|Sign or Symptom|Medications|10433,10442|false|false|false|C0018681|Headache|headaches
Procedure|Therapeutic or Preventive Procedure|Medications|10447,10457|false|false|false|C0184898|Surgical incisions|incisional
Finding|Sign or Symptom|Medications|10447,10462|false|false|false|C1717947|Incisional pain|incisional pain
Attribute|Clinical Attribute|Medications|10458,10462|false|false|false|C2598155||pain
Event|Event|Medications|10458,10462|false|false|false|||pain
Finding|Functional Concept|Medications|10458,10462|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Medications|10458,10462|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Medications|10481,10491|false|false|false|||experience
Finding|Finding|Medications|10512,10520|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|Medications|10512,10520|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Event|Event|Medications|10521,10527|false|false|false|||around
Anatomy|Body Location or Region|Medications|10534,10538|false|false|false|C0015450;C4266571|Face;Head>Face|face
Disorder|Disease or Syndrome|Medications|10534,10538|false|false|false|C3160739|FANCONI ANEMIA, COMPLEMENTATION GROUP E|face
Event|Event|Medications|10534,10538|false|false|false|||face
Finding|Gene or Genome|Medications|10534,10538|false|false|false|C1414531;C1423759;C2828055|ELOVL6 gene;FANCE gene;FANCE wt Allele|face
Anatomy|Body Part, Organ, or Organ Component|Medications|10543,10547|false|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|Medications|10543,10547|false|false|false|C5848506||eyes
Event|Event|Medications|10557,10563|false|false|false|||normal
Finding|Finding|Medications|10564,10577|false|false|false|C0241311|post operative (finding)|after surgery
Event|Event|Medications|10570,10577|false|false|false|||surgery
Finding|Finding|Medications|10570,10577|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Medications|10570,10577|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Medications|10570,10577|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Medications|10570,10577|false|false|false|C0543467|Operative Surgical Procedures|surgery
Finding|Functional Concept|Medications|10606,10612|false|false|false|C1522484;C1561503;C1705190|Precision - second;Second Suffix;metastatic qualifier|second
Finding|Idea or Concept|Medications|10606,10612|false|false|false|C1522484;C1561503;C1705190|Precision - second;Second Suffix;metastatic qualifier|second
Finding|Intellectual Product|Medications|10606,10612|false|false|false|C1522484;C1561503;C1705190|Precision - second;Second Suffix;metastatic qualifier|second
Finding|Idea or Concept|Medications|10623,10626|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Medications|10623,10626|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Medications|10630,10637|false|false|false|||surgery
Finding|Finding|Medications|10630,10637|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Medications|10630,10637|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Medications|10630,10637|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Medications|10630,10637|false|false|false|C0543467|Operative Surgical Procedures|surgery
Finding|Functional Concept|Medications|10644,10649|false|false|false|C1632850;C1879355;C4048755;C4521676|Apply;Apply (administration method);Apply (instruction)|apply
Anatomy|Body Part, Organ, or Organ Component|Medications|10651,10654|false|false|false|C0228434;C3496566|Structure of inferior central nucleus of pons;intracentral fissure|ice
Anatomy|Body Space or Junction|Medications|10651,10654|false|false|false|C0228434;C3496566|Structure of inferior central nucleus of pons;intracentral fissure|ice
Drug|Amino Acid, Peptide, or Protein|Medications|10651,10654|false|false|false|C0020746;C0025611;C1873773;C4721557|Caspase-1, human;Ice;Ice Pharmaceutical;methamphetamine|ice
Drug|Enzyme|Medications|10651,10654|false|false|false|C0020746;C0025611;C1873773;C4721557|Caspase-1, human;Ice;Ice Pharmaceutical;methamphetamine|ice
Drug|Hazardous or Poisonous Substance|Medications|10651,10654|false|false|false|C0020746;C0025611;C1873773;C4721557|Caspase-1, human;Ice;Ice Pharmaceutical;methamphetamine|ice
Drug|Inorganic Chemical|Medications|10651,10654|false|false|false|C0020746;C0025611;C1873773;C4721557|Caspase-1, human;Ice;Ice Pharmaceutical;methamphetamine|ice
Drug|Organic Chemical|Medications|10651,10654|false|false|false|C0020746;C0025611;C1873773;C4721557|Caspase-1, human;Ice;Ice Pharmaceutical;methamphetamine|ice
Drug|Pharmacologic Substance|Medications|10651,10654|false|false|false|C0020746;C0025611;C1873773;C4721557|Caspase-1, human;Ice;Ice Pharmaceutical;methamphetamine|ice
Event|Event|Medications|10651,10654|false|false|false|||ice
Finding|Gene or Genome|Medications|10651,10654|false|false|false|C1150137;C1366479;C1413348;C1705786;C3889432|CASP1 gene;CASP1 wt Allele;CES2 gene;CES2 wt Allele;caspase-1 activity|ice
Finding|Molecular Function|Medications|10651,10654|false|false|false|C1150137;C1366479;C1413348;C1705786;C3889432|CASP1 gene;CASP1 wt Allele;CES2 gene;CES2 wt Allele;caspase-1 activity|ice
Procedure|Therapeutic or Preventive Procedure|Medications|10651,10654|false|false|false|C0249492;C0280697;C0556917;C1879508|AIE Regimen;carboplatin/etoposide/ifosfamide;cryotherapy using ice;cytarabine/etoposide/idarubicin|ice
Phenomenon|Natural Phenomenon or Process|Medications|10660,10664|false|false|false|C0678568||cool
Event|Event|Medications|10668,10672|false|false|false|||warm
Finding|Finding|Medications|10668,10672|false|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|Medications|10668,10672|false|false|false|C0687712|warming process|warm
Anatomy|Body Part, Organ, or Organ Component|Medications|10691,10695|false|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|Medications|10691,10695|false|false|false|C5848506||eyes
Event|Event|Medications|10699,10703|false|false|false|||help
Event|Event|Medications|10714,10722|false|false|false|||swelling
Finding|Finding|Medications|10714,10722|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|Medications|10714,10722|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Event|Event|Medications|10728,10736|false|false|false|||swelling
Finding|Finding|Medications|10728,10736|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|Medications|10728,10736|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Event|Event|Medications|10749,10754|false|false|false|||worse
Finding|Finding|Medications|10749,10754|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Idea or Concept|Medications|10749,10754|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Drug|Organic Chemical|Medications|10762,10775|false|false|false|C4019028|Morning After|morning after
Drug|Pharmacologic Substance|Medications|10762,10775|false|false|false|C4019028|Morning After|morning after
Event|Event|Medications|10770,10775|false|false|false|||after
Event|Event|Medications|10777,10783|false|false|false|||laying
Event|Event|Medications|10794,10802|false|false|false|||sleeping
Event|Event|Medications|10807,10815|false|false|false|||decrease
Event|Event|Medications|10837,10847|false|false|false|||experience
Event|Event|Medications|10848,10856|false|false|false|||soreness
Finding|Sign or Symptom|Medications|10848,10856|false|false|false|C0234233|Sore to touch|soreness
Event|Event|Medications|10862,10869|false|false|false|||chewing
Finding|Finding|Medications|10862,10869|false|false|false|C0024888;C2015927|Chewing;outcomes otolaryngology chewing|chewing
Finding|Organism Function|Medications|10862,10869|false|false|false|C0024888;C2015927|Chewing;outcomes otolaryngology chewing|chewing
Event|Event|Medications|10879,10885|false|false|false|||normal
Event|Event|Medications|10896,10903|false|false|false|||surgery
Finding|Finding|Medications|10896,10903|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Medications|10896,10903|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Medications|10896,10903|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Medications|10896,10903|false|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Event|Medications|10913,10920|false|false|false|||improve
Finding|Finding|Medications|10926,10930|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Medications|10926,10930|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Medications|10926,10930|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Drug|Food|Medications|10939,10944|false|false|false|C0016452|Food|foods
Event|Event|Medications|10939,10944|false|false|false|||foods
Finding|Finding|Medications|10972,10976|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Medications|10972,10976|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Medications|10972,10976|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|Medications|10995,11000|false|false|false|||tired
Finding|Finding|Medications|10995,11000|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Finding|Intellectual Product|Medications|10995,11000|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Finding|Sign or Symptom|Medications|10995,11000|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Event|Event|Medications|11004,11016|false|false|false|||restlessness
Finding|Finding|Medications|11004,11016|false|false|false|C0085631;C3887611;C3887612|Agitation;Psychomotor Agitation;Restlessness|restlessness
Finding|Sign or Symptom|Medications|11004,11016|false|false|false|C0085631;C3887611;C3887612|Agitation;Psychomotor Agitation;Restlessness|restlessness
Event|Event|Medications|11025,11031|false|false|false|||common
Finding|Functional Concept|Medications|11025,11031|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Finding|Intellectual Product|Medications|11025,11031|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Event|Event|Medications|11036,11048|false|false|false|||Constipation
Finding|Sign or Symptom|Medications|11036,11048|false|false|false|C0009806|Constipation|Constipation
Event|Event|Medications|11052,11058|false|false|false|||common
Finding|Functional Concept|Medications|11052,11058|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Finding|Intellectual Product|Medications|11052,11058|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Event|Event|Medications|11063,11067|false|false|false|||sure
Finding|Intellectual Product|Medications|11063,11067|false|false|false|C4724437|SURE Test|sure
Drug|Food|Medications|11071,11076|false|false|false|C0452428|Drink (dietary substance)|drink
Event|Event|Medications|11071,11076|false|false|false|||drink
Event|Event|Medications|11077,11083|false|false|false|||plenty
Drug|Substance|Medications|11087,11093|false|false|false|C0302908|Liquid substance|fluids
Event|Event|Medications|11087,11093|false|false|false|||fluids
Finding|Body Substance|Medications|11087,11093|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|Medications|11087,11093|false|false|false|C0016286|Fluid Therapy|fluids
Finding|Finding|Medications|11105,11109|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|Medications|11105,11109|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|Medications|11105,11109|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Procedure|Therapeutic or Preventive Procedure|Medications|11105,11120|false|false|false|C0301568|High residue diet|high-fiber diet
Anatomy|Tissue|Medications|11110,11115|false|false|false|C1304649|Tissue fiber|fiber
Drug|Organic Chemical|Medications|11110,11115|false|false|false|C0225326;C1321801|Fiber brand of calcium polycarbophil;fiber|fiber
Drug|Pharmacologic Substance|Medications|11110,11115|false|false|false|C0225326;C1321801|Fiber brand of calcium polycarbophil;fiber|fiber
Drug|Food|Medications|11116,11120|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|Medications|11116,11120|false|false|false|||diet
Finding|Functional Concept|Medications|11116,11120|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|Medications|11116,11120|false|false|false|C0012159|Diet therapy|diet
Drug|Hazardous or Poisonous Substance|Medications|11140,11149|false|false|false|C0027415|Narcotics|narcotics
Drug|Pharmacologic Substance|Medications|11140,11149|false|false|false|C0027415|Narcotics|narcotics
Event|Event|Medications|11140,11149|false|false|false|||narcotics
Attribute|Clinical Attribute|Medications|11151,11163|false|false|false|C5886759|Prescription (attribute)|prescription
Event|Event|Medications|11151,11163|false|false|false|||prescription
Finding|Intellectual Product|Medications|11151,11163|false|false|false|C1521941|prescription document|prescription
Procedure|Health Care Activity|Medications|11151,11163|false|false|false|C0033080|Prescription (procedure)|prescription
Attribute|Clinical Attribute|Medications|11165,11169|false|false|false|C2598155||pain
Finding|Functional Concept|Medications|11165,11169|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Medications|11165,11169|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|Medications|11170,11181|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Medications|11170,11181|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Medications|11170,11181|false|false|false|||medications
Finding|Intellectual Product|Medications|11170,11181|false|false|false|C4284232|Medications|medications
Event|Event|Medications|11184,11187|false|false|false|||try
Drug|Pharmacologic Substance|Medications|11191,11207|false|false|false|C0013231|Drugs, Non-Prescription|over-the-counter
Drug|Hazardous or Poisonous Substance|Medications|11200,11207|false|false|false|C0702263|Counter brand of Terbufos|counter
Drug|Organic Chemical|Medications|11200,11207|false|false|false|C0702263|Counter brand of Terbufos|counter
Event|Event|Medications|11208,11213|false|false|false|||stool
Finding|Body Substance|Medications|11208,11213|false|false|false|C0015733|Feces|stool
Drug|Organic Chemical|Medications|11208,11222|false|false|false|C0301470;C1154263|Stool Softener;Stool Softener brand of docusate sodium|stool softener
Drug|Pharmacologic Substance|Medications|11208,11222|false|false|false|C0301470;C1154263|Stool Softener;Stool Softener brand of docusate sodium|stool softener
Event|Event|Medications|11214,11222|false|false|false|||softener
Event|Event|Medications|11233,11237|false|false|false|||Call
Event|Event|Medications|11243,11249|false|false|false|||Doctor
Finding|Intellectual Product|Medications|11243,11249|false|false|false|C2348314|Doctor - Title|Doctor
Finding|Finding|Medications|11265,11271|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Finding|Intellectual Product|Medications|11265,11271|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Finding|Finding|Medications|11265,11276|false|false|false|C0278140;C4050465;C4521229|Neck Pain Score 6;Severe Extremity Pain;Severe pain|Severe pain
Attribute|Clinical Attribute|Medications|11272,11276|false|false|false|C2598155||pain
Event|Event|Medications|11272,11276|false|false|false|||pain
Finding|Functional Concept|Medications|11272,11276|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Medications|11272,11276|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Medications|11278,11286|false|false|false|||swelling
Finding|Finding|Medications|11278,11286|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|Medications|11278,11286|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Disorder|Disease or Syndrome|Medications|11288,11295|false|false|false|C0041834|Erythema|redness
Event|Event|Medications|11288,11295|false|false|false|||redness
Finding|Finding|Medications|11288,11295|false|false|false|C0332575|Redness|redness
Event|Event|Medications|11299,11307|false|false|false|||drainage
Finding|Body Substance|Medications|11299,11307|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|Medications|11299,11307|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|Medications|11299,11307|false|false|false|C0013103|Drainage procedure|drainage
Anatomy|Body Location or Region|Medications|11317,11325|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Medications|11317,11325|false|false|false|C0332803|Surgical wound|incision
Event|Event|Medications|11317,11325|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|Medications|11317,11325|false|false|false|C0184898|Surgical incisions|incision
Anatomy|Body Location or Region|Medications|11327,11331|false|false|false|C1515974|Anatomic Site|site
Finding|Intellectual Product|Medications|11327,11331|false|false|false|C1546778||site
Finding|Finding|Medications|11337,11342|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Finding|Sign or Symptom|Medications|11337,11342|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Finding|Intellectual Product|Medications|11362,11369|false|false|false|C0542560|Academic degree|degrees
Attribute|Clinical Attribute|Medications|11384,11390|false|false|false|C4255480||Nausea
Event|Event|Medications|11384,11390|false|false|false|||Nausea
Finding|Sign or Symptom|Medications|11384,11390|false|false|false|C0027497|Nausea|Nausea
Event|Event|Medications|11398,11406|true|false|false|||vomiting
Finding|Sign or Symptom|Medications|11398,11406|true|false|false|C0042963|Vomiting|vomiting
Finding|Finding|Medications|11410,11417|true|false|false|C4085555|Extreme Response|Extreme
Disorder|Mental or Behavioral Dysfunction|Medications|11418,11428|true|false|false|C2830004|Somnolence|sleepiness
Event|Event|Medications|11418,11428|true|false|false|||sleepiness
Finding|Finding|Medications|11418,11428|true|false|false|C0013144|Drowsiness|sleepiness
Event|Event|Medications|11443,11447|true|false|false|||able
Finding|Finding|Medications|11443,11447|true|true|false|C1299581|Able (qualifier value)|able
Event|Event|Medications|11451,11455|true|false|false|||stay
Drug|Organic Chemical|Medications|11451,11461|true|false|false|C0723446|Stay Awake|stay awake
Drug|Pharmacologic Substance|Medications|11451,11461|true|false|false|C0723446|Stay Awake|stay awake
Event|Event|Medications|11456,11461|true|false|false|||awake
Finding|Finding|Medications|11456,11461|true|false|false|C0234422|Awake (finding)|awake
Finding|Finding|Medications|11465,11471|true|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Finding|Intellectual Product|Medications|11465,11471|true|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Event|Event|Medications|11472,11481|true|false|false|||headaches
Finding|Sign or Symptom|Medications|11472,11481|true|false|false|C0018681|Headache|headaches
Event|Event|Medications|11486,11494|true|false|false|||relieved
Attribute|Clinical Attribute|Medications|11498,11502|true|true|false|C2598155||pain
Finding|Functional Concept|Medications|11498,11502|true|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Medications|11498,11502|true|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Hazardous or Poisonous Substance|Medications|11498,11512|true|false|false|C0002771;C0722425|Analgesics;Pain Relieve brand of acetaminophen|pain relievers
Drug|Organic Chemical|Medications|11498,11512|true|false|false|C0002771;C0722425|Analgesics;Pain Relieve brand of acetaminophen|pain relievers
Drug|Pharmacologic Substance|Medications|11498,11512|true|false|false|C0002771;C0722425|Analgesics;Pain Relieve brand of acetaminophen|pain relievers
Event|Event|Medications|11503,11512|true|false|false|||relievers
Event|Event|Medications|11516,11524|true|false|false|||Seizures
Finding|Sign or Symptom|Medications|11516,11524|true|false|false|C0036572|Seizures|Seizures
Finding|Finding|Medications|11532,11535|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Medications|11532,11535|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Event|Event|Medications|11536,11544|true|false|false|||problems
Finding|Idea or Concept|Medications|11536,11544|true|false|false|C1546466|Problems - What subject filter|problems
Attribute|Clinical Attribute|Medications|11555,11561|true|false|false|C2707266||vision
Event|Event|Medications|11555,11561|true|false|false|||vision
Finding|Organism Function|Medications|11555,11561|true|false|false|C0042789|Vision|vision
Event|Event|Medications|11565,11572|true|false|false|||ability
Finding|Functional Concept|Medications|11565,11572|true|false|false|C5891046|Oral Intake Ability|ability
Finding|Intellectual Product|Medications|11565,11575|true|false|false|C5420000|Ability Question|ability to
Finding|Finding|Medications|11565,11581|true|false|false|C0564214|Ability to speak|ability to speak
Event|Event|Medications|11576,11581|false|false|false|||speak
Finding|Finding|Medications|11576,11581|false|false|false|C0234856;C0600116;C1547187|Does speak;Speak - language ability;Speaking (function)|speak
Finding|Idea or Concept|Medications|11576,11581|false|false|false|C0234856;C0600116;C1547187|Does speak;Speak - language ability;Speaking (function)|speak
Finding|Individual Behavior|Medications|11576,11581|false|false|false|C0234856;C0600116;C1547187|Does speak;Speak - language ability;Speaking (function)|speak
Event|Event|Medications|11585,11593|false|false|false|||Weakness
Finding|Sign or Symptom|Medications|11585,11593|false|false|false|C0004093;C3714552|Asthenia;Weakness|Weakness
Event|Event|Medications|11597,11604|false|false|false|||changes
Finding|Functional Concept|Medications|11597,11604|false|false|false|C0392747|Changing|changes
Event|Event|Medications|11608,11617|false|false|false|||sensation
Finding|Finding|Medications|11608,11617|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|Medications|11608,11617|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|Medications|11608,11617|false|false|false|C2229507|sensory exam|sensation
Anatomy|Body Location or Region|Medications|11626,11630|false|false|false|C0015450;C4266571|Face;Head>Face|face
Disorder|Disease or Syndrome|Medications|11626,11630|false|false|false|C3160739|FANCONI ANEMIA, COMPLEMENTATION GROUP E|face
Finding|Gene or Genome|Medications|11626,11630|false|false|false|C1414531;C1423759;C2828055|ELOVL6 gene;FANCE gene;FANCE wt Allele|face
Anatomy|Body Part, Organ, or Organ Component|Medications|11632,11636|false|false|false|C0446516|Upper arm|arms
Attribute|Clinical Attribute|Medications|11632,11636|false|false|false|C5782111||arms
Disorder|Neoplastic Process|Medications|11632,11636|false|false|false|C0206655|Alveolar rhabdomyosarcoma|arms
Event|Event|Medications|11632,11636|false|false|false|||arms
Finding|Gene or Genome|Medications|11632,11636|false|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Finding|Intellectual Product|Medications|11632,11636|false|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Anatomy|Body Part, Organ, or Organ Component|Medications|11641,11644|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Functional Concept|Medications|11646,11650|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|Call
Finding|Gene or Genome|Medications|11646,11650|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|Call
Finding|Intellectual Product|Medications|11646,11650|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|Call
Finding|Mental Process|Medications|11646,11650|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|Call
Finding|Finding|Medications|11677,11686|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Idea or Concept|Medications|11677,11686|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Intellectual Product|Medications|11677,11686|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Pathologic Function|Medications|11677,11686|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Phenomenon|Phenomenon or Process|Medications|11677,11686|false|false|false|C0013956|Emergency Situation|Emergency
Procedure|Health Care Activity|Medications|11677,11686|false|false|false|C1553500|emergency encounter|Emergency
Finding|Idea or Concept|Medications|11677,11691|false|false|false|C1546435|Encounter Referral Source - emergency room|Emergency Room
Finding|Mental Process|Medications|11699,11709|true|false|false|C0237607;C0596545|Experience;Experience (Practice)|experience
Event|Event|Medications|11743,11751|false|false|false|||numbness
Finding|Finding|Medications|11743,11751|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|Medications|11743,11751|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Event|Event|Medications|11755,11763|false|false|false|||weakness
Finding|Sign or Symptom|Medications|11755,11763|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Anatomy|Body Location or Region|Medications|11771,11775|false|false|false|C0015450;C4266571|Face;Head>Face|face
Disorder|Disease or Syndrome|Medications|11771,11775|false|false|false|C3160739|FANCONI ANEMIA, COMPLEMENTATION GROUP E|face
Finding|Gene or Genome|Medications|11771,11775|false|false|false|C1414531;C1423759;C2828055|ELOVL6 gene;FANCE gene;FANCE wt Allele|face
Anatomy|Body Part, Organ, or Organ Component|Medications|11777,11780|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|Medications|11777,11780|false|false|false|C3495676|Anorectal Malformations|arm
Event|Event|Medications|11777,11780|false|false|false|||arm
Finding|Gene or Genome|Medications|11777,11780|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|Medications|11777,11780|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|Medications|11777,11780|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|Medications|11777,11780|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Anatomy|Body Part, Organ, or Organ Component|Medications|11785,11788|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Disorder|Mental or Behavioral Dysfunction|Medications|11799,11808|false|false|false|C0009676|Confusion|confusion
Event|Event|Medications|11799,11808|false|false|false|||confusion
Finding|Finding|Medications|11799,11808|false|false|false|C0683369|Clouded consciousness|confusion
Event|Event|Medications|11812,11819|false|false|false|||trouble
Event|Event|Medications|11820,11828|false|false|false|||speaking
Event|Event|Medications|11832,11845|false|false|false|||understanding
Finding|Mental Process|Medications|11832,11845|false|false|false|C0162340|Comprehension|understanding
Event|Event|Medications|11864,11871|false|false|false|||walking
Event|Event|Medications|11873,11882|false|false|false|||dizziness
Finding|Sign or Symptom|Medications|11873,11882|false|false|false|C0012833;C0042571|Dizziness;Vertigo|dizziness
Event|Event|Medications|11887,11891|false|false|false|||loss
Finding|Finding|Medications|11887,11891|false|false|false|C5890125|Loss (adaptation)|loss
Finding|Finding|Medications|11887,11902|false|false|false|C0241981|Impairment of balance|loss of balance
Drug|Organic Chemical|Medications|11895,11902|false|false|false|C4319618|Balance (substance)|balance
Drug|Pharmacologic Substance|Medications|11895,11902|false|false|false|C4319618|Balance (substance)|balance
Event|Event|Medications|11895,11902|false|false|false|||balance
Finding|Finding|Medications|11895,11902|false|false|false|C0014653;C0560184|Ability to balance;Equilibrium|balance
Finding|Organism Function|Medications|11895,11902|false|false|false|C0014653;C0560184|Ability to balance;Equilibrium|balance
Procedure|Diagnostic Procedure|Medications|11895,11902|false|false|false|C2174421|examination of balance|balance
Event|Event|Medications|11907,11919|false|false|false|||coordination
Finding|Functional Concept|Medications|11907,11919|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|coordination
Finding|Idea or Concept|Medications|11907,11919|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|coordination
Finding|Physiologic Function|Medications|11907,11919|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|coordination
Finding|Finding|Medications|11930,11936|true|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Medications|11930,11936|true|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Event|Event|Medications|11937,11946|true|false|false|||headaches
Finding|Sign or Symptom|Medications|11937,11946|true|false|false|C0018681|Headache|headaches
Event|Event|Medications|11961,11967|true|false|false|||reason
Finding|Idea or Concept|Medications|11961,11967|true|false|false|C0392360|Indication of (contextual qualifier)|reason
Procedure|Health Care Activity|Medications|11971,11979|true|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Medications|11980,11992|true|false|false|C3263700||Instructions
Event|Event|Medications|11980,11992|true|false|false|||Instructions
Finding|Intellectual Product|Medications|11980,11992|true|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

