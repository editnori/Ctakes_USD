 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|25,29
No|30,32
:|32,33
_|36,37
_|37,38
_|38,39
<EOL>|39,40
<EOL>|41,42
Admission|42,51
Date|52,56
:|56,57
_|59,60
_|60,61
_|61,62
Discharge|76,85
Date|86,90
:|90,91
_|94,95
_|95,96
_|96,97
<EOL>|97,98
<EOL>|99,100
Date|100,104
of|105,107
Birth|108,113
:|113,114
_|116,117
_|117,118
_|118,119
Sex|132,135
:|135,136
F|139,140
<EOL>|140,141
<EOL>|142,143
Service|143,150
:|150,151
MEDICINE|152,160
<EOL>|160,161
<EOL>|162,163
IV|175,177
Dye|178,181
,|181,182
Iodine|183,189
Containing|190,200
Contrast|201,209
Media|210,215
/|216,217
Oxycodone|218,227
/|228,229
<EOL>|230,231
cilostazol|231,241
/|242,243
Varenicline|244,255
<EOL>|255,256
<EOL>|257,258
Attending|258,267
:|267,268
_|269,270
_|270,271
_|271,272
.|272,273
<EOL>|273,274
<EOL>|275,276
cough|293,298
,|298,299
dyspnea|300,307
<EOL>|307,308
<EOL>|309,310
Major|310,315
Surgical|316,324
or|325,327
Invasive|328,336
Procedure|337,346
:|346,347
<EOL>|347,348
None|348,352
<EOL>|352,353
<EOL>|353,354
<EOL>|355,356
HPI|384,387
:|387,388
_|389,390
_|390,391
_|391,392
year|393,397
old|398,401
female|402,408
with|409,413
history|414,421
of|422,424
COPD|425,429
(|430,431
on|431,433
home|434,438
O2|439,441
)|441,442
,|442,443
HTN|444,447
,|447,448
<EOL>|449,450
Afib|450,454
admitted|455,463
with|464,468
dyspnea|469,476
and|477,480
cough|481,486
.|486,487
<EOL>|489,490
Pt|491,493
states|494,500
inc|501,504
dyspnea|505,512
since|513,518
this|519,523
am|524,526
,|526,527
also|528,532
one|533,536
episode|537,544
of|545,547
<EOL>|548,549
retrosternal|549,561
chest|562,567
pressure|568,576
lasting|577,584
2minuts|585,592
on|593,595
way|596,599
to|600,602
ED|603,605
.|605,606
No|607,609
cp|610,612
<EOL>|613,614
currently|614,623
.|623,624
on|625,627
home|628,632
O2|633,635
.|635,636
no|637,639
fevers|640,646
/|646,647
chills|647,653
or|654,656
abd|657,660
sx|661,663
.|663,664
<EOL>|666,667
Patient|668,675
was|676,679
recently|680,688
admitted|689,697
from|698,702
_|703,704
_|704,705
_|705,706
with|707,711
COPD|712,716
flare|717,722
<EOL>|723,724
and|724,727
afib|728,732
with|733,737
RVR|738,741
.|741,742
She|743,746
could|747,752
not|753,756
receive|757,764
azithromycin|765,777
due|778,781
to|782,784
<EOL>|785,786
concern|786,793
for|794,797
QTc|798,801
prolongation|802,814
and|815,818
so|819,821
was|822,825
treated|826,833
with|834,838
<EOL>|839,840
ceftriaxone|840,851
/|851,852
cefpodoxime|852,863
.|863,864
She|865,868
was|869,872
treated|873,880
with|881,885
60mg|886,890
PO|891,893
prednisone|894,904
<EOL>|905,906
and|906,909
discharged|910,920
with|921,925
a|926,927
prednisone|928,938
taper|939,944
of|945,947
10|948,950
mg|951,953
decrease|954,962
q3d|963,966
<EOL>|967,968
until|968,973
at|974,976
10|977,979
mg|980,982
,|982,983
then|984,988
stay|989,993
at|994,996
10|997,999
mg|1000,1002
until|1003,1008
pulm|1009,1013
follow|1014,1020
up|1021,1023
.|1023,1024
She|1025,1028
was|1029,1032
<EOL>|1033,1034
also|1034,1038
counseled|1039,1048
to|1049,1051
do|1052,1054
pulmonary|1055,1064
rehab|1065,1070
and|1071,1074
follow|1075,1081
up|1082,1084
with|1085,1089
Dr|1090,1092
.|1092,1093
<EOL>|1094,1095
_|1095,1096
_|1096,1097
_|1097,1098
.|1098,1099
She|1100,1103
was|1104,1107
discharged|1108,1118
on|1119,1121
2L|1122,1124
supplemental|1125,1137
O2|1138,1140
to|1141,1143
be|1144,1146
worn|1147,1151
at|1152,1154
<EOL>|1155,1156
all|1156,1159
times|1160,1165
.|1165,1166
He|1167,1169
theophylline|1170,1182
was|1183,1186
decreased|1187,1196
from|1197,1201
300|1202,1205
mg|1206,1208
BID|1209,1212
to|1213,1215
_|1216,1217
_|1217,1218
_|1218,1219
<EOL>|1220,1221
mg|1221,1223
BID|1224,1227
due|1228,1231
to|1232,1234
her|1235,1238
afib|1239,1243
with|1244,1248
RVR|1249,1252
.|1252,1253
<EOL>|1255,1256
She|1257,1260
was|1261,1264
also|1265,1269
seen|1270,1274
in|1275,1277
the|1278,1281
ED|1282,1284
on|1285,1287
_|1288,1289
_|1289,1290
_|1290,1291
and|1292,1295
_|1296,1297
_|1297,1298
_|1298,1299
due|1300,1303
to|1304,1306
dyspnea|1307,1314
<EOL>|1315,1316
which|1316,1321
was|1322,1325
felt|1326,1330
to|1331,1333
be|1334,1336
a|1337,1338
continuation|1339,1351
of|1352,1354
her|1355,1358
COPD|1359,1363
flare|1364,1369
in|1370,1372
the|1373,1376
<EOL>|1377,1378
setting|1378,1385
of|1386,1388
patient|1389,1396
not|1397,1400
taking|1401,1407
her|1408,1411
home|1412,1416
medications|1417,1428
.|1428,1429
She|1430,1433
was|1434,1437
<EOL>|1438,1439
given|1439,1444
nebulizers|1445,1455
and|1456,1459
improved|1460,1468
.|1468,1469
She|1470,1473
was|1474,1477
DCed|1478,1482
home|1483,1487
with|1488,1492
_|1493,1494
_|1494,1495
_|1495,1496
for|1497,1500
<EOL>|1501,1502
assistance|1502,1512
with|1513,1517
medications|1518,1529
.|1529,1530
She|1531,1534
declined|1535,1543
pulmonary|1544,1553
rehab|1554,1559
<EOL>|1560,1561
facility|1561,1569
disposition|1570,1581
.|1581,1582
<EOL>|1584,1585
<EOL>|1585,1586
In|1586,1588
the|1589,1592
ED|1593,1595
,|1595,1596
initial|1597,1604
vitals|1605,1611
:|1611,1612
<EOL>|1614,1615
-|1615,1616
Exam|1617,1621
notable|1622,1629
for|1630,1633
:|1633,1634
diffuse|1635,1642
insp|1643,1647
/|1647,1648
esp|1648,1651
wheezing|1652,1660
,|1660,1661
dry|1662,1665
oropharynx|1666,1676
<EOL>|1678,1679
-|1679,1680
Labs|1681,1685
notable|1686,1693
for|1694,1697
:|1697,1698
nl|1699,1701
WBC|1702,1705
.|1705,1706
Trop|1707,1711
X1|1712,1714
neg|1715,1718
.|1718,1719
EKG|1720,1723
in|1724,1726
sinus|1727,1732
.|1732,1733
<EOL>|1733,1734
-|1734,1735
Imaging|1736,1743
notable|1744,1751
for|1752,1755
:|1755,1756
CXR|1757,1760
no|1761,1763
acute|1764,1769
process|1770,1777
.|1777,1778
<EOL>|1779,1780
-|1780,1781
Pt|1782,1784
given|1785,1790
:|1790,1791
duoneb|1792,1798
X|1799,1800
3.|1801,1803
methylpred|1804,1814
125mg|1815,1820
.|1820,1821
Aspirin|1822,1829
325mg|1830,1835
,|1835,1836
1L|1837,1839
NS|1840,1842
,|1842,1843
<EOL>|1844,1845
and|1845,1848
azithromycin|1849,1861
500mg|1862,1867
.|1867,1868
Peak|1869,1873
flow|1874,1878
150|1879,1882
,|1882,1883
baseline|1884,1892
per|1893,1896
pt|1897,1899
.|1899,1900
Symptoms|1901,1909
<EOL>|1910,1911
overall|1911,1918
improved|1919,1927
after|1928,1933
nebs|1934,1938
.|1938,1939
<EOL>|1940,1941
-|1941,1942
Vitals|1943,1949
prior|1950,1955
to|1956,1958
transfer|1959,1967
:|1967,1968
98.2|1969,1973
76|1974,1976
138|1977,1980
/|1980,1981
72|1981,1983
20|1984,1986
97NC|1987,1991
.|1991,1992
<EOL>|1994,1995
<EOL>|1995,1996
On|1996,1998
arrival|1999,2006
to|2007,2009
the|2010,2013
floor|2014,2019
,|2019,2020
pt|2021,2023
reports|2024,2031
feeling|2032,2039
much|2040,2044
improved|2045,2053
and|2054,2057
<EOL>|2058,2059
minimal|2059,2066
wheezing|2067,2075
.|2075,2076
<EOL>|2076,2077
<EOL>|2077,2078
No|2085,2087
fevers|2088,2094
,|2094,2095
chills|2096,2102
,|2102,2103
night|2104,2109
sweats|2110,2116
,|2116,2117
or|2118,2120
weight|2121,2127
changes|2128,2135
.|2135,2136
No|2137,2139
changes|2140,2147
<EOL>|2148,2149
in|2149,2151
vision|2152,2158
or|2159,2161
hearing|2162,2169
,|2169,2170
no|2171,2173
changes|2174,2181
in|2182,2184
balance|2185,2192
.|2192,2193
No|2194,2196
cough|2197,2202
,|2202,2203
no|2204,2206
<EOL>|2207,2208
shortness|2208,2217
of|2218,2220
breath|2221,2227
,|2227,2228
no|2229,2231
dyspnea|2232,2239
on|2240,2242
exertion|2243,2251
.|2251,2252
No|2253,2255
chest|2256,2261
pain|2262,2266
or|2267,2269
<EOL>|2270,2271
palpitations|2271,2283
.|2283,2284
No|2285,2287
nausea|2288,2294
or|2295,2297
vomiting|2298,2306
.|2306,2307
No|2308,2310
diarrhea|2311,2319
or|2320,2322
<EOL>|2323,2324
constipation|2324,2336
.|2336,2337
No|2338,2340
dysuria|2341,2348
or|2349,2351
hematuria|2352,2361
.|2361,2362
No|2363,2365
hematochezia|2366,2378
,|2378,2379
no|2380,2382
<EOL>|2383,2384
melena|2384,2390
.|2390,2391
No|2392,2394
numbness|2395,2403
or|2404,2406
weakness|2407,2415
,|2415,2416
no|2417,2419
focal|2420,2425
deficits|2426,2434
.|2434,2435
<EOL>|2437,2438
<EOL>|2438,2439
<EOL>|2440,2441
ASTHMA|2463,2469
/|2469,2470
COPD|2470,2474
<EOL>|2476,2477
ATYPICAL|2478,2486
CHEST|2487,2492
PAIN|2493,2497
<EOL>|2499,2500
CERVICAL|2501,2509
RADICULITIS|2510,2521
<EOL>|2523,2524
CERVICAL|2525,2533
SPONDYLOSIS|2534,2545
<EOL>|2547,2548
CORONARY|2549,2557
ARTERY|2558,2564
DISEASE|2565,2572
<EOL>|2574,2575
HEADACHE|2576,2584
<EOL>|2586,2587
HIP|2588,2591
REPLACEMENT|2592,2603
<EOL>|2605,2606
HYPERLIPIDEMIA|2607,2621
<EOL>|2623,2624
HYPERTENSION|2625,2637
<EOL>|2639,2640
OSTEOARTHRITIS|2641,2655
<EOL>|2657,2658
HERPES|2659,2665
ZOSTER|2666,2672
<EOL>|2674,2675
ATRIAL|2676,2682
FIBRILLATION|2683,2695
<EOL>|2697,2698
ANXIETY|2699,2706
<EOL>|2708,2709
GASTROINTESTINAL|2710,2726
BLEEDING|2727,2735
<EOL>|2737,2738
OSTEOARTHRITIS|2739,2753
<EOL>|2755,2756
ATHEROSCLEROTIC|2757,2772
CARDIOVASCULAR|2773,2787
DISEASE|2788,2795
<EOL>|2797,2798
PERIPHERAL|2799,2809
VASCULAR|2810,2818
DISEASE|2819,2826
<EOL>|2826,2827
<EOL>|2828,2829
:|2843,2844
<EOL>|2844,2845
_|2845,2846
_|2846,2847
_|2847,2848
<EOL>|2848,2849
:|2863,2864
<EOL>|2864,2865
Mother|2865,2871
:|2871,2872
_|2873,2874
_|2874,2875
_|2875,2876
,|2876,2877
HTN|2878,2881
<EOL>|2883,2884
Father|2884,2890
:|2890,2891
_|2892,2893
_|2893,2894
_|2894,2895
CA|2896,2898
<EOL>|2900,2901
Brother|2901,2908
:|2908,2909
CA|2910,2912
?|2912,2913
<EOL>|2915,2916
Brother|2916,2923
:|2923,2924
_|2925,2926
_|2926,2927
_|2927,2928
<EOL>|2929,2930
<EOL>|2931,2932
Physical|2932,2940
_|2941,2942
_|2942,2943
_|2943,2944
:|2944,2945
<EOL>|2945,2946
Admission|2946,2955
<EOL>|2955,2956
<EOL>|2956,2957
Vitals|2957,2963
:|2963,2964
99|2965,2967
142|2968,2971
/|2971,2972
80|2972,2974
77|2975,2977
20|2978,2980
95|2981,2983
/|2983,2984
2L|2984,2986
<EOL>|2987,2988
General|2988,2995
:|2995,2996
Alert|2997,3002
,|3002,3003
oriented|3004,3012
,|3012,3013
no|3014,3016
acute|3017,3022
distress|3023,3031
,|3031,3032
appears|3033,3040
very|3041,3045
calm|3046,3050
<EOL>|3051,3052
and|3052,3055
can|3056,3059
talk|3060,3064
in|3065,3067
full|3068,3072
sentences|3073,3082
<EOL>|3083,3084
HEENT|3084,3089
:|3089,3090
Sclerae|3091,3098
anicteric|3099,3108
,|3108,3109
MMM|3110,3113
,|3113,3114
oropharynx|3115,3125
clear|3126,3131
<EOL>|3133,3134
Neck|3134,3138
:|3138,3139
supple|3140,3146
,|3146,3147
JVP|3148,3151
not|3152,3155
elevated|3156,3164
,|3164,3165
no|3166,3168
LAD|3169,3172
<EOL>|3174,3175
Lungs|3175,3180
:|3180,3181
scattered|3182,3191
wheezing|3192,3200
<EOL>|3202,3203
CV|3203,3205
:|3205,3206
II|3207,3209
/|3209,3210
VI|3210,3212
RUSB|3213,3217
systolic|3218,3226
murmur|3227,3233
,|3233,3234
Nl|3235,3237
S1|3238,3240
,|3240,3241
S2|3242,3244
,|3244,3245
No|3246,3248
MRG|3249,3252
<EOL>|3254,3255
Abdomen|3255,3262
:|3262,3263
soft|3264,3268
,|3268,3269
NT|3270,3272
/|3272,3273
ND|3273,3275
bowel|3276,3281
sounds|3282,3288
present|3289,3296
,|3296,3297
no|3298,3300
rebound|3301,3308
tenderness|3309,3319
<EOL>|3320,3321
or|3321,3323
guarding|3324,3332
,|3332,3333
no|3334,3336
organomegaly|3337,3349
<EOL>|3351,3352
GU|3352,3354
:|3354,3355
no|3356,3358
foley|3359,3364
<EOL>|3366,3367
Ext|3367,3370
:|3370,3371
warm|3372,3376
,|3376,3377
well|3378,3382
perfused|3383,3391
,|3391,3392
2|3393,3394
+|3394,3395
pulses|3396,3402
,|3402,3403
no|3404,3406
clubbing|3407,3415
,|3415,3416
cyanosis|3417,3425
,|3425,3426
2|3427,3428
+|3428,3429
<EOL>|3430,3431
edema|3431,3436
b|3437,3438
/|3438,3439
l|3439,3440
<EOL>|3440,3441
Neuro|3441,3446
:|3446,3447
CN2|3448,3451
-|3451,3452
12|3452,3454
intact|3455,3461
,|3461,3462
no|3463,3465
focal|3466,3471
deficits|3472,3480
<EOL>|3481,3482
<EOL>|3482,3483
Vitals|3483,3489
:|3489,3490
98.5|3491,3495
122|3496,3499
/|3499,3500
69|3500,3502
(|3502,3503
130|3503,3506
-|3506,3507
150|3507,3510
)|3510,3511
76|3512,3514
(|3514,3515
70s|3515,3518
)|3518,3519
18|3520,3522
100|3523,3526
/|3526,3527
2L|3527,3529
<EOL>|3530,3531
General|3531,3538
:|3538,3539
Alert|3540,3545
,|3545,3546
oriented|3547,3555
,|3555,3556
no|3557,3559
acute|3560,3565
distress|3566,3574
,|3574,3575
appears|3576,3583
very|3584,3588
calm|3589,3593
<EOL>|3594,3595
and|3595,3598
can|3599,3602
talk|3603,3607
in|3608,3610
full|3611,3615
sentences|3616,3625
<EOL>|3626,3627
HEENT|3627,3632
:|3632,3633
Sclerae|3634,3641
anicteric|3642,3651
,|3651,3652
MMM|3653,3656
,|3656,3657
oropharynx|3658,3668
clear|3669,3674
<EOL>|3676,3677
Neck|3677,3681
:|3681,3682
supple|3683,3689
,|3689,3690
JVP|3691,3694
not|3695,3698
elevated|3699,3707
,|3707,3708
no|3709,3711
LAD|3712,3715
<EOL>|3717,3718
Lungs|3718,3723
:|3723,3724
scattered|3725,3734
wheezing|3735,3743
<EOL>|3745,3746
CV|3746,3748
:|3748,3749
II|3750,3752
/|3752,3753
VI|3753,3755
RUSB|3756,3760
systolic|3761,3769
murmur|3770,3776
,|3776,3777
Nl|3778,3780
S1|3781,3783
,|3783,3784
S2|3785,3787
,|3787,3788
No|3789,3791
MRG|3792,3795
<EOL>|3797,3798
Abdomen|3798,3805
:|3805,3806
soft|3807,3811
,|3811,3812
NT|3813,3815
/|3815,3816
ND|3816,3818
bowel|3819,3824
sounds|3825,3831
present|3832,3839
,|3839,3840
no|3841,3843
rebound|3844,3851
tenderness|3852,3862
<EOL>|3863,3864
or|3864,3866
guarding|3867,3875
,|3875,3876
no|3877,3879
organomegaly|3880,3892
<EOL>|3894,3895
GU|3895,3897
:|3897,3898
no|3899,3901
foley|3902,3907
<EOL>|3909,3910
Ext|3910,3913
:|3913,3914
warm|3915,3919
,|3919,3920
well|3921,3925
perfused|3926,3934
,|3934,3935
2|3936,3937
+|3937,3938
pulses|3939,3945
,|3945,3946
no|3947,3949
clubbing|3950,3958
,|3958,3959
cyanosis|3960,3968
,|3968,3969
2|3970,3971
+|3971,3972
<EOL>|3973,3974
edema|3974,3979
b|3980,3981
/|3981,3982
l|3982,3983
<EOL>|3983,3984
Neuro|3984,3989
:|3989,3990
CN2|3991,3994
-|3994,3995
12|3995,3997
intact|3998,4004
,|4004,4005
no|4006,4008
focal|4009,4014
deficits|4015,4023
<EOL>|4023,4024
<EOL>|4025,4026
Pertinent|4026,4035
Results|4036,4043
:|4043,4044
<EOL>|4044,4045
Admission|4045,4054
<EOL>|4054,4055
<EOL>|4055,4056
_|4056,4057
_|4057,4058
_|4058,4059
01|4060,4062
:|4062,4063
46PM|4063,4067
BLOOD|4068,4073
WBC|4074,4077
-|4077,4078
8.3|4078,4081
RBC|4082,4085
-|4085,4086
4|4086,4087
.|4087,4088
52|4088,4090
Hgb|4091,4094
-|4094,4095
10|4095,4097
.|4097,4098
8|4098,4099
*|4099,4100
Hct|4101,4104
-|4104,4105
36.2|4105,4109
<EOL>|4110,4111
MCV|4111,4114
-|4114,4115
80|4115,4117
*|4117,4118
MCH|4119,4122
-|4122,4123
23|4123,4125
.|4125,4126
9|4126,4127
*|4127,4128
MCHC|4129,4133
-|4133,4134
29|4134,4136
.|4136,4137
8|4137,4138
*|4138,4139
RDW|4140,4143
-|4143,4144
21|4144,4146
.|4146,4147
6|4147,4148
*|4148,4149
RDWSD|4150,4155
-|4155,4156
52|4156,4158
.|4158,4159
4|4159,4160
*|4160,4161
Plt|4162,4165
_|4166,4167
_|4167,4168
_|4168,4169
<EOL>|4169,4170
_|4170,4171
_|4171,4172
_|4172,4173
01|4174,4176
:|4176,4177
46PM|4177,4181
BLOOD|4182,4187
Neuts|4188,4193
-|4193,4194
93|4194,4196
.|4196,4197
4|4197,4198
*|4198,4199
Lymphs|4200,4206
-|4206,4207
4|4207,4208
.|4208,4209
0|4209,4210
*|4210,4211
Monos|4212,4217
-|4217,4218
1|4218,4219
.|4219,4220
8|4220,4221
*|4221,4222
<EOL>|4223,4224
Eos|4224,4227
-|4227,4228
0|4228,4229
.|4229,4230
1|4230,4231
*|4231,4232
Baso|4233,4237
-|4237,4238
0.1|4238,4241
Im|4242,4244
_|4245,4246
_|4246,4247
_|4247,4248
AbsNeut|4249,4256
-|4256,4257
7|4257,4258
.|4258,4259
77|4259,4261
*|4261,4262
AbsLymp|4263,4270
-|4270,4271
0|4271,4272
.|4272,4273
33|4273,4275
*|4275,4276
<EOL>|4277,4278
AbsMono|4278,4285
-|4285,4286
0|4286,4287
.|4287,4288
15|4288,4290
*|4290,4291
AbsEos|4292,4298
-|4298,4299
0|4299,4300
.|4300,4301
01|4301,4303
*|4303,4304
AbsBaso|4305,4312
-|4312,4313
0.01|4313,4317
<EOL>|4317,4318
_|4318,4319
_|4319,4320
_|4320,4321
01|4322,4324
:|4324,4325
46PM|4325,4329
BLOOD|4330,4335
_|4336,4337
_|4337,4338
_|4338,4339
PTT|4340,4343
-|4343,4344
31.9|4344,4348
_|4349,4350
_|4350,4351
_|4351,4352
<EOL>|4352,4353
_|4353,4354
_|4354,4355
_|4355,4356
01|4357,4359
:|4359,4360
46PM|4360,4364
BLOOD|4365,4370
Glucose|4371,4378
-|4378,4379
121|4379,4382
*|4382,4383
UreaN|4384,4389
-|4389,4390
19|4390,4392
Creat|4393,4398
-|4398,4399
1.1|4399,4402
Na|4403,4405
-|4405,4406
134|4406,4409
<EOL>|4410,4411
K|4411,4412
-|4412,4413
3.7|4413,4416
Cl|4417,4419
-|4419,4420
91|4420,4422
*|4422,4423
HCO3|4424,4428
-|4428,4429
31|4429,4431
AnGap|4432,4437
-|4437,4438
16|4438,4440
<EOL>|4440,4441
_|4441,4442
_|4442,4443
_|4443,4444
01|4445,4447
:|4447,4448
46PM|4448,4452
BLOOD|4453,4458
cTropnT|4459,4466
-|4466,4467
<|4467,4468
0|4468,4469
.|4469,4470
01|4470,4472
<EOL>|4472,4473
_|4473,4474
_|4474,4475
_|4475,4476
01|4477,4479
:|4479,4480
46PM|4480,4484
BLOOD|4485,4490
Calcium|4491,4498
-|4498,4499
10.1|4499,4503
Phos|4504,4508
-|4508,4509
2.7|4509,4512
Mg|4513,4515
-|4515,4516
2.1|4516,4519
<EOL>|4519,4520
_|4520,4521
_|4521,4522
_|4522,4523
01|4524,4526
:|4526,4527
58PM|4527,4531
BLOOD|4532,4537
Lactate|4538,4545
-|4545,4546
1.6|4546,4549
<EOL>|4549,4550
<EOL>|4550,4551
DISCHARGE|4551,4560
<EOL>|4560,4561
<EOL>|4561,4562
_|4562,4563
_|4563,4564
_|4564,4565
05|4566,4568
:|4568,4569
52AM|4569,4573
BLOOD|4574,4579
WBC|4580,4583
-|4583,4584
14|4584,4586
.|4586,4587
1|4587,4588
*|4588,4589
#|4589,4590
RBC|4591,4594
-|4594,4595
3|4595,4596
.|4596,4597
81|4597,4599
*|4599,4600
Hgb|4601,4604
-|4604,4605
9|4605,4606
.|4606,4607
4|4607,4608
*|4608,4609
Hct|4610,4613
-|4613,4614
30|4614,4616
.|4616,4617
8|4617,4618
*|4618,4619
<EOL>|4620,4621
MCV|4621,4624
-|4624,4625
81|4625,4627
*|4627,4628
MCH|4629,4632
-|4632,4633
24|4633,4635
.|4635,4636
7|4636,4637
*|4637,4638
MCHC|4639,4643
-|4643,4644
30|4644,4646
.|4646,4647
5|4647,4648
*|4648,4649
RDW|4650,4653
-|4653,4654
22|4654,4656
.|4656,4657
5|4657,4658
*|4658,4659
RDWSD|4660,4665
-|4665,4666
58|4666,4668
.|4668,4669
1|4669,4670
*|4670,4671
Plt|4672,4675
_|4676,4677
_|4677,4678
_|4678,4679
<EOL>|4679,4680
_|4680,4681
_|4681,4682
_|4682,4683
05|4684,4686
:|4686,4687
52AM|4687,4691
BLOOD|4692,4697
Glucose|4698,4705
-|4705,4706
107|4706,4709
*|4709,4710
UreaN|4711,4716
-|4716,4717
26|4717,4719
*|4719,4720
Creat|4721,4726
-|4726,4727
0.9|4727,4730
Na|4731,4733
-|4733,4734
136|4734,4737
<EOL>|4738,4739
K|4739,4740
-|4740,4741
3.5|4741,4744
Cl|4745,4747
-|4747,4748
94|4748,4750
*|4750,4751
HCO3|4752,4756
-|4756,4757
35|4757,4759
*|4759,4760
AnGap|4761,4766
-|4766,4767
11|4767,4769
<EOL>|4769,4770
<EOL>|4770,4771
CXR|4771,4774
_|4775,4776
_|4776,4777
_|4777,4778
<EOL>|4778,4779
<EOL>|4779,4780
No|4797,4799
acute|4800,4805
cardiopulmonary|4806,4821
process|4822,4829
.|4829,4830
<EOL>|4831,4832
<EOL>|4832,4833
<EOL>|4834,4835
_|4858,4859
_|4859,4860
_|4860,4861
year|4862,4866
old|4867,4870
female|4871,4877
with|4878,4882
history|4883,4890
of|4891,4893
COPD|4894,4898
(|4899,4900
on|4900,4902
home|4903,4907
O2|4908,4910
)|4910,4911
,|4911,4912
HTN|4913,4916
,|4916,4917
Afib|4918,4922
<EOL>|4923,4924
admitted|4924,4932
with|4933,4937
dyspnea|4938,4945
and|4946,4949
cough|4950,4955
.|4955,4956
<EOL>|4958,4959
<EOL>|4959,4960
#|4960,4961
COPD|4963,4967
exacerbation|4968,4980
:|4980,4981
Presenting|4982,4992
with|4993,4997
cough|4998,5003
,|5003,5004
significant|5005,5016
<EOL>|5017,5018
wheezing|5018,5026
and|5027,5030
poor|5031,5035
air|5036,5039
movement|5040,5048
initially|5049,5058
consistent|5059,5069
with|5070,5074
COPD|5075,5079
<EOL>|5080,5081
exacerbation|5081,5093
.|5093,5094
No|5095,5097
PNA|5098,5101
on|5102,5104
CXR|5105,5108
.|5108,5109
No|5110,5112
ischemic|5113,5121
EKG|5122,5125
changes|5126,5133
.|5133,5134
Symptoms|5135,5143
<EOL>|5144,5145
improved|5145,5153
with|5154,5158
duonebs|5159,5166
,|5166,5167
prednisone|5168,5178
and|5179,5182
doxycycline|5183,5194
.|5194,5195
Evaluated|5196,5205
by|5206,5208
<EOL>|5209,5210
_|5210,5211
_|5211,5212
_|5212,5213
and|5214,5217
discharged|5218,5228
to|5229,5231
rehab|5232,5237
facility|5238,5246
for|5247,5250
physical|5251,5259
strengthening|5260,5273
<EOL>|5274,5275
and|5275,5278
respiratory|5279,5290
rehab|5291,5296
.|5296,5297
Discharged|5298,5308
on|5309,5311
home|5312,5316
COPD|5317,5321
meds|5322,5326
and|5327,5330
steroid|5331,5338
<EOL>|5339,5340
taper|5340,5345
and|5346,5349
abx|5350,5353
course|5354,5360
.|5360,5361
<EOL>|5361,5362
<EOL>|5362,5363
#|5363,5364
pAfib|5365,5370
:|5370,5371
currently|5372,5381
rate|5382,5386
well|5387,5391
controlled|5392,5402
.|5402,5403
on|5404,5406
apixaban|5407,5415
<EOL>|5415,5416
<EOL>|5416,5417
-|5417,5418
continued|5419,5428
diltiazam|5429,5438
<EOL>|5438,5439
-|5439,5440
continued|5441,5450
apixaban|5451,5459
<EOL>|5459,5460
-|5460,5461
continued|5462,5471
amiodarone|5472,5482
<EOL>|5482,5483
<EOL>|5483,5484
#|5484,5485
Anemia|5486,5492
:|5492,5493
Fe|5494,5496
def|5497,5500
anemia|5501,5507
on|5508,5510
recent|5511,5517
admission|5518,5527
,|5527,5528
discharged|5529,5539
on|5540,5542
Fe|5543,5545
,|5545,5546
<EOL>|5547,5548
continued|5548,5557
iron|5558,5562
supplement|5563,5573
<EOL>|5573,5574
<EOL>|5574,5575
#|5575,5576
CAD|5577,5580
:|5580,5581
continue|5582,5590
aspirin|5591,5598
,|5598,5599
atorvastatin|5600,5612
<EOL>|5612,5613
#|5613,5614
Constipation|5615,5627
:|5627,5628
continue|5629,5637
home|5638,5642
bowel|5643,5648
reg|5649,5652
<EOL>|5652,5653
#|5653,5654
Anxiety|5655,5662
:|5662,5663
continued|5664,5673
home|5674,5678
meds|5679,5683
<EOL>|5683,5684
<EOL>|5684,5685
TRANSITIONAL|5685,5697
<EOL>|5698,5699
<EOL>|5699,5700
-|5700,5701
Discharged|5702,5712
on|5713,5715
steroid|5716,5723
taper|5724,5729
with|5730,5734
maintenance|5735,5746
dose|5747,5751
of|5752,5754
10mg|5755,5759
<EOL>|5760,5761
daily|5761,5766
until|5767,5772
she|5773,5776
sees|5777,5781
PCP|5782,5785
<EOL>|5785,5786
*|5786,5787
Take|5788,5792
_|5793,5794
_|5794,5795
_|5795,5796
-|5796,5797
<EOL>|5797,5798
<EOL>|5798,5799
-|5799,5800
Doxycycline|5801,5812
100mg|5813,5818
BID|5819,5822
to|5823,5825
_|5826,5827
_|5827,5828
_|5828,5829
<EOL>|5829,5830
<EOL>|5831,5832
Medications|5832,5843
on|5844,5846
Admission|5847,5856
:|5856,5857
<EOL>|5857,5858
The|5858,5861
Preadmission|5862,5874
Medication|5875,5885
list|5886,5890
is|5891,5893
accurate|5894,5902
and|5903,5906
complete|5907,5915
.|5915,5916
<EOL>|5916,5917
1.|5917,5919
Acetaminophen|5920,5933
650|5934,5937
mg|5938,5940
PO|5941,5943
Q6H|5944,5947
:|5947,5948
PRN|5948,5951
pain|5952,5956
<EOL>|5957,5958
2.|5958,5960
Amiodarone|5961,5971
200|5972,5975
mg|5976,5978
PO|5979,5981
DAILY|5982,5987
<EOL>|5988,5989
3.|5989,5991
Apixaban|5992,6000
5|6001,6002
mg|6003,6005
PO|6006,6008
BID|6009,6012
<EOL>|6013,6014
4.|6014,6016
Albuterol|6017,6026
0.083|6027,6032
%|6032,6033
Neb|6034,6037
Soln|6038,6042
1|6043,6044
NEB|6045,6048
IH|6049,6051
Q2H|6052,6055
:|6055,6056
PRN|6056,6059
SOB|6060,6063
<EOL>|6064,6065
5.|6065,6067
Artificial|6068,6078
Tears|6079,6084
_|6085,6086
_|6086,6087
_|6087,6088
DROP|6089,6093
BOTH|6094,6098
EYES|6099,6103
PRN|6104,6107
irritation|6108,6118
<EOL>|6119,6120
6.|6120,6122
Aspirin|6123,6130
81|6131,6133
mg|6134,6136
PO|6137,6139
DAILY|6140,6145
<EOL>|6146,6147
7.|6147,6149
Atorvastatin|6150,6162
10|6163,6165
mg|6166,6168
PO|6169,6171
QPM|6172,6175
<EOL>|6176,6177
8.|6177,6179
Diltiazem|6180,6189
Extended|6190,6198
-|6198,6199
Release|6199,6206
180|6207,6210
mg|6211,6213
PO|6214,6216
BID|6217,6220
<EOL>|6221,6222
9.|6222,6224
Dorzolamide|6225,6236
2|6237,6238
%|6238,6239
Ophth|6240,6245
.|6245,6246
Soln.|6247,6252
1|6253,6254
DROP|6255,6259
BOTH|6260,6264
EYES|6265,6269
BID|6270,6273
<EOL>|6274,6275
10.|6275,6278
Fluticasone|6279,6290
Propionate|6291,6301
NASAL|6302,6307
1|6308,6309
SPRY|6310,6314
NU|6315,6317
BID|6318,6321
<EOL>|6322,6323
11.|6323,6326
Fluticasone|6327,6338
-|6338,6339
Salmeterol|6339,6349
Diskus|6350,6356
(|6357,6358
250|6358,6361
/|6361,6362
50|6362,6364
)|6364,6365
1|6367,6368
INH|6369,6372
IH|6373,6375
BID|6376,6379
<EOL>|6380,6381
12.|6381,6384
Hydrochlorothiazide|6385,6404
50|6405,6407
mg|6408,6410
PO|6411,6413
DAILY|6414,6419
<EOL>|6420,6421
13.|6421,6424
Isosorbide|6425,6435
Mononitrate|6436,6447
(|6448,6449
Extended|6449,6457
Release|6458,6465
)|6465,6466
240|6467,6470
mg|6471,6473
PO|6474,6476
DAILY|6477,6482
<EOL>|6483,6484
14.|6484,6487
Latanoprost|6488,6499
0.005|6500,6505
%|6505,6506
Ophth|6507,6512
.|6512,6513
Soln.|6514,6519
1|6520,6521
DROP|6522,6526
LEFT|6527,6531
EYE|6532,6535
QHS|6536,6539
<EOL>|6540,6541
15.|6541,6544
Lorazepam|6545,6554
0.5|6555,6558
mg|6559,6561
PO|6562,6564
QHS|6565,6568
:|6568,6569
PRN|6569,6572
insomnia|6573,6581
<EOL>|6582,6583
16|6583,6585
.|6585,6586
Multivitamins|6587,6600
W|6601,6602
/|6602,6603
minerals|6603,6611
1|6612,6613
TAB|6614,6617
PO|6618,6620
DAILY|6621,6626
<EOL>|6627,6628
17.|6628,6631
Ranitidine|6632,6642
300|6643,6646
mg|6647,6649
PO|6650,6652
DAILY|6653,6658
<EOL>|6659,6660
18.|6660,6663
Tiotropium|6664,6674
Bromide|6675,6682
1|6683,6684
CAP|6685,6688
IH|6689,6691
DAILY|6692,6697
<EOL>|6698,6699
19|6699,6701
.|6701,6702
Theophylline|6703,6715
SR|6716,6718
200|6719,6722
mg|6723,6725
PO|6726,6728
BID|6729,6732
<EOL>|6733,6734
20|6734,6736
.|6736,6737
Ferrous|6738,6745
Sulfate|6746,6753
325|6754,6757
mg|6758,6760
PO|6761,6763
DAILY|6764,6769
<EOL>|6770,6771
21|6771,6773
.|6773,6774
Docusate|6775,6783
Sodium|6784,6790
100|6791,6794
mg|6795,6797
PO|6798,6800
BID|6801,6804
<EOL>|6805,6806
22.|6806,6809
Polyethylene|6810,6822
Glycol|6823,6829
17|6830,6832
g|6833,6834
PO|6835,6837
DAILY|6838,6843
<EOL>|6844,6845
23|6845,6847
.|6847,6848
Ipratropium|6849,6860
Bromide|6861,6868
Neb|6869,6872
1|6873,6874
NEB|6875,6878
IH|6879,6881
Q6H|6882,6885
:|6885,6886
PRN|6886,6889
SOB|6890,6893
<EOL>|6894,6895
24|6895,6897
.|6897,6898
PredniSONE|6899,6909
30|6910,6912
mg|6913,6915
PO|6916,6918
DAILY|6919,6924
<EOL>|6925,6926
Start|6926,6931
:|6931,6932
_|6933,6934
_|6934,6935
_|6935,6936
,|6936,6937
First|6938,6943
Dose|6944,6948
:|6948,6949
Next|6950,6954
Routine|6955,6962
Administration|6963,6977
Time|6978,6982
<EOL>|6983,6984
This|6984,6988
is|6989,6991
dose|6992,6996
#|6997,6998
1|6999,7000
of|7001,7003
2|7004,7005
tapered|7006,7013
doses|7014,7019
<EOL>|7019,7020
25|7020,7022
.|7022,7023
PredniSONE|7024,7034
20|7035,7037
mg|7038,7040
PO|7041,7043
DAILY|7044,7049
<EOL>|7050,7051
Start|7051,7056
:|7056,7057
After|7058,7063
30|7064,7066
mg|7067,7069
DAILY|7070,7075
tapered|7076,7083
dose|7084,7088
<EOL>|7089,7090
This|7090,7094
is|7095,7097
dose|7098,7102
#|7103,7104
2|7105,7106
of|7107,7109
2|7110,7111
tapered|7112,7119
doses|7120,7125
<EOL>|7125,7126
26|7126,7128
.|7128,7129
PredniSONE|7130,7140
10|7141,7143
mg|7144,7146
PO|7147,7149
DAILY|7150,7155
<EOL>|7156,7157
Start|7157,7162
:|7162,7163
After|7164,7169
last|7170,7174
tapered|7175,7182
dose|7183,7187
completes|7188,7197
<EOL>|7198,7199
This|7199,7203
is|7204,7206
the|7207,7210
maintenance|7211,7222
dose|7223,7227
to|7228,7230
follow|7231,7237
the|7238,7241
last|7242,7246
tapered|7247,7254
dose|7255,7259
<EOL>|7259,7260
<EOL>|7260,7261
<EOL>|7262,7263
Discharge|7263,7272
Medications|7273,7284
:|7284,7285
<EOL>|7285,7286
1.|7286,7288
Acetaminophen|7289,7302
650|7303,7306
mg|7307,7309
PO|7310,7312
Q6H|7313,7316
:|7316,7317
PRN|7317,7320
pain|7321,7325
<EOL>|7326,7327
2.|7327,7329
Amiodarone|7330,7340
200|7341,7344
mg|7345,7347
PO|7348,7350
DAILY|7351,7356
<EOL>|7357,7358
3.|7358,7360
Apixaban|7361,7369
5|7370,7371
mg|7372,7374
PO|7375,7377
BID|7378,7381
<EOL>|7382,7383
4.|7383,7385
Artificial|7386,7396
Tears|7397,7402
_|7403,7404
_|7404,7405
_|7405,7406
DROP|7407,7411
BOTH|7412,7416
EYES|7417,7421
PRN|7422,7425
irritation|7426,7436
<EOL>|7437,7438
5.|7438,7440
Aspirin|7441,7448
81|7449,7451
mg|7452,7454
PO|7455,7457
DAILY|7458,7463
<EOL>|7464,7465
6.|7465,7467
Atorvastatin|7468,7480
10|7481,7483
mg|7484,7486
PO|7487,7489
QPM|7490,7493
<EOL>|7494,7495
7.|7495,7497
Diltiazem|7498,7507
Extended|7508,7516
-|7516,7517
Release|7517,7524
180|7525,7528
mg|7529,7531
PO|7532,7534
BID|7535,7538
<EOL>|7539,7540
8.|7540,7542
Docusate|7543,7551
Sodium|7552,7558
100|7559,7562
mg|7563,7565
PO|7566,7568
BID|7569,7572
<EOL>|7573,7574
9.|7574,7576
Dorzolamide|7577,7588
2|7589,7590
%|7590,7591
Ophth|7592,7597
.|7597,7598
Soln.|7599,7604
1|7605,7606
DROP|7607,7611
BOTH|7612,7616
EYES|7617,7621
BID|7622,7625
<EOL>|7626,7627
10.|7627,7630
Ferrous|7631,7638
Sulfate|7639,7646
325|7647,7650
mg|7651,7653
PO|7654,7656
DAILY|7657,7662
<EOL>|7663,7664
11.|7664,7667
Fluticasone|7668,7679
Propionate|7680,7690
NASAL|7691,7696
1|7697,7698
SPRY|7699,7703
NU|7704,7706
BID|7707,7710
<EOL>|7711,7712
12.|7712,7715
Fluticasone|7716,7727
-|7727,7728
Salmeterol|7728,7738
Diskus|7739,7745
(|7746,7747
250|7747,7750
/|7750,7751
50|7751,7753
)|7753,7754
1|7756,7757
INH|7758,7761
IH|7762,7764
BID|7765,7768
<EOL>|7769,7770
13.|7770,7773
Hydrochlorothiazide|7774,7793
50|7794,7796
mg|7797,7799
PO|7800,7802
DAILY|7803,7808
<EOL>|7809,7810
14.|7810,7813
Isosorbide|7814,7824
Mononitrate|7825,7836
(|7837,7838
Extended|7838,7846
Release|7847,7854
)|7854,7855
240|7856,7859
mg|7860,7862
PO|7863,7865
DAILY|7866,7871
<EOL>|7872,7873
15.|7873,7876
Latanoprost|7877,7888
0.005|7889,7894
%|7894,7895
Ophth|7896,7901
.|7901,7902
Soln.|7903,7908
1|7909,7910
DROP|7911,7915
LEFT|7916,7920
EYE|7921,7924
QHS|7925,7928
<EOL>|7929,7930
16|7930,7932
.|7932,7933
Lorazepam|7934,7943
0.5|7944,7947
mg|7948,7950
PO|7951,7953
QHS|7954,7957
:|7957,7958
PRN|7958,7961
insomnia|7962,7970
<EOL>|7971,7972
17.|7972,7975
Multivitamins|7976,7989
W|7990,7991
/|7991,7992
minerals|7992,8000
1|8001,8002
TAB|8003,8006
PO|8007,8009
DAILY|8010,8015
<EOL>|8016,8017
18.|8017,8020
Polyethylene|8021,8033
Glycol|8034,8040
17|8041,8043
g|8044,8045
PO|8046,8048
DAILY|8049,8054
<EOL>|8055,8056
19|8056,8058
.|8058,8059
Ranitidine|8060,8070
300|8071,8074
mg|8075,8077
PO|8078,8080
DAILY|8081,8086
<EOL>|8087,8088
20|8088,8090
.|8090,8091
Theophylline|8092,8104
SR|8105,8107
200|8108,8111
mg|8112,8114
PO|8115,8117
BID|8118,8121
<EOL>|8122,8123
21|8123,8125
.|8125,8126
Tiotropium|8127,8137
Bromide|8138,8145
1|8146,8147
CAP|8148,8151
IH|8152,8154
DAILY|8155,8160
<EOL>|8161,8162
22.|8162,8165
Albuterol|8166,8175
Inhaler|8176,8183
_|8184,8185
_|8185,8186
_|8186,8187
PUFF|8188,8192
IH|8193,8195
Q6H|8196,8199
:|8199,8200
PRN|8200,8203
SOB|8204,8207
<EOL>|8208,8209
23|8209,8211
.|8211,8212
Ipratropium|8213,8224
Bromide|8225,8232
Neb|8233,8236
1|8237,8238
NEB|8239,8242
IH|8243,8245
Q6H|8246,8249
:|8249,8250
PRN|8250,8253
SOB|8254,8257
<EOL>|8258,8259
24|8259,8261
.|8261,8262
Albuterol|8263,8272
0.083|8273,8278
%|8278,8279
Neb|8280,8283
Soln|8284,8288
1|8289,8290
NEB|8291,8294
IH|8295,8297
Q2H|8298,8301
:|8301,8302
PRN|8302,8305
SOB|8306,8309
<EOL>|8310,8311
25|8311,8313
.|8313,8314
Doxycycline|8315,8326
Hyclate|8327,8334
100|8335,8338
mg|8339,8341
PO|8342,8344
Q12H|8345,8349
Duration|8350,8358
:|8358,8359
2|8360,8361
Days|8362,8366
<EOL>|8367,8368
to|8368,8370
end|8371,8374
_|8375,8376
_|8376,8377
_|8377,8378
<EOL>|8379,8380
26|8380,8382
.|8382,8383
PredniSONE|8384,8394
10|8395,8397
mg|8398,8400
PO|8401,8403
ASDIR|8404,8409
<EOL>|8410,8411
Take|8411,8415
_|8416,8417
_|8417,8418
_|8418,8419
-|8419,8420
<EOL>|8421,8422
Tapered|8422,8429
dose|8430,8434
-|8435,8436
DOWN|8437,8441
<EOL>|8442,8443
<EOL>|8443,8444
<EOL>|8445,8446
Discharge|8446,8455
Disposition|8456,8467
:|8467,8468
<EOL>|8468,8469
Extended|8469,8477
Care|8478,8482
<EOL>|8482,8483
<EOL>|8484,8485
Facility|8485,8493
:|8493,8494
<EOL>|8494,8495
_|8495,8496
_|8496,8497
_|8497,8498
<EOL>|8498,8499
<EOL>|8500,8501
Discharge|8501,8510
Diagnosis|8511,8520
:|8520,8521
<EOL>|8521,8522
Primary|8522,8529
<EOL>|8529,8530
<EOL>|8530,8531
COPD|8531,8535
exacerbation|8536,8548
<EOL>|8548,8549
<EOL>|8549,8550
Secondary|8550,8559
<EOL>|8559,8560
<EOL>|8560,8561
CORONARY|8562,8570
ARTERY|8571,8577
DISEASE|8578,8585
<EOL>|8587,8588
HYPERLIPIDEMIA|8589,8603
<EOL>|8605,8606
HYPERTENSION|8607,8619
<EOL>|8621,8622
OSTEOARTHRITIS|8623,8637
<EOL>|8639,8640
ATRIAL|8641,8647
FIBRILLATION|8648,8660
<EOL>|8662,8663
ANXIETY|8664,8671
<EOL>|8673,8674
GASTROINTESTINAL|8675,8691
BLEEDING|8692,8700
<EOL>|8702,8703
OSTEOARTHRITIS|8704,8718
<EOL>|8720,8721
<EOL>|8721,8722
<EOL>|8723,8724
Mental|8745,8751
Status|8752,8758
:|8758,8759
Clear|8760,8765
and|8766,8769
coherent|8770,8778
.|8778,8779
<EOL>|8779,8780
Level|8780,8785
of|8786,8788
Consciousness|8789,8802
:|8802,8803
Alert|8804,8809
and|8810,8813
interactive|8814,8825
.|8825,8826
<EOL>|8826,8827
Activity|8827,8835
Status|8836,8842
:|8842,8843
Ambulatory|8844,8854
-|8855,8856
requires|8857,8865
assistance|8866,8876
or|8877,8879
aid|8880,8883
(|8884,8885
walker|8885,8891
<EOL>|8892,8893
or|8893,8895
cane|8896,8900
)|8900,8901
.|8901,8902
<EOL>|8902,8903
<EOL>|8903,8904
<EOL>|8905,8906
Dear|8930,8934
_|8935,8936
_|8936,8937
_|8937,8938
,|8938,8939
<EOL>|8939,8940
<EOL>|8940,8941
_|8945,8946
_|8946,8947
_|8947,8948
were|8949,8953
admitted|8954,8962
with|8963,8967
exacerbation|8968,8980
of|8981,8983
your|8984,8988
COPD|8989,8993
.|8993,8994
We|8995,8997
gave|8998,9002
<EOL>|9003,9004
_|9004,9005
_|9005,9006
_|9006,9007
some|9008,9012
treatments|9013,9023
and|9024,9027
_|9028,9029
_|9029,9030
_|9030,9031
improved.|9032,9041
_|9042,9043
_|9043,9044
_|9044,9045
were|9046,9050
evaluated|9051,9060
by|9061,9063
the|9064,9067
<EOL>|9068,9069
physical|9069,9077
therapy|9078,9085
team|9086,9090
who|9091,9094
recommended|9095,9106
a|9107,9108
rehab|9109,9114
stay|9115,9119
for|9120,9123
<EOL>|9124,9125
strengthening|9125,9138
and|9139,9142
improve|9143,9150
your|9151,9155
breathing|9156,9165
.|9165,9166
Please|9167,9173
take|9174,9178
your|9179,9183
<EOL>|9184,9185
medications|9185,9196
as|9197,9199
prescribed|9200,9210
and|9211,9214
follow|9215,9221
up|9222,9224
with|9225,9229
your|9230,9234
providers|9235,9244
.|9244,9245
<EOL>|9245,9246
<EOL>|9246,9247
Sincerely|9247,9256
,|9256,9257
<EOL>|9257,9258
_|9258,9259
_|9259,9260
_|9260,9261
medical|9262,9269
team|9270,9274
<EOL>|9274,9275
<EOL>|9276,9277
Followup|9277,9285
Instructions|9286,9298
:|9298,9299
<EOL>|9299,9300
_|9300,9301
_|9301,9302
_|9302,9303
<EOL>|9303,9304

