 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Procedure|Health Care Activity|SIMPLE_SEGMENT|48,57|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|48,62|false|false|false|C2598112||Admission Date
Finding|Body Substance|SIMPLE_SEGMENT|82,91|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|82,91|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|82,91|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|82,91|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|82,96|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|114,119|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|114,119|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|114,119|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|138,141|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|138,141|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|138,141|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|138,141|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|138,141|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|149,156|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|149,156|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Attribute|Clinical Attribute|SIMPLE_SEGMENT|173,182|false|false|false|C1717415||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|173,182|false|false|false|C0020517|Hypersensitivity|Allergies
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|185,190|false|false|false|C0749139|sulfa|Sulfa
Drug|Antibiotic|SIMPLE_SEGMENT|192,203|false|false|false|C0038760;C0599503;C3536763|Sulfonamide Anti-Infective Agents;Sulfonamide [EPC];Sulfonamides|Sulfonamide
Drug|Organic Chemical|SIMPLE_SEGMENT|192,203|false|false|false|C0038760;C0599503;C3536763|Sulfonamide Anti-Infective Agents;Sulfonamide [EPC];Sulfonamides|Sulfonamide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|192,203|false|false|false|C0038760;C0599503;C3536763|Sulfonamide Anti-Infective Agents;Sulfonamide [EPC];Sulfonamides|Sulfonamide
Drug|Antibiotic|SIMPLE_SEGMENT|204,215|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|Antibiotics
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|219,230|false|false|false|C0161486;C2876539|Poisoning by penicillin;Poisoning by, adverse effect of and underdosing of penicillins|Penicillins
Drug|Antibiotic|SIMPLE_SEGMENT|219,230|false|false|false|C0030842|penicillins|Penicillins
Drug|Organic Chemical|SIMPLE_SEGMENT|219,230|false|false|false|C0030842|penicillins|Penicillins
Finding|Pathologic Function|SIMPLE_SEGMENT|219,230|false|false|false|C0413443|Adverse reaction to penicillins|Penicillins
Finding|Functional Concept|SIMPLE_SEGMENT|233,242|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|251,266|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|257,266|false|false|false|C3864418||Complaint
Finding|Finding|SIMPLE_SEGMENT|257,266|false|false|false|C5441521|Complaint (finding)|Complaint
Anatomy|Body Location or Region|SIMPLE_SEGMENT|268,272|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|SIMPLE_SEGMENT|268,272|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|SIMPLE_SEGMENT|268,272|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Finding|Sign or Symptom|SIMPLE_SEGMENT|268,277|false|false|false|C0007859|Neck Pain|neck pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|273,277|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|273,277|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|273,277|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|SIMPLE_SEGMENT|282,286|false|false|false|C0085639|Falls|fall
Finding|Classification|SIMPLE_SEGMENT|289,294|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|295,303|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|295,303|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|307,325|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|316,325|false|false|false|C0945766||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|316,325|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|316,325|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|316,325|false|false|false|C0184661|Interventional procedure|Procedure
Procedure|Health Care Activity|SIMPLE_SEGMENT|340,349|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Finding|Conceptual Entity|SIMPLE_SEGMENT|352,359|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|352,359|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|352,359|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|352,362|false|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|352,378|false|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|352,378|false|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|363,370|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|363,370|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|363,378|false|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|371,378|false|false|false|C0221423|Illness (finding)|Illness
Finding|Finding|SIMPLE_SEGMENT|384,388|false|false|false|C1706180|Male Gender|male
Finding|Idea or Concept|SIMPLE_SEGMENT|414,422|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Idea or Concept|SIMPLE_SEGMENT|428,438|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|SIMPLE_SEGMENT|428,438|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Anatomy|Body Location or Region|SIMPLE_SEGMENT|442,450|false|false|false|C0027530|Neck|cervical
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|455,463|false|false|false|C0016658|Fracture|fracture
Finding|Body Substance|SIMPLE_SEGMENT|475,482|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|475,482|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|475,482|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|SIMPLE_SEGMENT|545,552|false|false|false|C0596020|Does hit (finding)|hitting
Anatomy|Body Location or Region|SIMPLE_SEGMENT|570,574|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|570,574|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|570,574|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|570,574|false|false|false|C0876917|Procedure on head|head
Finding|Finding|SIMPLE_SEGMENT|589,593|true|false|false|C5890125|Loss (adaptation)|loss
Finding|Finding|SIMPLE_SEGMENT|589,610|true|false|false|C0041657|Unconscious State|loss of consciousness
Finding|Finding|SIMPLE_SEGMENT|597,610|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|consciousness
Finding|Mental Process|SIMPLE_SEGMENT|597,610|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|consciousness
Finding|Body Substance|SIMPLE_SEGMENT|617,624|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|617,624|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|617,624|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Sign or Symptom|SIMPLE_SEGMENT|638,646|false|false|false|C0018681|Headache|headache
Anatomy|Body Location or Region|SIMPLE_SEGMENT|651,655|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|SIMPLE_SEGMENT|651,655|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|SIMPLE_SEGMENT|651,655|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Finding|Sign or Symptom|SIMPLE_SEGMENT|651,660|false|false|false|C0007859|Neck Pain|neck pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|656,660|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|656,660|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|656,660|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Idea or Concept|SIMPLE_SEGMENT|675,683|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Body Substance|SIMPLE_SEGMENT|688,695|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|688,695|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|688,695|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Anatomy|Body Location or Region|SIMPLE_SEGMENT|704,708|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|704,708|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|704,708|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|704,708|false|false|false|C0876917|Procedure on head|head
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|704,719|false|false|false|C0856548|Laceration of head|head laceration
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|709,719|false|false|false|C0043246|Laceration|laceration
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|731,738|false|false|false|C0040405|X-Ray Computed Tomography|CT scan
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|734,738|false|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|760,768|false|false|false|C0016658|Fracture|fracture
Finding|Body Substance|SIMPLE_SEGMENT|774,781|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|774,781|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|774,781|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|SIMPLE_SEGMENT|793,801|true|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|SIMPLE_SEGMENT|793,801|true|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|804,812|false|false|false|C0030554|Paresthesia|tingling
Finding|Sign or Symptom|SIMPLE_SEGMENT|804,812|false|false|false|C2242996|Has tingling sensation|tingling
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|820,824|false|false|false|C0446516|Upper arm|arms
Attribute|Clinical Attribute|SIMPLE_SEGMENT|820,824|false|false|false|C5782111||arms
Disorder|Neoplastic Process|SIMPLE_SEGMENT|820,824|false|false|false|C0206655|Alveolar rhabdomyosarcoma|arms
Finding|Gene or Genome|SIMPLE_SEGMENT|820,824|false|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Finding|Intellectual Product|SIMPLE_SEGMENT|820,824|false|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|828,832|false|false|false|C1140621|Leg|legs
Attribute|Clinical Attribute|SIMPLE_SEGMENT|828,832|false|false|false|C5781420||legs
Finding|Sign or Symptom|SIMPLE_SEGMENT|837,845|true|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|853,857|false|false|false|C0446516|Upper arm|arms
Attribute|Clinical Attribute|SIMPLE_SEGMENT|853,857|true|false|false|C5782111||arms
Disorder|Neoplastic Process|SIMPLE_SEGMENT|853,857|true|false|false|C0206655|Alveolar rhabdomyosarcoma|arms
Finding|Gene or Genome|SIMPLE_SEGMENT|853,857|true|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Finding|Intellectual Product|SIMPLE_SEGMENT|853,857|true|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|861,865|false|false|false|C1140621|Leg|legs
Attribute|Clinical Attribute|SIMPLE_SEGMENT|861,865|false|false|false|C5781420||legs
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|879,884|false|false|false|C0021853|Intestines|bowel
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|879,897|true|false|false|C0015732|Fecal Incontinence|bowel incontinence
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|885,897|true|false|false|C0021167|Incontinence|incontinence
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|901,908|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|901,908|true|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|901,908|true|false|false|C0872388|Procedures on bladder|bladder
Finding|Functional Concept|SIMPLE_SEGMENT|901,918|true|false|false|C0080274|Urinary Retention|bladder retention
Attribute|Clinical Attribute|SIMPLE_SEGMENT|909,918|false|false|false|C1318143|Retention - dental|retention
Finding|Cell Function|SIMPLE_SEGMENT|909,918|false|false|false|C0035280;C0080274;C0333117;C1753315|Retention (Psychology);Retention of content;Urinary Retention;cellular entity retention|retention
Finding|Functional Concept|SIMPLE_SEGMENT|909,918|false|false|false|C0035280;C0080274;C0333117;C1753315|Retention (Psychology);Retention of content;Urinary Retention;cellular entity retention|retention
Finding|Mental Process|SIMPLE_SEGMENT|909,918|false|false|false|C0035280;C0080274;C0333117;C1753315|Retention (Psychology);Retention of content;Urinary Retention;cellular entity retention|retention
Attribute|Clinical Attribute|SIMPLE_SEGMENT|931,941|false|false|false|C2926599||anesthesia
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|931,941|false|false|false|C4049933|Anesthesia substance|anesthesia
Finding|Finding|SIMPLE_SEGMENT|931,941|false|false|false|C0278134;C2219802|Absence of sensation|anesthesia
Finding|Sign or Symptom|SIMPLE_SEGMENT|931,941|false|false|false|C0278134;C2219802|Absence of sensation|anesthesia
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|931,941|false|false|false|C0002903;C0002912|Anesthesia procedures;Dental anesthesia|anesthesia
Anatomy|Body Location or Region|SIMPLE_SEGMENT|954,959|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|954,959|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|954,964|true|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|954,964|true|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|960,964|true|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|960,964|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|960,964|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|966,985|true|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|SIMPLE_SEGMENT|966,985|true|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|SIMPLE_SEGMENT|979,985|false|false|false|C0225386|Breath|breath
Anatomy|Body Location or Region|SIMPLE_SEGMENT|990,999|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|SIMPLE_SEGMENT|990,1004|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1000,1004|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1000,1004|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1000,1004|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|SIMPLE_SEGMENT|1012,1032|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Finding|Functional Concept|SIMPLE_SEGMENT|1017,1024|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|1017,1024|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|1017,1024|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1017,1024|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|1017,1032|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1025,1032|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1025,1032|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1025,1032|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1034,1037|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|PMH
Finding|Gene or Genome|SIMPLE_SEGMENT|1042,1045|false|false|false|C1414538|FBL gene|fib
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1047,1052|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1047,1052|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1047,1052|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Finding|Finding|SIMPLE_SEGMENT|1047,1052|false|false|false|C0750873|COLON PROBLEM|colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1047,1055|false|true|false|C0007102|Malignant tumor of colon|colon ca
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1057,1060|false|false|false|C0020538|Hypertensive disease|htn
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1062,1066|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|copd
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1062,1066|false|false|false|C1647218|COPD pharmacologic substance|copd
Finding|Gene or Genome|SIMPLE_SEGMENT|1062,1066|false|false|false|C1412502|ARCN1 gene|copd
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|1070,1073|false|false|false|C0026760|Multiple Epiphyseal Dysplasia|MED
Finding|Gene or Genome|SIMPLE_SEGMENT|1070,1073|false|false|false|C1413596;C1413597;C1419866;C1456376;C1549978;C4321267;C5781216|COL9A2 gene;COL9A3 gene;COMP gene;COMP wt Allele;Master of Education;SCN8A gene;SCN8A wt Allele|MED
Finding|Intellectual Product|SIMPLE_SEGMENT|1070,1073|false|false|false|C1413596;C1413597;C1419866;C1456376;C1549978;C4321267;C5781216|COL9A2 gene;COL9A3 gene;COMP gene;COMP wt Allele;Master of Education;SCN8A gene;SCN8A wt Allele|MED
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|1075,1083|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|SIMPLE_SEGMENT|1075,1083|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1075,1083|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|SIMPLE_SEGMENT|1085,1096|false|false|false|C0002144|allopurinol|allopurinol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1085,1096|false|false|false|C0002144|allopurinol|allopurinol
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1098,1104|false|false|false|C0678172|Asacol|asacol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1098,1104|false|false|false|C0678172|Asacol|asacol
Drug|Organic Chemical|SIMPLE_SEGMENT|1113,1116|false|false|false|C0033017|Pregnenolone Carbonitrile|pcn
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1113,1116|false|false|false|C0033017|Pregnenolone Carbonitrile|pcn
Finding|Gene or Genome|SIMPLE_SEGMENT|1113,1116|false|false|false|C1418643;C1826553;C4050150|PCNT gene;PLEC gene;PLEC wt Allele|pcn
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1118,1123|false|false|false|C0749139|sulfa|sulfa
Finding|Functional Concept|SIMPLE_SEGMENT|1127,1133|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|1127,1141|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1134,1141|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1134,1141|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1134,1141|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|1147,1153|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|1147,1153|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|1147,1153|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|1147,1153|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|1147,1161|false|false|false|C0241889|Family Medical History|Family History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1154,1161|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1154,1161|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1154,1161|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1168,1176|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|1168,1176|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1168,1176|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|1168,1181|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1168,1181|false|false|false|C0031809|Physical Examination|Physical Exam
Finding|Functional Concept|SIMPLE_SEGMENT|1177,1181|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1177,1181|false|false|false|C0582103|Medical Examination|Exam
Event|Activity|SIMPLE_SEGMENT|1195,1200|false|false|false|C1882509|put - instruction imperative|place
Finding|Functional Concept|SIMPLE_SEGMENT|1195,1200|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|SIMPLE_SEGMENT|1195,1200|false|false|false|C1533810||place
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1216,1219|false|false|false|C1366678;C1433371;C4049852|L-Type Amino Acid Transporter;LAT protein, human;ORC3 protein, human|lat
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1216,1219|false|false|false|C1366678;C1433371;C4049852|L-Type Amino Acid Transporter;LAT protein, human;ORC3 protein, human|lat
Drug|Immunologic Factor|SIMPLE_SEGMENT|1216,1219|false|false|false|C1366678;C1433371;C4049852|L-Type Amino Acid Transporter;LAT protein, human;ORC3 protein, human|lat
Finding|Gene or Genome|SIMPLE_SEGMENT|1216,1219|false|false|false|C1335085;C1425844;C1705279;C2240043|LAT gene;ORC3 gene;ORC3 wt Allele;SPNS1 gene|lat
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1220,1223|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|1220,1223|false|false|false|C3495676|Anorectal Malformations|arm
Finding|Gene or Genome|SIMPLE_SEGMENT|1220,1223|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1220,1223|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|SIMPLE_SEGMENT|1220,1223|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1220,1223|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1227,1232|false|false|false|C0040067|Thumb structure|thumb
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1249,1255|false|false|false|C0016129;C0851278;C4299059|Fingers;Fingers not including thumb;Upper extremity>Finger|finger
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|1258,1261|false|false|false|C0026760|Multiple Epiphyseal Dysplasia|med
Finding|Gene or Genome|SIMPLE_SEGMENT|1258,1261|false|false|false|C1413596;C1413597;C1419866;C1456376;C1549978;C4321267;C5781216|COL9A2 gene;COL9A3 gene;COMP gene;COMP wt Allele;Master of Education;SCN8A gene;SCN8A wt Allele|med
Finding|Intellectual Product|SIMPLE_SEGMENT|1258,1261|false|false|false|C1413596;C1413597;C1419866;C1456376;C1549978;C4321267;C5781216|COL9A2 gene;COL9A3 gene;COMP gene;COMP wt Allele;Master of Education;SCN8A gene;SCN8A wt Allele|med
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1262,1265|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|1262,1265|false|false|false|C3495676|Anorectal Malformations|arm
Finding|Gene or Genome|SIMPLE_SEGMENT|1262,1265|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1262,1265|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|SIMPLE_SEGMENT|1262,1265|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1262,1265|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Finding|Finding|SIMPLE_SEGMENT|1280,1286|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Finding|SIMPLE_SEGMENT|1294,1300|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Finding|SIMPLE_SEGMENT|1308,1314|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Finding|SIMPLE_SEGMENT|1322,1328|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Finding|SIMPLE_SEGMENT|1342,1348|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Finding|SIMPLE_SEGMENT|1356,1362|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Finding|SIMPLE_SEGMENT|1370,1376|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Finding|SIMPLE_SEGMENT|1384,1390|false|false|false|C1554187|Gender Status - Intact|intact
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1399,1404|false|false|false|C0225442;C0460005;C1523842|Trunk of elephant;Trunk structure;dendritic shaft|Trunk
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1399,1404|false|false|false|C0225442;C0460005;C1523842|Trunk of elephant;Trunk structure;dendritic shaft|Trunk
Anatomy|Cell Component|SIMPLE_SEGMENT|1399,1404|false|false|false|C0225442;C0460005;C1523842|Trunk of elephant;Trunk structure;dendritic shaft|Trunk
Finding|Finding|SIMPLE_SEGMENT|1406,1412|false|false|false|C1554187|Gender Status - Intact|intact
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1449,1454|false|false|false|C0018246;C0816951;C4266533|Inguinal part of abdomen;Inguinal region;Pelvis>Groin|Groin
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1456,1460|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|Knee
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1456,1460|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|Knee
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|1456,1460|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|Knee
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1456,1460|false|false|false|C0562271|Examination of knee joint|Knee
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|1466,1469|false|false|false|C0026760|Multiple Epiphyseal Dysplasia|Med
Finding|Gene or Genome|SIMPLE_SEGMENT|1466,1469|false|false|false|C1413596;C1413597;C1419866;C1456376;C1549978;C4321267;C5781216|COL9A2 gene;COL9A3 gene;COMP gene;COMP wt Allele;Master of Education;SCN8A gene;SCN8A wt Allele|Med
Finding|Intellectual Product|SIMPLE_SEGMENT|1466,1469|false|false|false|C1413596;C1413597;C1419866;C1456376;C1549978;C4321267;C5781216|COL9A2 gene;COL9A3 gene;COMP gene;COMP wt Allele;Master of Education;SCN8A gene;SCN8A wt Allele|Med
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1470,1474|false|false|false|C0230445;C1305418|Structure of calf of leg|Calf
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1470,1474|false|false|false|C0230445;C1305418|Structure of calf of leg|Calf
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1477,1480|false|false|false|C0228547|Clava structure (body structure)|Grt
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1481,1484|false|false|false|C0040357;C4299090|Lower extremity>Toes;Toes|Toe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1490,1493|false|false|false|C0040357;C4299090|Lower extremity>Toes;Toes|Toe
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1501,1506|false|false|false|C0039866;C4299091|Lower extremity>Thigh;Thigh structure|Thigh
Finding|Functional Concept|SIMPLE_SEGMENT|1599,1604|false|false|false|C1513492|motor movement|Motor
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1615,1618|false|false|false|C0175372;C3495985|Structure of inferior brachium of corpora quadrigemina;nucleus of the brachium of the inferior colliculus|Bic
Drug|Organic Chemical|SIMPLE_SEGMENT|1615,1618|false|false|false|C0063382|imidazole mustard|Bic
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1615,1618|false|false|false|C0063382|imidazole mustard|Bic
Finding|Gene or Genome|SIMPLE_SEGMENT|1615,1618|false|false|false|C1537811;C2681931|MIR155 gene;MIR155HG gene|Bic
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1615,1618|false|false|false|C5202575|BIC Regimen|Bic
Finding|Gene or Genome|SIMPLE_SEGMENT|1628,1631|false|false|false|C0814229;C3891460|TRI-AAT9-1 gene;Temptation and Restraint Inventory|Tri
Finding|Intellectual Product|SIMPLE_SEGMENT|1628,1631|false|false|false|C0814229;C3891460|TRI-AAT9-1 gene;Temptation and Restraint Inventory|Tri
Finding|Finding|SIMPLE_SEGMENT|1840,1848|false|false|false|C0034935|Babinski Reflex|Babinski
Finding|Classification|SIMPLE_SEGMENT|1851,1859|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|1851,1859|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1851,1859|false|false|false|C5237010|Expression Negative|negative
Finding|Sign or Symptom|SIMPLE_SEGMENT|1861,1867|false|false|false|C0009024|Clonus|Clonus
Finding|Finding|SIMPLE_SEGMENT|1873,1880|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|SIMPLE_SEGMENT|1873,1880|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Intellectual Product|SIMPLE_SEGMENT|1887,1892|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|1893,1901|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1893,1908|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|1893,1908|false|false|false|C0489547|Hospital course|Hospital Course
Finding|Body Substance|SIMPLE_SEGMENT|1910,1917|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1910,1917|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1910,1917|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Finding|SIMPLE_SEGMENT|1946,1953|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Finding|Functional Concept|SIMPLE_SEGMENT|1946,1953|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|1946,1953|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1946,1953|false|false|false|C0543467|Operative Surgical Procedures|Surgery
Event|Occupational Activity|SIMPLE_SEGMENT|1954,1961|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|1954,1961|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Finding|Finding|SIMPLE_SEGMENT|1967,1978|false|false|false|C0478530;C1548358;C1554188;C5890437|Examination and observation for unspecified reason;Observation (finding)|observation
Finding|Idea or Concept|SIMPLE_SEGMENT|1967,1978|false|false|false|C0478530;C1548358;C1554188;C5890437|Examination and observation for unspecified reason;Observation (finding)|observation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1967,1978|false|false|false|C0302523;C0700325;C1964257|Observation - diagnostic procedure;Observation in research;Patient observation|observation
Procedure|Health Care Activity|SIMPLE_SEGMENT|1967,1978|false|false|false|C0302523;C0700325;C1964257|Observation - diagnostic procedure;Observation in research;Patient observation|observation
Procedure|Research Activity|SIMPLE_SEGMENT|1967,1978|false|false|false|C0302523;C0700325;C1964257|Observation - diagnostic procedure;Observation in research;Patient observation|observation
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|1990,1998|false|false|false|C0016658|Fracture|fracture
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2032,2049|false|false|false|C0589110|Postoperative deep vein thrombosis|postoperative DVT
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2046,2049|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2046,2049|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2046,2049|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2046,2061|false|false|false|C0853245|DVT prophylaxis|DVT prophylaxis
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2050,2061|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Drug|Food|SIMPLE_SEGMENT|2064,2068|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|Diet
Finding|Functional Concept|SIMPLE_SEGMENT|2064,2068|false|false|false|C1549512|diet - supply|Diet
Procedure|Health Care Activity|SIMPLE_SEGMENT|2064,2068|false|false|false|C0012159|Diet therapy|Diet
Finding|Body Substance|SIMPLE_SEGMENT|2102,2109|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|2102,2109|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|2102,2109|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|2124,2128|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2124,2128|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|2124,2128|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|2124,2128|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Sign or Symptom|SIMPLE_SEGMENT|2124,2133|false|false|false|C0221776|Oral pain|oral pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2129,2133|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|2129,2133|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2129,2133|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2134,2144|false|false|false|C0013227|Pharmaceutical Preparations|medication
Finding|Intellectual Product|SIMPLE_SEGMENT|2134,2144|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Finding|Finding|SIMPLE_SEGMENT|2146,2154|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|2146,2154|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2146,2154|false|false|false|C0031809|Physical Examination|Physical
Finding|Intellectual Product|SIMPLE_SEGMENT|2146,2162|false|false|false|C1547999|Diagnostic Service Section ID - Physical Therapy|Physical therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2146,2162|false|false|false|C0949766|Physical therapy|Physical therapy
Finding|Finding|SIMPLE_SEGMENT|2155,2162|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|SIMPLE_SEGMENT|2155,2162|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2155,2162|false|false|false|C0087111|Therapeutic procedure|therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2182,2194|false|false|false|C0185112;C2080791|Mobilization (procedure);physical therapy mobilization (treatment)|mobilization
Finding|Finding|SIMPLE_SEGMENT|2202,2210|false|false|false|C4036205|Ambulate|ambulate
Finding|Finding|SIMPLE_SEGMENT|2226,2238|false|false|false|C0857121|Hypertensive (finding)|hypertensive
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2257,2265|false|false|false|C0013227|Pharmaceutical Preparations|Medicine
Procedure|Health Care Activity|SIMPLE_SEGMENT|2257,2273|false|false|false|C0746478|MEDICINE CONSULT|Medicine consult
Procedure|Health Care Activity|SIMPLE_SEGMENT|2266,2273|false|false|false|C0009818|Consultation|consult
Finding|Gene or Genome|SIMPLE_SEGMENT|2331,2334|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2335,2352|false|false|false|C0003364|Antihypertensive Agents|antihypertensives
Finding|Finding|SIMPLE_SEGMENT|2385,2393|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|2385,2393|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|2385,2393|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|2385,2393|false|false|false|C0033095||pressure
Finding|Finding|SIMPLE_SEGMENT|2394,2401|false|false|false|C4036057|Too low|too low
Finding|Finding|SIMPLE_SEGMENT|2398,2401|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|SIMPLE_SEGMENT|2398,2401|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Finding|SIMPLE_SEGMENT|2402,2413|false|false|false|C4036056|Too quickly|too quickly
Finding|Idea or Concept|SIMPLE_SEGMENT|2417,2425|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2417,2432|false|false|false|C0488549||Hospital course
Finding|Finding|SIMPLE_SEGMENT|2417,2432|false|false|false|C0489547|Hospital course|Hospital course
Finding|Idea or Concept|SIMPLE_SEGMENT|2469,2472|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|2469,2472|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Body Substance|SIMPLE_SEGMENT|2477,2486|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|2477,2486|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|2477,2486|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|2477,2486|false|false|false|C0030685|Patient Discharge|discharge
Finding|Body Substance|SIMPLE_SEGMENT|2491,2498|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|2491,2498|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|2491,2498|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|SIMPLE_SEGMENT|2503,2511|false|false|false|C0277797|Apyrexial|afebrile
Finding|Intellectual Product|SIMPLE_SEGMENT|2517,2523|false|false|false|C1547311|Patient Condition Code - Stable|stable
Drug|Food|SIMPLE_SEGMENT|2524,2529|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|vital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2524,2535|false|false|false|C0488614;C0518766|Vital signs|vital signs
Procedure|Health Care Activity|SIMPLE_SEGMENT|2524,2535|false|false|false|C0150404|Taking vital signs|vital signs
Finding|Finding|SIMPLE_SEGMENT|2530,2535|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|2530,2535|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Finding|SIMPLE_SEGMENT|2538,2549|false|false|false|C5546696|Feeling comfortable|comfortable
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|2553,2557|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2553,2557|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|2553,2557|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|2553,2557|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Sign or Symptom|SIMPLE_SEGMENT|2553,2562|false|false|false|C0221776|Oral pain|oral pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2558,2562|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|2558,2562|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2558,2562|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|SIMPLE_SEGMENT|2558,2570|false|false|false|C5548091|Demonstrates adequate pain control|pain control
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2558,2570|false|false|false|C0002766;C1304888|Pain control;Pain management (procedure)|pain control
Drug|Organic Chemical|SIMPLE_SEGMENT|2563,2570|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2563,2570|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|SIMPLE_SEGMENT|2563,2570|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Finding|Conceptual Entity|SIMPLE_SEGMENT|2563,2570|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|SIMPLE_SEGMENT|2563,2570|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|SIMPLE_SEGMENT|2563,2570|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|2588,2600|false|false|false|C0184625||regular diet
Drug|Food|SIMPLE_SEGMENT|2596,2600|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Finding|Functional Concept|SIMPLE_SEGMENT|2596,2600|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|SIMPLE_SEGMENT|2596,2600|false|false|false|C0012159|Diet therapy|diet
Finding|Body Substance|SIMPLE_SEGMENT|2605,2614|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|2605,2614|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|2605,2614|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|2605,2614|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|2605,2626|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2615,2626|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2615,2626|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|2615,2626|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|2631,2644|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2631,2644|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2631,2644|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|SIMPLE_SEGMENT|2659,2662|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2663,2667|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|2663,2667|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2663,2667|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Gene or Genome|SIMPLE_SEGMENT|2669,2673|false|false|false|C1823816|C1orf210 gene|temp
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2669,2673|false|false|false|C0279848|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|temp
Finding|Sign or Symptom|SIMPLE_SEGMENT|2682,2690|false|false|false|C0018681|Headache|headache
Drug|Organic Chemical|SIMPLE_SEGMENT|2695,2706|false|false|false|C0002144|allopurinol|Allopurinol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2695,2706|false|false|false|C0002144|allopurinol|Allopurinol
Drug|Organic Chemical|SIMPLE_SEGMENT|2727,2737|false|false|false|C0127615|mesalamine|Mesalamine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2727,2737|false|false|false|C0127615|mesalamine|Mesalamine
Drug|Organic Chemical|SIMPLE_SEGMENT|2760,2770|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2760,2770|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|2760,2779|false|false|false|C0700548|metoprolol tartrate|Metoprolol Tartrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2760,2779|false|false|false|C0700548|metoprolol tartrate|Metoprolol Tartrate
Drug|Organic Chemical|SIMPLE_SEGMENT|2771,2779|false|false|false|C0039328;C0144544|Tartrates;tartrate|Tartrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2771,2779|false|false|false|C0039328;C0144544|Tartrates;tartrate|Tartrate
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2789,2792|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2789,2792|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2789,2792|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|2789,2792|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|2797,2807|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2797,2807|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|2827,2835|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|SIMPLE_SEGMENT|2827,2835|false|false|false|C0043031|warfarin|Warfarin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2827,2835|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|SIMPLE_SEGMENT|2854,2863|false|false|false|C0030049|oxycodone|OxycoDONE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2854,2863|false|false|false|C0030049|oxycodone|OxycoDONE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2854,2863|false|false|false|C0524222|Oxycodone measurement|OxycoDONE
Finding|Idea or Concept|SIMPLE_SEGMENT|2865,2874|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Finding|Intellectual Product|SIMPLE_SEGMENT|2865,2874|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2865,2882|false|false|false|C1708470|Immediate Release Dosage Form|Immediate Release
Finding|Functional Concept|SIMPLE_SEGMENT|2875,2882|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|2875,2882|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2875,2882|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Finding|Gene or Genome|SIMPLE_SEGMENT|2901,2904|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2905,2909|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|2905,2909|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2905,2909|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|2914,2922|false|false|false|C0012010|diazepam|Diazepam
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2914,2922|false|false|false|C0012010|diazepam|Diazepam
Finding|Gene or Genome|SIMPLE_SEGMENT|2936,2939|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Sign or Symptom|SIMPLE_SEGMENT|2940,2946|false|false|false|C0037763|Spasm|spasms
Finding|Body Substance|SIMPLE_SEGMENT|2951,2960|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|2951,2960|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|2951,2960|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|2951,2960|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2951,2972|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|2951,2972|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2961,2972|false|false|false|C2926604||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|2961,2972|false|false|false|C0184758|Patient disposition|Disposition
Finding|Idea or Concept|SIMPLE_SEGMENT|2974,2978|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|2974,2978|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|2974,2978|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|SIMPLE_SEGMENT|2984,2991|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|2984,2991|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Finding|Intellectual Product|SIMPLE_SEGMENT|2994,3002|false|false|false|C4695111|ADMIN.FACILITY|Facility
Finding|Body Substance|SIMPLE_SEGMENT|3010,3019|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|3010,3019|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|3010,3019|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|3010,3019|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|3010,3029|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3020,3029|false|false|false|C0945731||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|3020,3029|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|3020,3029|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3020,3029|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|3034,3042|false|false|false|C0016658|Fracture|fracture
Finding|Body Substance|SIMPLE_SEGMENT|3045,3054|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|3045,3054|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|3045,3054|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|3045,3054|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3055,3064|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3055,3064|false|false|false|C0012634|Disease|Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|3055,3064|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|3066,3072|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3066,3079|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|3066,3079|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3073,3079|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|3073,3079|false|false|false|C1546481|What subject filter - Status|Status
Finding|Idea or Concept|SIMPLE_SEGMENT|3081,3086|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Finding|SIMPLE_SEGMENT|3091,3099|false|false|false|C4068804|Coherent|coherent
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3101,3123|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|3101,3123|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|3110,3123|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|3110,3123|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3125,3130|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|3125,3130|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3125,3130|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|SIMPLE_SEGMENT|3125,3130|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|3125,3130|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|3125,3130|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|3135,3146|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|3148,3156|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|3148,3156|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|3148,3156|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3157,3163|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|3157,3163|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|SIMPLE_SEGMENT|3165,3175|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|3165,3175|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|3165,3175|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|3165,3175|false|false|false|C1561560|ambulatory encounter|Ambulatory
Finding|Finding|SIMPLE_SEGMENT|3178,3189|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|SIMPLE_SEGMENT|3178,3189|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Body Substance|SIMPLE_SEGMENT|3193,3202|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|3193,3202|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|3193,3202|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|3193,3202|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3193,3215|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|3193,3215|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|3193,3215|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3203,3215|false|false|false|C3263700||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|3203,3215|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Event|Activity|SIMPLE_SEGMENT|3250,3259|false|false|false|C3241922|Operation Activity|operation
Procedure|Machine Activity|SIMPLE_SEGMENT|3250,3259|false|false|false|C0543467;C1880161|Computer Operation;Operative Surgical Procedures|operation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3250,3259|false|false|false|C0543467;C1880161|Computer Operation;Operative Surgical Procedures|operation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3261,3269|false|false|false|C0751437|Adenohypophyseal Diseases|Anterior
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3270,3278|false|false|false|C0027530|Neck|Cervical
Finding|Functional Concept|SIMPLE_SEGMENT|3280,3293|false|false|false|C1965697|Decompression - action (qualifier value)|Decompression
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|3280,3293|false|false|false|C0011117|external decompression|Decompression
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3280,3293|false|false|false|C0021153;C1829459|Decompression;Decompressive incision|Decompression
Finding|Functional Concept|SIMPLE_SEGMENT|3298,3304|false|false|false|C0332466|Fused structure|Fusion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3298,3304|false|false|false|C1293131|Fusion procedure|Fusion
Event|Activity|SIMPLE_SEGMENT|3328,3337|false|false|false|C3241922|Operation Activity|operation
Procedure|Machine Activity|SIMPLE_SEGMENT|3328,3337|false|false|false|C0543467;C1880161|Computer Operation;Operative Surgical Procedures|operation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3328,3337|false|false|false|C0543467;C1880161|Computer Operation;Operative Surgical Procedures|operation
Event|Activity|SIMPLE_SEGMENT|3340,3348|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|3340,3348|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|3340,3348|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3394,3397|false|false|false|C3161851|liquid-based cytology (procedure)|lbs
Finding|Finding|SIMPLE_SEGMENT|3429,3440|false|false|false|C5546696|Feeling comfortable|comfortable
Anatomy|Cell Component|SIMPLE_SEGMENT|3464,3467|false|false|false|C1166663|actomyosin contractile ring|car
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3464,3467|false|false|false|C0406810|Carney Complex|car
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3464,3467|false|false|false|C3539542;C4039583;C5890846|Chimeric antigen receptor;Coxsackievirus and Adenovirus Receptor, human;Extracellular Calcium-Sensing Receptor, Human|car
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3464,3467|false|false|false|C3539542;C4039583;C5890846|Chimeric antigen receptor;Coxsackievirus and Adenovirus Receptor, human;Extracellular Calcium-Sensing Receptor, Human|car
Drug|Immunologic Factor|SIMPLE_SEGMENT|3464,3467|false|false|false|C3539542;C4039583;C5890846|Chimeric antigen receptor;Coxsackievirus and Adenovirus Receptor, human;Extracellular Calcium-Sensing Receptor, Human|car
Finding|Gene or Genome|SIMPLE_SEGMENT|3464,3467|false|false|false|C1413828;C1417827;C1420354;C1547285;C1706434;C1858724;C2239319;C3273602;C3540475;C3811749;C4039583;C5890846;C5890847;C5960871|CASR wt Allele;CXADR gene;CXADR wt Allele;CXADRP1 gene;Car - Mode of Arrival Code;Caronte Gene;Chimeric antigen receptor;Extracellular Calcium-Sensing Receptor, Human;NR1I3 gene;NR1I3 wt Allele;PRKAR1A wt Allele;SPG7 gene;SPG7 wt Allele;TRIM13 wt Allele|car
Finding|Intellectual Product|SIMPLE_SEGMENT|3464,3467|false|false|false|C1413828;C1417827;C1420354;C1547285;C1706434;C1858724;C2239319;C3273602;C3540475;C3811749;C4039583;C5890846;C5890847;C5960871|CASR wt Allele;CXADR gene;CXADR wt Allele;CXADRP1 gene;Car - Mode of Arrival Code;Caronte Gene;Chimeric antigen receptor;Extracellular Calcium-Sensing Receptor, Human;NR1I3 gene;NR1I3 wt Allele;PRKAR1A wt Allele;SPG7 gene;SPG7 wt Allele;TRIM13 wt Allele|car
Finding|Receptor|SIMPLE_SEGMENT|3464,3467|false|false|false|C1413828;C1417827;C1420354;C1547285;C1706434;C1858724;C2239319;C3273602;C3540475;C3811749;C4039583;C5890846;C5890847;C5960871|CASR wt Allele;CXADR gene;CXADR wt Allele;CXADRP1 gene;Car - Mode of Arrival Code;Caronte Gene;Chimeric antigen receptor;Extracellular Calcium-Sensing Receptor, Human;NR1I3 gene;NR1I3 wt Allele;PRKAR1A wt Allele;SPG7 gene;SPG7 wt Allele;TRIM13 wt Allele|car
Finding|Finding|SIMPLE_SEGMENT|3546,3560|false|false|false|C0007237;C0034992|Encounter due to care involving use of rehabilitation procedures;Rehabilitation aspects|Rehabilitation
Finding|Functional Concept|SIMPLE_SEGMENT|3546,3560|false|false|false|C0007237;C0034992|Encounter due to care involving use of rehabilitation procedures;Rehabilitation aspects|Rehabilitation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3546,3560|false|false|false|C0034991|Rehabilitation therapy|Rehabilitation
Finding|Finding|SIMPLE_SEGMENT|3562,3570|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|3562,3570|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|3562,3570|false|false|false|C0031809|Physical Examination|Physical
Finding|Intellectual Product|SIMPLE_SEGMENT|3562,3578|false|false|false|C1547999|Diagnostic Service Section ID - Physical Therapy|Physical Therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3562,3578|false|false|false|C0949766|Physical therapy|Physical Therapy
Finding|Finding|SIMPLE_SEGMENT|3571,3578|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|Therapy
Finding|Functional Concept|SIMPLE_SEGMENT|3571,3578|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|Therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3571,3578|false|false|false|C0087111|Therapeutic procedure|Therapy
Finding|Finding|SIMPLE_SEGMENT|3584,3591|false|false|false|C4035626|3 times|3 times
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3586,3591|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|SIMPLE_SEGMENT|3594,3597|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|3594,3597|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|3618,3622|false|false|false|C0080331|Walking (function)|walk
Finding|Idea or Concept|SIMPLE_SEGMENT|3643,3647|false|false|false|C1552020|Role Class - part|part
Event|Activity|SIMPLE_SEGMENT|3656,3664|false|false|false|C0237820||recovery
Finding|Organism Function|SIMPLE_SEGMENT|3656,3664|false|false|false|C2004454|Recovery - healing process|recovery
Finding|Finding|SIMPLE_SEGMENT|3683,3687|false|false|false|C4281574|Much|much
Finding|Conceptual Entity|SIMPLE_SEGMENT|3723,3732|false|false|false|C0231448;C1880641|Extension;Telephone Extension Number|Extension
Finding|Functional Concept|SIMPLE_SEGMENT|3723,3732|false|false|false|C0231448;C1880641|Extension;Telephone Extension Number|Extension
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|3733,3741|false|false|false|C0015259|Exercise|Exercise
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3733,3741|false|false|false|C1522704|Exercise Pain Management|Exercise
Finding|Idea or Concept|SIMPLE_SEGMENT|3760,3763|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|3760,3763|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3795,3805|false|false|false|C2598159||Swallowing
Finding|Finding|SIMPLE_SEGMENT|3795,3805|false|false|false|C0011167;C0740170;C4281783|Deglutition;Does swallow;Swallowing G-code|Swallowing
Finding|Intellectual Product|SIMPLE_SEGMENT|3795,3805|false|false|false|C0011167;C0740170;C4281783|Deglutition;Does swallow;Swallowing G-code|Swallowing
Finding|Organism Function|SIMPLE_SEGMENT|3795,3805|false|false|false|C0011167;C0740170;C4281783|Deglutition;Does swallow;Swallowing G-code|Swallowing
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3795,3805|false|false|false|C3665547|outcomes otolaryngology swallowing (treatment)|Swallowing
Finding|Finding|SIMPLE_SEGMENT|3807,3817|false|false|false|C1299586|Has difficulty doing (qualifier value)|Difficulty
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3807,3828|true|false|false|C0011168|Deglutition Disorders|Difficulty swallowing
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3818,3828|false|false|false|C2598159||swallowing
Finding|Finding|SIMPLE_SEGMENT|3818,3828|false|false|false|C0011167;C0740170;C4281783|Deglutition;Does swallow;Swallowing G-code|swallowing
Finding|Intellectual Product|SIMPLE_SEGMENT|3818,3828|false|false|false|C0011167;C0740170;C4281783|Deglutition;Does swallow;Swallowing G-code|swallowing
Finding|Organism Function|SIMPLE_SEGMENT|3818,3828|false|false|false|C0011167;C0740170;C4281783|Deglutition;Does swallow;Swallowing G-code|swallowing
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3818,3828|false|false|false|C3665547|outcomes otolaryngology swallowing (treatment)|swallowing
Finding|Gene or Genome|SIMPLE_SEGMENT|3857,3861|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Intellectual Product|SIMPLE_SEGMENT|3857,3861|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Finding|SIMPLE_SEGMENT|3865,3872|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|3865,3872|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|3865,3872|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3865,3872|false|false|false|C0543467|Operative Surgical Procedures|surgery
Finding|Finding|SIMPLE_SEGMENT|3899,3903|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|3899,3903|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|3899,3903|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|3925,3930|false|false|false|C0005658|bite injury|bites
Finding|Organism Function|SIMPLE_SEGMENT|4026,4034|false|false|false|C0026649|Movement|movement
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4044,4048|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|SIMPLE_SEGMENT|4044,4048|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|SIMPLE_SEGMENT|4044,4048|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4091,4099|false|false|false|C0027530|Neck|Cervical
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4109,4113|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|SIMPLE_SEGMENT|4109,4113|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|SIMPLE_SEGMENT|4109,4113|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4114,4119|false|false|false|C1828220|Application of brace (procedure)|Brace
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4142,4147|false|false|false|C1828220|Application of brace (procedure)|brace
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4156,4161|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Functional Concept|SIMPLE_SEGMENT|4173,4179|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|4173,4179|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|SIMPLE_SEGMENT|4173,4182|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|SIMPLE_SEGMENT|4173,4182|false|false|false|C1522577|follow-up|follow-up
Event|Activity|SIMPLE_SEGMENT|4183,4194|false|false|false|C0003629|Appointments|appointment
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|4254,4267|false|false|false|C2937301|take a shower|take a shower
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|4282,4288|false|false|false|C0026597|Motion|motion
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4297,4301|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|SIMPLE_SEGMENT|4297,4301|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|SIMPLE_SEGMENT|4297,4301|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Event|Activity|SIMPLE_SEGMENT|4327,4332|false|false|false|C1882509|put - instruction imperative|Place
Finding|Functional Concept|SIMPLE_SEGMENT|4327,4332|false|false|false|C1704765|Place - dosing instruction imperative|Place
Procedure|Health Care Activity|SIMPLE_SEGMENT|4327,4332|false|false|false|C1533810||Place
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4358,4362|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|SIMPLE_SEGMENT|4358,4362|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|SIMPLE_SEGMENT|4358,4362|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|4395,4400|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|Wound
Finding|Body Substance|SIMPLE_SEGMENT|4395,4400|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|Wound
Finding|Functional Concept|SIMPLE_SEGMENT|4395,4400|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|Wound
Finding|Intellectual Product|SIMPLE_SEGMENT|4395,4400|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|Wound
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4395,4405|false|false|false|C0886052;C1272654|Wound care management;wound care|Wound Care
Event|Activity|SIMPLE_SEGMENT|4401,4405|false|false|false|C1947933|care activity|Care
Finding|Finding|SIMPLE_SEGMENT|4401,4405|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|SIMPLE_SEGMENT|4401,4405|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|4415,4425|false|false|false|C0043246|Laceration|laceration
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4429,4434|false|false|false|C0036270|Scalp structure|scalp
Finding|Body Substance|SIMPLE_SEGMENT|4439,4447|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|SIMPLE_SEGMENT|4439,4447|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4439,4447|false|false|false|C0013103|Drainage procedure|drainage
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4448,4455|false|false|false|C0041834|Erythema|redness
Finding|Finding|SIMPLE_SEGMENT|4448,4455|false|false|false|C0332575|Redness|redness
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4464,4467|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|4464,4467|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4464,4467|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4464,4467|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|4464,4467|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|4464,4467|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|4464,4467|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4464,4467|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|4464,4467|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|4464,4467|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Idea or Concept|SIMPLE_SEGMENT|4535,4539|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|4535,4539|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|4535,4539|false|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4540,4551|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4540,4551|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|SIMPLE_SEGMENT|4540,4551|false|false|false|C4284232|Medications|medications
Finding|Functional Concept|SIMPLE_SEGMENT|4580,4590|false|false|false|C1524062|Additional|Additional
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4591,4602|false|false|true|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4591,4602|false|false|true|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|4591,4602|false|false|true|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|4606,4613|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4606,4613|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|SIMPLE_SEGMENT|4606,4613|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Finding|Conceptual Entity|SIMPLE_SEGMENT|4606,4613|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|SIMPLE_SEGMENT|4606,4613|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|SIMPLE_SEGMENT|4606,4613|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4620,4624|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|4620,4624|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|4620,4624|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Idea or Concept|SIMPLE_SEGMENT|4653,4659|false|false|false|C0807726|refill|refill
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|4663,4671|false|false|false|C0027415|Narcotics|narcotic
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4663,4671|false|false|false|C0027415|Narcotics|narcotic
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4673,4686|false|false|false|C2741652||prescriptions
Procedure|Health Care Activity|SIMPLE_SEGMENT|4673,4686|false|false|false|C0033080|Prescription (procedure)|prescriptions
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4691,4695|false|false|false|C0270724|Infantile Neuroaxonal Dystrophy|plan
Finding|Functional Concept|SIMPLE_SEGMENT|4691,4695|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Intellectual Product|SIMPLE_SEGMENT|4691,4695|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Mental Process|SIMPLE_SEGMENT|4691,4695|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Idea or Concept|SIMPLE_SEGMENT|4745,4749|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|4745,4749|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|4745,4749|false|false|false|C1553498|home health encounter|home
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|4828,4836|false|false|false|C0027415|Narcotics|narcotic
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4828,4836|false|false|false|C0027415|Narcotics|narcotic
Drug|Organic Chemical|SIMPLE_SEGMENT|4838,4847|false|false|false|C0722364|Oxycontin|oxycontin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4838,4847|false|false|false|C0722364|Oxycontin|oxycontin
Drug|Organic Chemical|SIMPLE_SEGMENT|4849,4858|false|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4849,4858|false|false|false|C0030049|oxycodone|oxycodone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4849,4858|false|false|false|C0524222|Oxycodone measurement|oxycodone
Drug|Organic Chemical|SIMPLE_SEGMENT|4861,4869|false|false|false|C0086787|Percocet|percocet
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4861,4869|false|false|false|C0086787|Percocet|percocet
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4871,4884|false|false|false|C2741652||prescriptions
Procedure|Health Care Activity|SIMPLE_SEGMENT|4871,4884|false|false|false|C0033080|Prescription (procedure)|prescriptions
Finding|Intellectual Product|SIMPLE_SEGMENT|4892,4900|false|false|false|C1547997;C3244303|Diagnostic Service Section ID - Pharmacy;Pharmacy domain|pharmacy
Procedure|Health Care Activity|SIMPLE_SEGMENT|4892,4900|false|false|false|C0031321|Pharmaceutical Services|pharmacy
Finding|Functional Concept|SIMPLE_SEGMENT|4907,4915|false|false|false|C0332287;C1883712|Add - instruction imperative;In addition to|addition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4951,4955|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|4951,4955|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|4951,4955|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4956,4967|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4956,4967|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|SIMPLE_SEGMENT|4956,4967|false|false|false|C4284232|Medications|medications
Finding|Finding|SIMPLE_SEGMENT|4998,5005|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|4998,5005|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|4998,5005|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4998,5005|false|false|false|C0543467|Operative Surgical Procedures|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|5009,5015|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|Follow
Finding|Intellectual Product|SIMPLE_SEGMENT|5009,5015|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|Follow
Finding|Finding|SIMPLE_SEGMENT|5009,5018|false|false|false|C0589120|Follow-up status|Follow up
Procedure|Health Care Activity|SIMPLE_SEGMENT|5009,5018|false|false|false|C1522577|follow-up|Follow up
Finding|Idea or Concept|SIMPLE_SEGMENT|5037,5043|false|false|false|C1549636|Address type - Office|office
Event|Activity|SIMPLE_SEGMENT|5060,5071|false|false|false|C0003629|Appointments|appointment
Finding|Idea or Concept|SIMPLE_SEGMENT|5104,5107|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|5104,5107|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Activity|SIMPLE_SEGMENT|5116,5125|false|false|false|C3241922|Operation Activity|operation
Procedure|Machine Activity|SIMPLE_SEGMENT|5116,5125|false|false|false|C0543467;C1880161|Computer Operation;Operative Surgical Procedures|operation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5116,5125|false|false|false|C0543467;C1880161|Computer Operation;Operative Surgical Procedures|operation
Finding|Intellectual Product|SIMPLE_SEGMENT|5172,5176|false|false|false|C1561540|Transaction counts and value totals - week|week
Finding|Social Behavior|SIMPLE_SEGMENT|5177,5182|false|false|false|C0545082|Visit|visit
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5202,5210|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|5202,5210|false|false|false|C0332803|Surgical wound|incision
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5202,5210|false|false|false|C0184898|Surgical incisions|incision
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5217,5225|false|false|false|C0168634|BaseLine dental cement|baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|5217,5225|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|5227,5233|false|false|false|C0043309|Roentgen Rays|x rays
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5227,5233|false|false|false|C1306645|Plain x-ray|x rays
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|5229,5233|false|false|false|C0851346|Radiation|rays
Finding|Intellectual Product|SIMPLE_SEGMENT|5269,5273|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Idea or Concept|SIMPLE_SEGMENT|5302,5305|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|5302,5305|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Activity|SIMPLE_SEGMENT|5313,5322|false|false|false|C3241922|Operation Activity|operation
Procedure|Machine Activity|SIMPLE_SEGMENT|5313,5322|false|false|false|C0543467;C1880161|Computer Operation;Operative Surgical Procedures|operation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5313,5322|false|false|false|C0543467;C1880161|Computer Operation;Operative Surgical Procedures|operation
Finding|Finding|SIMPLE_SEGMENT|5333,5337|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|5333,5337|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|5333,5337|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|5346,5357|false|false|false|C0750501|most likely|most likely
Finding|Finding|SIMPLE_SEGMENT|5351,5357|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|5351,5357|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5365,5372|false|false|false|C1525443|W flexion|Flexion
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5365,5372|false|false|false|C0231452||Flexion
Finding|Conceptual Entity|SIMPLE_SEGMENT|5373,5382|false|false|false|C0231448;C1880641|Extension;Telephone Extension Number|Extension
Finding|Functional Concept|SIMPLE_SEGMENT|5373,5382|false|false|false|C0231448;C1880641|Extension;Telephone Extension Number|Extension
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5383,5389|false|false|false|C0885876|X-rays, Homeopathic Preparations|X-rays
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|5383,5389|false|false|false|C0043309|Roentgen Rays|X-rays
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5383,5389|false|false|false|C0043299;C1306645|Diagnostic radiologic examination;Plain x-ray|X-rays
Finding|Intellectual Product|SIMPLE_SEGMENT|5395,5400|false|false|false|C4050225|Often - answer to question|often
Finding|Finding|SIMPLE_SEGMENT|5401,5405|false|false|false|C1299581|Able (qualifier value)|able
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5424,5428|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Finding|Intellectual Product|SIMPLE_SEGMENT|5471,5475|false|false|false|C1561540|Transaction counts and value totals - week|week
Finding|Idea or Concept|SIMPLE_SEGMENT|5496,5502|false|false|false|C1549636|Address type - Office|office
Finding|Finding|SIMPLE_SEGMENT|5517,5522|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|5517,5522|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Intellectual Product|SIMPLE_SEGMENT|5529,5536|false|false|false|C0542560|Academic degree|degrees
Finding|Body Substance|SIMPLE_SEGMENT|5550,5558|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|SIMPLE_SEGMENT|5550,5558|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5550,5558|false|false|false|C0013103|Drainage procedure|drainage
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|5569,5574|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Finding|Body Substance|SIMPLE_SEGMENT|5569,5574|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|SIMPLE_SEGMENT|5569,5574|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|SIMPLE_SEGMENT|5569,5574|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Finding|SIMPLE_SEGMENT|5600,5608|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|5600,5608|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|5600,5608|false|false|false|C0031809|Physical Examination|Physical
Finding|Intellectual Product|SIMPLE_SEGMENT|5600,5616|false|false|false|C1547999|Diagnostic Service Section ID - Physical Therapy|Physical Therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5600,5616|false|false|false|C0949766|Physical therapy|Physical Therapy
Finding|Finding|SIMPLE_SEGMENT|5609,5616|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|Therapy
Finding|Functional Concept|SIMPLE_SEGMENT|5609,5616|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|Therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5609,5616|false|false|false|C0087111|Therapeutic procedure|Therapy
Event|Activity|SIMPLE_SEGMENT|5618,5626|false|false|false|C0441655|Activities|activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|5618,5626|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Finding|Finding|SIMPLE_SEGMENT|5618,5626|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Finding|Finding|SIMPLE_SEGMENT|5649,5658|false|false|false|C0682295|Full-time employment (finding)|full time
Finding|Finding|SIMPLE_SEGMENT|5654,5658|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|5654,5658|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|5654,5658|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Functional Concept|SIMPLE_SEGMENT|5680,5690|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|5680,5690|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|5680,5690|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|5680,5690|false|false|false|C1561560|ambulatory encounter|ambulatory
Phenomenon|Human-caused Phenomenon or Process|SIMPLE_SEGMENT|5713,5719|false|true|false|C0036043|Safety|safety
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5724,5731|false|false|false|C0011119|Decompression Sickness|bending
Finding|Finding|SIMPLE_SEGMENT|5724,5731|false|false|false|C0700231;C2584296|Bending - Changing basic body position;Does bend|bending
Finding|Physiologic Function|SIMPLE_SEGMENT|5724,5731|false|false|false|C0700231;C2584296|Bending - Changing basic body position;Does bend|bending
Finding|Pathologic Function|SIMPLE_SEGMENT|5732,5740|true|false|false|C0040480;C1265748|Musculoskeletal torsion (function);Torsion (malposition)|twisting
Finding|Physiologic Function|SIMPLE_SEGMENT|5732,5740|true|false|false|C0040480;C1265748|Musculoskeletal torsion (function);Torsion (malposition)|twisting
Finding|Conceptual Entity|SIMPLE_SEGMENT|5759,5768|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|Treatment
Finding|Functional Concept|SIMPLE_SEGMENT|5759,5768|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|Treatment
Procedure|Health Care Activity|SIMPLE_SEGMENT|5759,5768|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|Treatment
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5759,5768|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|Treatment
Finding|Intellectual Product|SIMPLE_SEGMENT|5769,5778|false|false|false|C3898838;C4321352|Frequency;How Often|Frequency
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|5780,5787|false|false|false|C0728873|Monitor brand of insecticide|monitor
Drug|Organic Chemical|SIMPLE_SEGMENT|5780,5787|false|false|false|C0728873|Monitor brand of insecticide|monitor
Anatomy|Body System|SIMPLE_SEGMENT|5788,5792|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5788,5792|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5788,5792|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Finding|Body Substance|SIMPLE_SEGMENT|5788,5792|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|SIMPLE_SEGMENT|5788,5792|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5796,5800|false|false|false|C0008114|Chin|chin
Procedure|Health Care Activity|SIMPLE_SEGMENT|5796,5800|false|false|false|C2226982|examination of chin|chin
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5805,5817|false|false|false|C0230005|Occipital region|back of head
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5813,5817|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5813,5817|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5813,5817|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5813,5817|false|false|false|C0876917|Procedure on head|head
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|5822,5831|false|false|false|C1265875|Disintegration (morphologic abnormality)|breakdown
Finding|Organism Function|SIMPLE_SEGMENT|5822,5831|false|false|false|C0699900|Catabolism|breakdown
Procedure|Health Care Activity|SIMPLE_SEGMENT|5846,5854|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5855,5867|false|false|false|C3263700||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|5855,5867|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

