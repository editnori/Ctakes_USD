 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|26,30
No|31,33
:|33,34
_|37,38
_|38,39
_|39,40
<EOL>|40,41
<EOL>|42,43
Admission|43,52
Date|53,57
:|57,58
_|60,61
_|61,62
_|62,63
Discharge|77,86
Date|87,91
:|91,92
_|95,96
_|96,97
_|97,98
<EOL>|98,99
<EOL>|100,101
Date|101,105
of|106,108
Birth|109,114
:|114,115
_|117,118
_|118,119
_|119,120
Sex|133,136
:|136,137
M|140,141
<EOL>|141,142
<EOL>|143,144
Service|144,151
:|151,152
MEDICINE|153,161
<EOL>|161,162
<EOL>|163,164
Allergies|164,173
:|173,174
<EOL>|175,176
Corgard|176,183
/|184,185
_|186,187
_|187,188
_|188,189
<EOL>|189,190
<EOL>|191,192
Attending|192,201
:|201,202
_|203,204
_|204,205
_|205,206
.|206,207
<EOL>|207,208
<EOL>|209,210
Major|210,215
Surgical|216,224
or|225,227
Invasive|228,236
Procedure|237,246
:|246,247
<EOL>|247,248
None|248,252
<EOL>|252,253
<EOL>|253,254
attach|254,260
<EOL>|260,261
<EOL>|262,263
Pertinent|263,272
Results|273,280
:|280,281
<EOL>|281,282
ADMISSION|282,291
LABS|292,296
:|296,297
<EOL>|297,298
=|298,299
=|299,300
=|300,301
=|301,302
=|302,303
=|303,304
=|304,305
=|305,306
=|306,307
=|307,308
=|308,309
=|309,310
=|310,311
=|311,312
=|312,313
<EOL>|313,314
_|314,315
_|315,316
_|316,317
12|318,320
:|320,321
48AM|321,325
BLOOD|326,331
WBC|332,335
-|335,336
10|336,338
.|338,339
3|339,340
*|340,341
RBC|342,345
-|345,346
3|346,347
.|347,348
71|348,350
*|350,351
Hgb|352,355
-|355,356
10|356,358
.|358,359
6|359,360
*|360,361
Hct|362,365
-|365,366
36|366,368
.|368,369
6|369,370
*|370,371
<EOL>|372,373
MCV|373,376
-|376,377
99|377,379
*|379,380
MCH|381,384
-|384,385
28.6|385,389
MCHC|390,394
-|394,395
29|395,397
.|397,398
0|398,399
*|399,400
RDW|401,404
-|404,405
18|405,407
.|407,408
6|408,409
*|409,410
RDWSD|411,416
-|416,417
55|417,419
.|419,420
8|420,421
*|421,422
Plt|423,426
_|427,428
_|428,429
_|429,430
<EOL>|430,431
_|431,432
_|432,433
_|433,434
12|435,437
:|437,438
48AM|438,442
BLOOD|443,448
_|449,450
_|450,451
_|451,452
PTT|453,456
-|456,457
82|457,459
.|459,460
4|460,461
*|461,462
_|463,464
_|464,465
_|465,466
<EOL>|466,467
_|467,468
_|468,469
_|469,470
12|471,473
:|473,474
48AM|474,478
BLOOD|479,484
Glucose|485,492
-|492,493
128|493,496
*|496,497
UreaN|498,503
-|503,504
47|504,506
*|506,507
Creat|508,513
-|513,514
2|514,515
.|515,516
2|516,517
*|517,518
Na|519,521
-|521,522
144|522,525
<EOL>|526,527
K|527,528
-|528,529
3.8|529,532
Cl|533,535
-|535,536
105|536,539
HCO3|540,544
-|544,545
22|545,547
AnGap|548,553
-|553,554
17|554,556
<EOL>|556,557
_|557,558
_|558,559
_|559,560
12|561,563
:|563,564
48AM|564,568
BLOOD|569,574
ALT|575,578
-|578,579
75|579,581
*|581,582
AST|583,586
-|586,587
55|587,589
*|589,590
AlkPhos|591,598
-|598,599
150|599,602
*|602,603
TotBili|604,611
-|611,612
1.1|612,615
<EOL>|615,616
_|616,617
_|617,618
_|618,619
12|620,622
:|622,623
48AM|623,627
BLOOD|628,633
_|634,635
_|635,636
_|636,637
<EOL>|637,638
_|638,639
_|639,640
_|640,641
12|642,644
:|644,645
48AM|645,649
BLOOD|650,655
Calcium|656,663
-|663,664
9.2|664,667
Phos|668,672
-|672,673
4.0|673,676
Mg|677,679
-|679,680
2.3|680,683
<EOL>|683,684
_|684,685
_|685,686
_|686,687
01|688,690
:|690,691
19AM|691,695
BLOOD|696,701
_|702,703
_|703,704
_|704,705
pO2|706,709
-|709,710
59|710,712
*|712,713
pCO2|714,718
-|718,719
42|719,721
pH|722,724
-|724,725
7|725,726
.|726,727
34|727,729
*|729,730
<EOL>|731,732
calTCO2|732,739
-|739,740
24|740,742
Base|743,747
XS|748,750
-|750,751
-|751,752
2|752,753
<EOL>|753,754
<EOL>|754,755
RELEVANT|755,763
LABS|764,768
:|768,769
<EOL>|769,770
=|770,771
=|771,772
=|772,773
=|773,774
=|774,775
=|775,776
=|776,777
=|777,778
=|778,779
=|779,780
=|780,781
=|781,782
=|782,783
=|783,784
<EOL>|784,785
_|785,786
_|786,787
_|787,788
12|789,791
:|791,792
48AM|792,796
BLOOD|797,802
_|803,804
_|804,805
_|805,806
<EOL>|806,807
<EOL>|807,808
IMAGING|808,815
:|815,816
<EOL>|816,817
=|817,818
=|818,819
=|819,820
=|820,821
=|821,822
=|822,823
=|823,824
=|824,825
<EOL>|825,826
CXR|826,829
:|829,830
_|831,832
_|832,833
_|833,834
<EOL>|834,835
No|835,837
comparison|838,848
.|848,849
The|851,854
lung|855,859
volumes|860,867
are|868,871
low|872,875
.|875,876
Moderate|878,886
cardiomegaly|887,899
<EOL>|900,901
is|901,903
present|904,911
.|911,912
Normal|914,920
alignment|921,930
of|931,933
the|934,937
sternal|938,945
wires|946,951
after|952,957
CABG|958,962
.|962,963
<EOL>|965,966
Mild|966,970
bilateral|971,980
pleural|981,988
effusions|989,998
.|998,999
Signs|1001,1006
of|1007,1009
moderate|1010,1018
pulmonary|1019,1028
<EOL>|1029,1030
edema|1030,1035
.|1035,1036
Retrocardiac|1038,1050
atelectasis|1051,1062
,|1062,1063
no|1064,1066
evidence|1067,1075
of|1076,1078
pneumonia|1079,1088
.|1088,1089
<EOL>|1090,1091
<EOL>|1091,1092
CXR|1092,1095
:|1095,1096
_|1097,1098
_|1098,1099
_|1099,1100
<EOL>|1100,1101
There|1101,1106
are|1107,1110
stable|1111,1117
postsurgical|1118,1130
changes|1131,1138
following|1139,1148
wedge|1149,1154
resection|1155,1164
<EOL>|1165,1166
the|1166,1169
right|1170,1175
<EOL>|1176,1177
lower|1177,1182
lobe|1183,1187
.|1187,1188
Small|1190,1195
bilateral|1196,1205
effusions|1206,1215
right|1216,1221
greater|1222,1229
than|1230,1234
left|1235,1239
<EOL>|1240,1241
are|1241,1244
unchanged|1245,1254
.|1254,1255
Cardiomediastinal|1256,1273
silhouette|1274,1284
is|1285,1287
stable|1288,1294
.|1294,1295
There|1297,1302
is|1303,1305
<EOL>|1306,1307
moderate|1307,1315
cardiomegaly|1316,1328
.|1328,1329
No|1331,1333
pneumothorax|1334,1346
.|1346,1347
Mild|1349,1353
pulmonary|1354,1363
edema|1364,1369
<EOL>|1370,1371
is|1371,1373
unchanged|1374,1383
.|1383,1384
<EOL>|1385,1386
<EOL>|1386,1387
DISCARHGE|1387,1396
LABS|1397,1401
:|1401,1402
<EOL>|1402,1403
=|1403,1404
=|1404,1405
=|1405,1406
=|1406,1407
=|1407,1408
=|1408,1409
=|1409,1410
=|1410,1411
=|1411,1412
=|1412,1413
=|1413,1414
=|1414,1415
=|1415,1416
=|1416,1417
=|1417,1418
=|1418,1419
=|1419,1420
=|1420,1421
=|1421,1422
<EOL>|1422,1423
_|1423,1424
_|1424,1425
_|1425,1426
08|1427,1429
:|1429,1430
00AM|1430,1434
BLOOD|1435,1440
WBC|1441,1444
-|1444,1445
5.4|1445,1448
RBC|1449,1452
-|1452,1453
3|1453,1454
.|1454,1455
54|1455,1457
*|1457,1458
Hgb|1459,1462
-|1462,1463
10|1463,1465
.|1465,1466
3|1466,1467
*|1467,1468
Hct|1469,1472
-|1472,1473
34|1473,1475
.|1475,1476
1|1476,1477
*|1477,1478
<EOL>|1479,1480
MCV|1480,1483
-|1483,1484
96|1484,1486
MCH|1487,1490
-|1490,1491
29.1|1491,1495
MCHC|1496,1500
-|1500,1501
30|1501,1503
.|1503,1504
2|1504,1505
*|1505,1506
RDW|1507,1510
-|1510,1511
19|1511,1513
.|1513,1514
0|1514,1515
*|1515,1516
RDWSD|1517,1522
-|1522,1523
65|1523,1525
.|1525,1526
7|1526,1527
*|1527,1528
Plt|1529,1532
_|1533,1534
_|1534,1535
_|1535,1536
<EOL>|1536,1537
_|1537,1538
_|1538,1539
_|1539,1540
08|1541,1543
:|1543,1544
00AM|1544,1548
BLOOD|1549,1554
Glucose|1555,1562
-|1562,1563
94|1563,1565
UreaN|1566,1571
-|1571,1572
44|1572,1574
*|1574,1575
Creat|1576,1581
-|1581,1582
2|1582,1583
.|1583,1584
0|1584,1585
*|1585,1586
Na|1587,1589
-|1589,1590
140|1590,1593
<EOL>|1594,1595
K|1595,1596
-|1596,1597
3.6|1597,1600
Cl|1601,1603
-|1603,1604
99|1604,1606
HCO3|1607,1611
-|1611,1612
27|1612,1614
AnGap|1615,1620
-|1620,1621
14|1621,1623
<EOL>|1623,1624
_|1624,1625
_|1625,1626
_|1626,1627
08|1628,1630
:|1630,1631
00AM|1631,1635
BLOOD|1636,1641
ALT|1642,1645
-|1645,1646
38|1646,1648
AST|1649,1652
-|1652,1653
46|1653,1655
*|1655,1656
LD|1657,1659
(|1659,1660
LDH|1660,1663
)|1663,1664
-|1664,1665
198|1665,1668
AlkPhos|1669,1676
-|1676,1677
108|1677,1680
<EOL>|1681,1682
TotBili|1682,1689
-|1689,1690
0.5|1690,1693
<EOL>|1693,1694
_|1694,1695
_|1695,1696
_|1696,1697
08|1698,1700
:|1700,1701
00AM|1701,1705
BLOOD|1706,1711
Calcium|1712,1719
-|1719,1720
9.0|1720,1723
Phos|1724,1728
-|1728,1729
3.5|1729,1732
Mg|1733,1735
-|1735,1736
2.3|1736,1739
<EOL>|1739,1740
<EOL>|1741,1742
Brief|1742,1747
Hospital|1748,1756
Course|1757,1763
:|1763,1764
<EOL>|1764,1765
TRANSITIONAL|1765,1777
ISSUES|1778,1784
:|1784,1785
<EOL>|1785,1786
=|1786,1787
=|1787,1788
=|1788,1789
=|1789,1790
=|1790,1791
=|1791,1792
=|1792,1793
=|1793,1794
=|1794,1795
=|1795,1796
=|1796,1797
=|1797,1798
=|1798,1799
=|1799,1800
=|1800,1801
=|1801,1802
=|1802,1803
=|1803,1804
=|1804,1805
=|1805,1806
<EOL>|1806,1807
[|1807,1808
]|1808,1809
Consider|1810,1818
discontinuing|1819,1832
amiodarone|1833,1843
given|1844,1849
persistence|1850,1861
of|1862,1864
AF|1865,1867
<EOL>|1868,1869
despite|1869,1876
this|1877,1881
medication|1882,1892
<EOL>|1892,1893
[|1893,1894
]|1894,1895
Consider|1896,1904
starting|1905,1913
beta|1914,1918
blocker|1919,1926
,|1926,1927
if|1928,1930
BP|1931,1933
is|1934,1936
able|1937,1941
to|1942,1944
tolerate|1945,1953
.|1953,1954
<EOL>|1955,1956
Patient|1956,1963
previously|1964,1974
did|1975,1978
not|1979,1982
tolerate|1983,1991
this|1992,1996
medication|1997,2007
while|2008,2013
on|2014,2016
<EOL>|2017,2018
pembrolizumab|2018,2031
(|2032,2033
dizziness|2033,2042
and|2043,2046
_|2047,2048
_|2048,2049
_|2049,2050
,|2050,2051
but|2052,2055
patient|2056,2063
has|2064,2067
been|2068,2072
off|2073,2076
of|2077,2079
<EOL>|2080,2081
pembrolizumab|2081,2094
since|2095,2100
_|2101,2102
_|2102,2103
_|2103,2104
<EOL>|2104,2105
[|2105,2106
]|2106,2107
Consider|2108,2116
starting|2117,2125
spironolactone|2126,2140
and|2141,2144
_|2145,2146
_|2146,2147
_|2147,2148
pending|2149,2156
blood|2157,2162
<EOL>|2163,2164
pressures|2164,2173
;|2173,2174
trialed|2175,2182
losartan|2183,2191
and|2192,2195
spironolactone|2196,2210
during|2211,2217
this|2218,2222
<EOL>|2223,2224
admission|2224,2233
,|2233,2234
but|2235,2238
ultimately|2239,2249
held|2250,2254
due|2255,2258
to|2259,2261
hypotension|2262,2273
.|2273,2274
<EOL>|2275,2276
[|2276,2277
]|2277,2278
His|2279,2282
LFTs|2283,2287
should|2288,2294
be|2295,2297
rechecked|2298,2307
~|2308,2309
2|2309,2310
weeks|2311,2316
after|2317,2322
discharge|2323,2332
<EOL>|2333,2334
(|2334,2335
_|2335,2336
_|2336,2337
_|2337,2338
)|2338,2339
.|2339,2340
He|2341,2343
has|2344,2347
a|2348,2349
history|2350,2357
of|2358,2360
transaminitis|2361,2374
attributed|2375,2385
in|2386,2388
part|2389,2393
<EOL>|2394,2395
to|2395,2397
statin|2398,2404
use|2405,2408
in|2409,2411
the|2412,2415
past|2416,2420
;|2420,2421
he|2422,2424
was|2425,2428
restarted|2429,2438
on|2439,2441
rosuvastatin|2442,2454
this|2455,2459
<EOL>|2460,2461
admission|2461,2470
(|2471,2472
given|2472,2477
history|2478,2485
of|2486,2488
CAD|2489,2492
s|2493,2494
/|2494,2495
p|2495,2496
CABG|2497,2501
)|2501,2502
,|2502,2503
and|2504,2507
LFTs|2508,2512
on|2513,2515
day|2516,2519
of|2520,2522
<EOL>|2523,2524
admission|2524,2533
were|2534,2538
ALT|2539,2542
38|2543,2545
,|2545,2546
AST|2547,2550
46|2551,2553
,|2553,2554
Alk|2555,2558
phos|2559,2563
108|2564,2567
,|2567,2568
Tbili|2569,2574
0.5|2575,2578
.|2578,2579
<EOL>|2579,2580
[|2580,2581
]|2581,2582
Follow|2583,2589
up|2590,2592
with|2593,2597
Oncology|2598,2606
regarding|2607,2616
melanoma|2617,2625
.|2625,2626
<EOL>|2626,2627
[|2627,2628
]|2628,2629
Monitor|2630,2637
for|2638,2641
resolution|2642,2652
of|2653,2655
supplemental|2656,2668
O2|2669,2671
requirement|2672,2683
after|2684,2689
<EOL>|2690,2691
discharge|2691,2700
.|2700,2701
He|2702,2704
was|2705,2708
requiring|2709,2718
_|2719,2720
_|2720,2721
_|2721,2722
of|2723,2725
O2|2726,2728
by|2729,2731
NC|2732,2734
at|2735,2737
time|2738,2742
of|2743,2745
<EOL>|2746,2747
discharge|2747,2756
,|2756,2757
in|2758,2760
the|2761,2764
setting|2765,2772
of|2773,2775
recovering|2776,2786
from|2787,2791
pneumonia|2792,2801
.|2801,2802
<EOL>|2802,2803
<EOL>|2803,2804
DISCHARGE|2804,2813
WT|2814,2816
:|2816,2817
116.18|2818,2824
lbs|2825,2828
<EOL>|2828,2829
DISCHARTE|2829,2838
Cr|2839,2841
:|2841,2842
2.0|2843,2846
<EOL>|2846,2847
DISCHARGE|2847,2856
DIURETIC|2857,2865
:|2865,2866
torsemide|2867,2876
60|2877,2879
mg|2880,2882
PO|2883,2885
BID|2886,2889
<EOL>|2889,2890
<EOL>|2890,2891
SUMMARY|2891,2898
:|2898,2899
<EOL>|2899,2900
=|2900,2901
=|2901,2902
=|2902,2903
=|2903,2904
=|2904,2905
=|2905,2906
=|2906,2907
=|2907,2908
=|2908,2909
=|2909,2910
=|2910,2911
=|2911,2912
=|2912,2913
=|2913,2914
=|2914,2915
<EOL>|2915,2916
Mr.|2916,2919
_|2920,2921
_|2921,2922
_|2922,2923
is|2924,2926
a|2927,2928
_|2929,2930
_|2930,2931
_|2931,2932
man|2933,2936
with|2937,2941
PMH|2942,2945
of|2946,2948
HFrEF|2949,2954
(|2955,2956
35|2956,2958
%|2958,2959
<EOL>|2960,2961
_|2961,2962
_|2962,2963
_|2963,2964
,|2964,2965
<EOL>|2965,2966
CAD|2966,2969
s|2970,2971
/|2971,2972
p|2972,2973
3v|2974,2976
CABG|2977,2981
(|2982,2983
_|2983,2984
_|2984,2985
_|2985,2986
)|2986,2987
and|2988,2991
subsequent|2992,3002
PCI|3003,3006
to|3007,3009
the|3010,3013
LAD|3014,3017
(|3018,3019
_|3019,3020
_|3020,3021
_|3021,3022
)|3022,3023
,|3023,3024
<EOL>|3024,3025
moderate|3025,3033
tricuspid|3034,3043
regurgitation|3044,3057
,|3057,3058
right|3059,3064
ventricular|3065,3076
dysfunction|3077,3088
,|3088,3089
<EOL>|3089,3090
moderate|3090,3098
pulmonary|3099,3108
hypertension|3109,3121
,|3121,3122
and|3123,3126
paroxysmal|3127,3137
atrial|3138,3144
<EOL>|3145,3146
fibrillation|3146,3158
on|3159,3161
apixaban|3162,3170
,|3170,3171
stage|3172,3177
III|3178,3181
chronic|3182,3189
kidney|3190,3196
disease|3197,3204
<EOL>|3205,3206
(|3206,3207
Baseline|3207,3215
Cr|3216,3218
2.0|3219,3222
-|3222,3223
2.1|3223,3226
)|3226,3227
,|3227,3228
cerebrovascular|3229,3244
disease|3245,3252
,|3252,3253
and|3254,3257
metastatic|3258,3268
<EOL>|3269,3270
melanoma|3270,3278
of|3279,3281
unknown|3282,3289
primary|3290,3297
on|3298,3300
Pembrolizumab|3301,3314
(|3315,3316
on|3316,3318
hold|3319,3323
since|3324,3329
<EOL>|3330,3331
_|3331,3332
_|3332,3333
_|3333,3334
iso|3335,3338
worsening|3339,3348
transaminitis|3349,3362
and|3363,3366
concern|3367,3374
for|3375,3378
<EOL>|3379,3380
cardiotoxicity|3380,3394
)|3394,3395
.|3395,3396
He|3397,3399
was|3400,3403
admitted|3404,3412
with|3413,3417
volume|3418,3424
overload|3425,3433
from|3434,3438
heart|3439,3444
<EOL>|3445,3446
failure|3446,3453
exacerbation|3454,3466
and|3467,3470
pneumonia|3471,3480
with|3481,3485
high|3486,3490
oxygen|3491,3497
<EOL>|3498,3499
requirements|3499,3511
.|3511,3512
He|3513,3515
initially|3516,3525
required|3526,3534
CCU|3535,3538
admission|3539,3548
for|3549,3552
high|3553,3557
flow|3558,3562
<EOL>|3563,3564
oxygen|3564,3570
,|3570,3571
weaned|3572,3578
to|3579,3581
nasal|3582,3587
cannula|3588,3595
after|3596,3601
aggressive|3602,3612
IV|3613,3615
diuresis|3616,3624
and|3625,3628
<EOL>|3629,3630
treatment|3630,3639
of|3640,3642
pneumonia|3643,3652
with|3653,3657
5|3658,3659
day|3660,3663
course|3664,3670
of|3671,3673
Zosyn|3674,3679
after|3680,3685
<EOL>|3686,3687
receiving|3687,3696
vancomycin|3697,3707
at|3708,3710
OSH|3711,3714
.|3714,3715
He|3716,3718
was|3719,3722
transferred|3723,3734
to|3735,3737
cardiology|3738,3748
<EOL>|3749,3750
floor|3750,3755
where|3756,3761
he|3762,3764
continued|3765,3774
to|3775,3777
diurese|3778,3785
well|3786,3790
and|3791,3794
his|3795,3798
oxygen|3799,3805
<EOL>|3806,3807
requirement|3807,3818
was|3819,3822
weaned|3823,3829
to|3830,3832
_|3833,3834
_|3834,3835
_|3835,3836
.|3836,3837
He|3838,3840
was|3841,3844
transitioned|3845,3857
to|3858,3860
60|3861,3863
mg|3864,3866
<EOL>|3867,3868
torsemide|3868,3877
PO|3878,3880
BID|3881,3884
which|3885,3890
adequately|3891,3901
maintained|3902,3912
euvolemia|3913,3922
.|3922,3923
<EOL>|3924,3925
<EOL>|3925,3926
ACUTE|3926,3931
ISSUES|3932,3938
:|3938,3939
<EOL>|3940,3941
=|3941,3942
=|3942,3943
=|3943,3944
=|3944,3945
=|3945,3946
=|3946,3947
=|3947,3948
=|3948,3949
=|3949,3950
=|3950,3951
=|3951,3952
=|3952,3953
=|3953,3954
<EOL>|3955,3956
#|3956,3957
Acute|3958,3963
on|3964,3966
chronic|3967,3974
systolic|3975,3983
heart|3984,3989
failure|3990,3997
exacerbation|3998,4010
<EOL>|4010,4011
Patient|4011,4018
with|4019,4023
history|4024,4031
of|4032,4034
heart|4035,4040
failure|4041,4048
with|4049,4053
etiology|4054,4062
likely|4063,4069
<EOL>|4070,4071
ischemic|4071,4079
cardiomyopathy|4080,4094
given|4095,4100
history|4101,4108
of|4109,4111
CAD|4112,4115
s|4116,4117
/|4117,4118
p|4118,4119
CABG|4120,4124
and|4125,4128
PCI|4129,4132
.|4132,4133
<EOL>|4134,4135
Admitted|4135,4143
with|4144,4148
fluid|4149,4154
overload|4155,4163
and|4164,4167
pleural|4168,4175
effusion|4176,4184
.|4184,4185
Trigger|4186,4193
for|4194,4197
<EOL>|4198,4199
current|4199,4206
exacerbation|4207,4219
could|4220,4225
be|4226,4228
infectious|4229,4239
given|4240,4245
evidence|4246,4254
of|4255,4257
<EOL>|4258,4259
pneumonia|4259,4268
in|4269,4271
left|4272,4276
lower|4277,4282
lobe|4283,4287
on|4288,4290
admission|4291,4300
.|4300,4301
Patient|4302,4309
with|4310,4314
high|4315,4319
<EOL>|4320,4321
oxygen|4321,4327
requirements|4328,4340
prior|4341,4346
to|4347,4349
admission|4350,4359
but|4360,4363
responded|4364,4373
<EOL>|4374,4375
appropriately|4375,4388
to|4389,4391
diuresis|4392,4400
with|4401,4405
Lasix|4406,4411
.|4411,4412
After|4413,4418
IV|4419,4421
diuresis|4422,4430
,|4430,4431
patient|4432,4439
<EOL>|4440,4441
was|4441,4444
transitioned|4445,4457
PO|4458,4460
torsemide|4461,4470
and|4471,4474
maintained|4475,4485
at|4486,4488
euvolemia|4489,4498
.|4498,4499
With|4500,4504
<EOL>|4505,4506
effective|4506,4515
diuresis|4516,4524
,|4524,4525
the|4526,4529
patient|4530,4537
's|4537,4539
oxygen|4540,4546
requirement|4547,4558
gradually|4559,4568
<EOL>|4569,4570
lowered|4570,4577
from|4578,4582
4L|4583,4585
NC|4586,4588
to|4589,4591
_|4592,4593
_|4593,4594
_|4594,4595
NC|4596,4598
.|4598,4599
He|4600,4602
was|4603,4606
discharged|4607,4617
on|4618,4620
torsemide|4621,4630
60|4631,4633
<EOL>|4634,4635
mg|4635,4637
PO|4638,4640
BID|4641,4644
.|4644,4645
He|4646,4648
was|4649,4652
unable|4653,4659
to|4660,4662
tolerate|4663,4671
afterload|4672,4681
reducing|4682,4690
agents|4691,4697
<EOL>|4698,4699
or|4699,4701
neurohormonal|4702,4715
blockade|4716,4724
agents|4725,4731
due|4732,4735
to|4736,4738
hypotension|4739,4750
.|4750,4751
<EOL>|4752,4753
<EOL>|4753,4754
#|4754,4755
Lower|4756,4761
left|4762,4766
lobe|4767,4771
pneumonia|4772,4781
<EOL>|4781,4782
Patient|4782,4789
with|4790,4794
evidence|4795,4803
of|4804,4806
pneumonia|4807,4816
in|4817,4819
the|4820,4823
left|4824,4828
lower|4829,4834
lobe|4835,4839
,|4839,4840
<EOL>|4841,4842
received|4842,4850
vanc|4851,4855
/|4855,4856
zosyn|4856,4861
at|4862,4864
outside|4865,4872
hospital|4873,4881
and|4882,4885
continued|4886,4895
on|4896,4898
Zosyn|4899,4904
<EOL>|4905,4906
here|4906,4910
for|4911,4914
a|4915,4916
total|4917,4922
of|4923,4925
5|4926,4927
day|4928,4931
course|4932,4938
with|4939,4943
resolution|4944,4954
of|4955,4957
symptoms|4958,4966
.|4966,4967
We|4968,4970
<EOL>|4971,4972
suspect|4972,4979
that|4980,4984
his|4985,4988
lingering|4989,4998
O2|4999,5001
requirement|5002,5013
is|5014,5016
at|5017,5019
least|5020,5025
in|5026,5028
part|5029,5033
<EOL>|5034,5035
due|5035,5038
to|5039,5041
slowly|5042,5048
resorbing|5049,5058
consolidation|5059,5072
left|5073,5077
over|5078,5082
from|5083,5087
his|5088,5091
<EOL>|5092,5093
infection|5093,5102
.|5102,5103
He|5104,5106
was|5107,5110
requiring|5111,5120
_|5121,5122
_|5122,5123
_|5123,5124
of|5125,5127
supplemental|5128,5140
O2|5141,5143
by|5144,5146
NC|5147,5149
at|5150,5152
<EOL>|5153,5154
time|5154,5158
of|5159,5161
discharge|5162,5171
.|5171,5172
<EOL>|5172,5173
<EOL>|5173,5174
#|5174,5175
Pleural|5176,5183
effusion|5184,5192
,|5192,5193
bilateral|5194,5203
<EOL>|5203,5204
Patient|5204,5211
with|5212,5216
evidence|5217,5225
of|5226,5228
right|5229,5234
pleural|5235,5242
effusion|5243,5251
.|5251,5252
Etiology|5253,5261
likely|5262,5268
<EOL>|5269,5270
fluid|5270,5275
overload|5276,5284
given|5285,5290
heart|5291,5296
failure|5297,5304
with|5305,5309
reduced|5310,5317
ejection|5318,5326
<EOL>|5327,5328
fraction|5328,5336
.|5336,5337
Pleural|5338,5345
effusion|5346,5354
resolved|5355,5363
improved|5364,5372
with|5373,5377
diuresis|5378,5386
and|5387,5390
<EOL>|5391,5392
his|5392,5395
oxygen|5396,5402
requirement|5403,5414
trended|5415,5422
down|5423,5427
to|5428,5430
_|5431,5432
_|5432,5433
_|5433,5434
NC|5435,5437
.|5437,5438
Given|5439,5444
this|5445,5449
,|5449,5450
<EOL>|5451,5452
thoracentesis|5452,5465
was|5466,5469
deferred|5470,5478
.|5478,5479
<EOL>|5480,5481
<EOL>|5481,5482
#|5482,5483
Atrial|5484,5490
fibrillation|5491,5503
<EOL>|5503,5504
Patient|5504,5511
with|5512,5516
chronic|5517,5524
history|5525,5532
of|5533,5535
atrial|5536,5542
fibrillation|5543,5555
.|5555,5556
In|5557,5559
afib|5560,5564
<EOL>|5565,5566
throughout|5566,5576
this|5577,5581
admission|5582,5591
.|5591,5592
Continued|5593,5602
amiodarone|5603,5613
and|5614,5617
apixaban|5618,5626
.|5626,5627
<EOL>|5628,5629
Rates|5629,5634
appropriately|5635,5648
controlled|5649,5659
.|5659,5660
<EOL>|5660,5661
<EOL>|5661,5662
CHRONIC|5662,5669
ISSUES|5670,5676
<EOL>|5676,5677
=|5677,5678
=|5678,5679
=|5679,5680
=|5680,5681
=|5681,5682
=|5682,5683
=|5683,5684
=|5684,5685
=|5685,5686
=|5686,5687
=|5687,5688
=|5688,5689
=|5689,5690
=|5690,5691
=|5691,5692
=|5692,5693
<EOL>|5693,5694
#|5694,5695
Coronary|5696,5704
artery|5705,5711
disease|5712,5719
s|5720,5721
/|5721,5722
p|5722,5723
CABG|5724,5728
<EOL>|5728,5729
Patient|5729,5736
with|5737,5741
history|5742,5749
of|5750,5752
3|5753,5754
vessel|5755,5761
CABG|5762,5766
on|5767,5769
_|5770,5771
_|5771,5772
_|5772,5773
(|5774,5775
_|5775,5776
_|5776,5777
_|5777,5778
)|5778,5779
and|5780,5783
<EOL>|5783,5784
subsequent|5784,5794
PCI|5795,5798
to|5799,5801
LAD|5802,5805
(|5806,5807
_|5807,5808
_|5808,5809
_|5809,5810
)|5810,5811
.|5811,5812
Continued|5813,5822
home|5823,5827
aspirin|5828,5835
.|5835,5836
Patient|5837,5844
<EOL>|5845,5846
was|5846,5849
started|5850,5857
on|5858,5860
low|5861,5864
dose|5865,5869
rosuvastatin|5870,5882
5|5883,5884
mg|5885,5887
daily|5888,5893
.|5893,5894
On|5895,5897
review|5898,5904
,|5904,5905
it|5906,5908
<EOL>|5909,5910
appears|5910,5917
he|5918,5920
had|5921,5924
been|5925,5929
on|5930,5932
this|5933,5937
medication|5938,5948
at|5949,5951
this|5952,5956
dose|5957,5961
in|5962,5964
the|5965,5968
past|5969,5973
<EOL>|5974,5975
but|5975,5978
it|5979,5981
was|5982,5985
discontinued|5986,5998
due|5999,6002
to|6003,6005
transamnitis|6006,6018
;|6018,6019
however|6020,6027
,|6027,6028
at|6029,6031
the|6032,6035
<EOL>|6036,6037
time|6037,6041
it|6042,6044
was|6045,6048
unclear|6049,6056
whether|6057,6064
this|6065,6069
was|6070,6073
an|6074,6076
effect|6077,6083
of|6084,6086
the|6087,6090
statin|6091,6097
or|6098,6100
<EOL>|6101,6102
pembrolizumab|6102,6115
.|6115,6116
Given|6117,6122
that|6123,6127
the|6128,6131
patient|6132,6139
has|6140,6143
not|6144,6147
had|6148,6151
his|6152,6155
checkpoint|6156,6166
<EOL>|6167,6168
inhibitor|6168,6177
therapy|6178,6185
since|6186,6191
_|6192,6193
_|6193,6194
_|6194,6195
,|6195,6196
the|6197,6200
decision|6201,6209
was|6210,6213
to|6214,6216
restart|6217,6224
<EOL>|6225,6226
rosuvastatin|6226,6238
.|6238,6239
<EOL>|6240,6241
<EOL>|6241,6242
#|6242,6243
Chronic|6244,6251
kidney|6252,6258
disease|6259,6266
<EOL>|6266,6267
Baseline|6267,6275
Cr|6276,6278
appears|6279,6286
to|6287,6289
be|6290,6292
2.1|6293,6296
-|6296,6297
2.2|6297,6300
over|6301,6305
past|6306,6310
year|6311,6315
.|6315,6316
Cr|6317,6319
remained|6320,6328
<EOL>|6329,6330
between|6330,6337
1.8|6338,6341
-|6341,6342
2.4|6342,6345
throughout|6346,6356
admission|6357,6366
.|6366,6367
<EOL>|6368,6369
<EOL>|6369,6370
#|6370,6371
Anemia|6372,6378
<EOL>|6378,6379
Chronic|6379,6386
,|6386,6387
although|6388,6396
worsening|6397,6406
since|6407,6412
_|6413,6414
_|6414,6415
_|6415,6416
.|6416,6417
On|6418,6420
admission|6421,6430
<EOL>|6431,6432
hemoglobin|6432,6442
<EOL>|6442,6443
10.6|6443,6447
and|6448,6451
remained|6452,6460
stable|6461,6467
.|6467,6468
<EOL>|6469,6470
<EOL>|6470,6471
#|6471,6472
Thrombocytopenia|6473,6489
<EOL>|6489,6490
Uncertain|6490,6499
etiology|6500,6508
,|6508,6509
appears|6510,6517
subacute|6518,6526
/|6526,6527
chronic|6527,6534
.|6534,6535
On|6536,6538
admission|6539,6548
<EOL>|6548,6549
platelets|6549,6558
130|6559,6562
down|6563,6567
-|6567,6568
trended|6568,6575
to|6576,6578
100s|6579,6583
.|6583,6584
No|6585,6587
concern|6588,6595
for|6596,6599
bleeding|6600,6608
<EOL>|6609,6610
throughout|6610,6620
admission|6621,6630
.|6630,6631
<EOL>|6632,6633
<EOL>|6633,6634
#|6634,6635
Melanoma|6636,6644
<EOL>|6644,6645
Patient|6645,6652
with|6653,6657
history|6658,6665
of|6666,6668
metastatic|6669,6679
melanoma|6680,6688
with|6689,6693
unknown|6694,6701
<EOL>|6702,6703
primary|6703,6710
.|6710,6711
<EOL>|6711,6712
On|6712,6714
treatment|6715,6724
with|6725,6729
pembrolizumab|6730,6743
,|6743,6744
but|6745,6748
held|6749,6753
since|6754,6759
_|6760,6761
_|6761,6762
_|6762,6763
iso|6764,6767
<EOL>|6767,6768
toxicity|6768,6776
.|6776,6777
<EOL>|6778,6779
<EOL>|6779,6780
CODE|6780,6784
:|6784,6785
DNR|6786,6789
/|6789,6790
DNI|6790,6793
<EOL>|6793,6794
CONTACT|6794,6801
:|6801,6802
_|6803,6804
_|6804,6805
_|6805,6806
(|6807,6808
_|6808,6809
_|6809,6810
_|6810,6811
)|6811,6812
<EOL>|6812,6813
Relationship|6813,6825
:|6825,6826
Son|6827,6830
<EOL>|6831,6832
Phone|6832,6837
number|6838,6844
:|6844,6845
_|6846,6847
_|6847,6848
_|6848,6849
<EOL>|6849,6850
<EOL>|6851,6852
_|6852,6853
_|6853,6854
_|6854,6855
on|6856,6858
Admission|6859,6868
:|6868,6869
<EOL>|6869,6870
The|6870,6873
Preadmission|6874,6886
Medication|6887,6897
list|6898,6902
is|6903,6905
accurate|6906,6914
and|6915,6918
complete|6919,6927
.|6927,6928
<EOL>|6928,6929
1.|6929,6931
Amiodarone|6932,6942
200|6943,6946
mg|6947,6949
PO|6950,6952
DAILY|6953,6958
<EOL>|6959,6960
2.|6960,6962
Apixaban|6963,6971
2.5|6972,6975
mg|6976,6978
PO|6979,6981
BID|6982,6985
<EOL>|6986,6987
3.|6987,6989
Aspirin|6990,6997
81|6998,7000
mg|7001,7003
PO|7004,7006
DAILY|7007,7012
<EOL>|7013,7014
4.|7014,7016
Docusate|7017,7025
Sodium|7026,7032
100|7033,7036
mg|7037,7039
PO|7040,7042
BID|7043,7046
<EOL>|7047,7048
5.|7048,7050
Ferrous|7051,7058
Sulfate|7059,7066
325|7067,7070
mg|7071,7073
PO|7074,7076
DAILY|7077,7082
<EOL>|7083,7084
6.|7084,7086
Senna|7087,7092
17.2|7093,7097
mg|7098,7100
PO|7101,7103
HS|7104,7106
<EOL>|7107,7108
7.|7108,7110
Sertraline|7111,7121
50|7122,7124
mg|7125,7127
PO|7128,7130
DAILY|7131,7136
<EOL>|7137,7138
8.|7138,7140
Tamsulosin|7141,7151
0.4|7152,7155
mg|7156,7158
PO|7159,7161
QHS|7162,7165
<EOL>|7166,7167
9.|7167,7169
Torsemide|7170,7179
40|7180,7182
mg|7183,7185
PO|7186,7188
DAILY|7189,7194
<EOL>|7195,7196
10.|7196,7199
coenzyme|7200,7208
Q10|7209,7212
100|7213,7216
mg|7217,7219
oral|7220,7224
DAILY|7225,7230
<EOL>|7231,7232
11.|7232,7235
Align|7236,7241
(|7242,7243
bifidobacterium|7243,7258
infantis|7259,7267
)|7267,7268
4|7269,7270
mg|7271,7273
oral|7274,7278
DAILY|7279,7284
<EOL>|7285,7286
12.|7286,7289
Potassium|7290,7299
Chloride|7300,7308
40|7309,7311
mEq|7312,7315
PO|7316,7318
DAILY|7319,7324
<EOL>|7325,7326
<EOL>|7326,7327
<EOL>|7328,7329
Discharge|7329,7338
Medications|7339,7350
:|7350,7351
<EOL>|7351,7352
1.|7352,7354
Rosuvastatin|7356,7368
Calcium|7369,7376
5|7377,7378
mg|7379,7381
PO|7382,7384
QPM|7385,7388
<EOL>|7390,7391
2.|7391,7393
Vitamin|7395,7402
D|7403,7404
1000|7405,7409
UNIT|7410,7414
PO|7415,7417
DAILY|7418,7423
<EOL>|7425,7426
3.|7426,7428
Torsemide|7430,7439
60|7440,7442
mg|7443,7445
PO|7446,7448
BID|7449,7452
<EOL>|7454,7455
4.|7455,7457
Align|7459,7464
(|7465,7466
bifidobacterium|7466,7481
infantis|7482,7490
)|7490,7491
4|7492,7493
mg|7494,7496
oral|7497,7501
DAILY|7502,7507
<EOL>|7509,7510
5.|7510,7512
Amiodarone|7514,7524
200|7525,7528
mg|7529,7531
PO|7532,7534
DAILY|7535,7540
<EOL>|7542,7543
6.|7543,7545
Apixaban|7547,7555
2.5|7556,7559
mg|7560,7562
PO|7563,7565
BID|7566,7569
<EOL>|7571,7572
7.|7572,7574
Aspirin|7576,7583
81|7584,7586
mg|7587,7589
PO|7590,7592
DAILY|7593,7598
<EOL>|7600,7601
8.|7601,7603
coenzyme|7605,7613
Q10|7614,7617
100|7618,7621
mg|7622,7624
oral|7625,7629
DAILY|7630,7635
<EOL>|7637,7638
9.|7638,7640
Docusate|7642,7650
Sodium|7651,7657
100|7658,7661
mg|7662,7664
PO|7665,7667
BID|7668,7671
<EOL>|7673,7674
10.|7674,7677
Ferrous|7679,7686
Sulfate|7687,7694
325|7695,7698
mg|7699,7701
PO|7702,7704
DAILY|7705,7710
<EOL>|7712,7713
11.|7713,7716
Potassium|7718,7727
Chloride|7728,7736
40|7737,7739
mEq|7740,7743
PO|7744,7746
DAILY|7747,7752
<EOL>|7754,7755
12.|7755,7758
Senna|7760,7765
17.2|7766,7770
mg|7771,7773
PO|7774,7776
HS|7777,7779
<EOL>|7781,7782
13.|7782,7785
Sertraline|7787,7797
50|7798,7800
mg|7801,7803
PO|7804,7806
DAILY|7807,7812
<EOL>|7814,7815
14.|7815,7818
Tamsulosin|7820,7830
0.4|7831,7834
mg|7835,7837
PO|7838,7840
QHS|7841,7844
<EOL>|7846,7847
<EOL>|7847,7848
_|7848,7849
_|7849,7850
_|7850,7851
and|7852,7855
mineralocorticoid|7856,7873
receptor|7874,7882
antagonist|7883,7893
held|7894,7898
in|7899,7901
the|7902,7905
<EOL>|7906,7907
setting|7907,7914
of|7915,7917
hypotension|7918,7929
and|7930,7933
CKD|7934,7937
.|7937,7938
Patient|7939,7946
is|7947,7949
intolerant|7950,7960
of|7961,7963
beta|7964,7968
<EOL>|7969,7970
blockers|7970,7978
due|7979,7982
to|7983,7985
dizziness|7986,7995
/|7995,7996
hypotension|7996,8007
previously|8008,8018
.|8018,8019
<EOL>|8019,8020
<EOL>|8021,8022
Discharge|8022,8031
Disposition|8032,8043
:|8043,8044
<EOL>|8044,8045
Extended|8045,8053
Care|8054,8058
<EOL>|8058,8059
<EOL>|8060,8061
Facility|8061,8069
:|8069,8070
<EOL>|8070,8071
_|8071,8072
_|8072,8073
_|8073,8074
<EOL>|8074,8075
<EOL>|8076,8077
Discharge|8077,8086
Diagnosis|8087,8096
:|8096,8097
<EOL>|8097,8098
Primary|8098,8105
diagnosis|8106,8115
:|8115,8116
<EOL>|8116,8117
=|8117,8118
=|8118,8119
=|8119,8120
=|8120,8121
=|8121,8122
=|8122,8123
=|8123,8124
=|8124,8125
=|8125,8126
=|8126,8127
=|8127,8128
=|8128,8129
=|8129,8130
=|8130,8131
=|8131,8132
=|8132,8133
=|8133,8134
=|8134,8135
=|8135,8136
=|8136,8137
=|8137,8138
<EOL>|8138,8139
Acute|8139,8144
on|8145,8147
chronic|8148,8155
systolic|8156,8164
heart|8165,8170
failure|8171,8178
exacerbation|8179,8191
<EOL>|8191,8192
Lower|8192,8197
left|8198,8202
lobe|8203,8207
pneumonia|8208,8217
<EOL>|8217,8218
Bilateral|8218,8227
pleural|8228,8235
effusion|8236,8244
<EOL>|8244,8245
Atrial|8245,8251
fibrillation|8252,8264
<EOL>|8264,8265
<EOL>|8265,8266
Secondary|8266,8275
diagnosis|8276,8285
:|8285,8286
<EOL>|8286,8287
=|8287,8288
=|8288,8289
=|8289,8290
=|8290,8291
=|8291,8292
=|8292,8293
=|8293,8294
=|8294,8295
=|8295,8296
=|8296,8297
=|8297,8298
=|8298,8299
=|8299,8300
=|8300,8301
=|8301,8302
=|8302,8303
=|8303,8304
=|8304,8305
=|8305,8306
=|8306,8307
=|8307,8308
<EOL>|8308,8309
Coronary|8309,8317
artery|8318,8324
disease|8325,8332
status|8333,8339
post|8340,8344
CABG|8345,8349
<EOL>|8349,8350
Chronic|8350,8357
kidney|8358,8364
disease|8365,8372
<EOL>|8372,8373
Anemia|8373,8379
<EOL>|8379,8380
Thrombocytopenia|8380,8396
<EOL>|8396,8397
Metastatic|8397,8407
melanoma|8408,8416
<EOL>|8416,8417
<EOL>|8417,8418
<EOL>|8419,8420
Discharge|8420,8429
Condition|8430,8439
:|8439,8440
<EOL>|8440,8441
Mental|8441,8447
Status|8448,8454
:|8454,8455
Clear|8456,8461
and|8462,8465
coherent|8466,8474
.|8474,8475
<EOL>|8475,8476
Level|8476,8481
of|8482,8484
Consciousness|8485,8498
:|8498,8499
Alert|8500,8505
and|8506,8509
interactive|8510,8521
.|8521,8522
<EOL>|8522,8523
Activity|8523,8531
Status|8532,8538
:|8538,8539
Ambulatory|8540,8550
-|8551,8552
requires|8553,8561
assistance|8562,8572
or|8573,8575
aid|8576,8579
(|8580,8581
walker|8581,8587
<EOL>|8588,8589
or|8589,8591
cane|8592,8596
)|8596,8597
.|8597,8598
<EOL>|8598,8599
<EOL>|8599,8600
<EOL>|8601,8602
Discharge|8602,8611
Instructions|8612,8624
:|8624,8625
<EOL>|8625,8626
Dear|8626,8630
Mr.|8631,8634
_|8635,8636
_|8636,8637
_|8637,8638
,|8638,8639
<EOL>|8639,8640
<EOL>|8640,8641
It|8641,8643
was|8644,8647
a|8648,8649
pleasure|8650,8658
taking|8659,8665
care|8666,8670
of|8671,8673
you|8674,8677
at|8678,8680
the|8681,8684
_|8685,8686
_|8686,8687
_|8687,8688
<EOL>|8689,8690
_|8690,8691
_|8691,8692
_|8692,8693
.|8693,8694
<EOL>|8695,8696
<EOL>|8696,8697
WHY|8697,8700
WAS|8701,8704
I|8705,8706
IN|8707,8709
THE|8710,8713
HOSPITAL|8714,8722
?|8722,8723
<EOL>|8725,8726
=|8726,8727
=|8727,8728
=|8728,8729
=|8729,8730
=|8730,8731
=|8731,8732
=|8732,8733
=|8733,8734
=|8734,8735
=|8735,8736
=|8736,8737
=|8737,8738
=|8738,8739
=|8739,8740
=|8740,8741
=|8741,8742
=|8742,8743
=|8743,8744
=|8744,8745
=|8745,8746
=|8746,8747
=|8747,8748
=|8748,8749
=|8749,8750
=|8750,8751
=|8751,8752
<EOL>|8755,8756
-|8756,8757
You|8758,8761
were|8762,8766
admitted|8767,8775
because|8776,8783
of|8784,8786
you|8787,8790
were|8791,8795
short|8796,8801
of|8802,8804
breath|8805,8811
<EOL>|8812,8813
<EOL>|8813,8814
WHAT|8814,8818
HAPPENED|8819,8827
IN|8828,8830
THE|8831,8834
HOSPITAL|8835,8843
?|8843,8844
<EOL>|8846,8847
=|8847,8848
=|8848,8849
=|8849,8850
=|8850,8851
=|8851,8852
=|8852,8853
=|8853,8854
=|8854,8855
=|8855,8856
=|8856,8857
=|8857,8858
=|8858,8859
=|8859,8860
=|8860,8861
=|8861,8862
=|8862,8863
=|8863,8864
=|8864,8865
=|8865,8866
=|8866,8867
=|8867,8868
=|8868,8869
=|8869,8870
=|8870,8871
=|8871,8872
=|8872,8873
=|8873,8874
=|8874,8875
=|8875,8876
=|8876,8877
<EOL>|8879,8880
-|8880,8881
You|8882,8885
were|8886,8890
found|8891,8896
to|8897,8899
have|8900,8904
fluid|8905,8910
on|8911,8913
your|8914,8918
lungs|8919,8924
.|8924,8925
This|8926,8930
was|8931,8934
because|8935,8942
<EOL>|8943,8944
you|8944,8947
have|8948,8952
a|8953,8954
medical|8955,8962
condition|8963,8972
called|8973,8979
heart|8980,8985
failure|8986,8993
,|8993,8994
where|8995,9000
your|9001,9005
<EOL>|9006,9007
heart|9007,9012
does|9013,9017
not|9018,9021
pump|9022,9026
hard|9027,9031
enough|9032,9038
and|9039,9042
fluid|9043,9048
backs|9049,9054
up|9055,9057
into|9058,9062
your|9063,9067
<EOL>|9068,9069
lungs|9069,9074
.|9074,9075
<EOL>|9076,9077
-|9077,9078
You|9079,9082
were|9083,9087
given|9088,9093
a|9094,9095
diuretic|9096,9104
medication|9105,9115
to|9116,9118
help|9119,9123
get|9124,9127
the|9128,9131
fluid|9132,9137
<EOL>|9138,9139
out|9139,9142
.|9142,9143
You|9144,9147
improved|9148,9156
considerably|9157,9169
and|9170,9173
are|9174,9177
ready|9178,9183
to|9184,9186
leave|9187,9192
the|9193,9196
<EOL>|9197,9198
hospital|9198,9206
.|9206,9207
<EOL>|9209,9210
<EOL>|9210,9211
WHAT|9211,9215
SHOULD|9216,9222
I|9223,9224
DO|9225,9227
WHEN|9228,9232
I|9233,9234
GO|9235,9237
HOME|9238,9242
?|9242,9243
<EOL>|9245,9246
=|9246,9247
=|9247,9248
=|9248,9249
=|9249,9250
=|9250,9251
=|9251,9252
=|9252,9253
=|9253,9254
=|9254,9255
=|9255,9256
=|9256,9257
=|9257,9258
=|9258,9259
=|9259,9260
=|9260,9261
=|9261,9262
=|9262,9263
=|9263,9264
=|9264,9265
=|9265,9266
=|9266,9267
=|9267,9268
=|9268,9269
=|9269,9270
=|9270,9271
=|9271,9272
=|9272,9273
=|9273,9274
=|9274,9275
=|9275,9276
=|9276,9277
=|9277,9278
<EOL>|9280,9281
-|9281,9282
Be|9283,9285
sure|9286,9290
to|9291,9293
take|9294,9298
all|9299,9302
your|9303,9307
medications|9308,9319
and|9320,9323
attend|9324,9330
all|9331,9334
of|9335,9337
your|9338,9342
<EOL>|9343,9344
appointments|9344,9356
listed|9357,9363
below|9364,9369
.|9369,9370
<EOL>|9371,9372
-|9372,9373
Your|9374,9378
weight|9379,9385
at|9386,9388
discharge|9389,9398
is|9399,9401
116.18|9402,9408
lbs|9409,9412
.|9412,9413
Please|9414,9420
weigh|9421,9426
yourself|9427,9435
<EOL>|9436,9437
today|9437,9442
at|9443,9445
home|9446,9450
and|9451,9454
use|9455,9458
this|9459,9463
as|9464,9466
your|9467,9471
new|9472,9475
baseline|9476,9484
<EOL>|9486,9487
-|9487,9488
Please|9489,9495
weigh|9496,9501
yourself|9502,9510
every|9511,9516
day|9517,9520
in|9521,9523
the|9524,9527
morning|9528,9535
.|9535,9536
Call|9537,9541
your|9542,9546
<EOL>|9547,9548
doctor|9548,9554
or|9555,9557
the|9558,9561
HeartLine|9562,9571
at|9572,9574
_|9575,9576
_|9576,9577
_|9577,9578
if|9579,9581
your|9582,9586
weight|9587,9593
goes|9594,9598
up|9599,9601
<EOL>|9602,9603
by|9603,9605
more|9606,9610
than|9611,9615
3|9616,9617
lbs|9618,9621
or|9622,9624
you|9625,9628
experience|9629,9639
significant|9640,9651
chest|9652,9657
pain|9658,9662
and|9663,9666
<EOL>|9667,9668
shortness|9668,9677
of|9678,9680
breath|9681,9687
.|9687,9688
<EOL>|9690,9691
<EOL>|9691,9692
Thank|9692,9697
you|9698,9701
for|9702,9705
allowing|9706,9714
us|9715,9717
to|9718,9720
be|9721,9723
involved|9724,9732
in|9733,9735
your|9736,9740
care|9741,9745
,|9745,9746
we|9747,9749
wish|9750,9754
<EOL>|9755,9756
you|9756,9759
all|9760,9763
the|9764,9767
best|9768,9772
!|9772,9773
<EOL>|9775,9776
<EOL>|9776,9777
Sincerely|9777,9786
,|9786,9787
<EOL>|9787,9788
Your|9788,9792
_|9793,9794
_|9794,9795
_|9795,9796
Team|9797,9801
<EOL>|9803,9804
<EOL>|9805,9806
Followup|9806,9814
Instructions|9815,9827
:|9827,9828
<EOL>|9828,9829
_|9829,9830
_|9830,9831
_|9831,9832
<EOL>|9832,9833

