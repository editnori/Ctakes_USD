 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|32,36
No|37,39
:|39,40
_|43,44
_|44,45
_|45,46
<EOL>|46,47
<EOL>|48,49
Admission|49,58
Date|59,63
:|63,64
_|66,67
_|67,68
_|68,69
Discharge|83,92
Date|93,97
:|97,98
_|101,102
_|102,103
_|103,104
<EOL>|104,105
<EOL>|106,107
Date|107,111
of|112,114
Birth|115,120
:|120,121
_|123,124
_|124,125
_|125,126
Sex|139,142
:|142,143
F|146,147
<EOL>|147,148
<EOL>|149,150
Service|150,157
:|157,158
MEDICINE|159,167
<EOL>|167,168
<EOL>|169,170
_|182,183
_|183,184
_|184,185
<EOL>|185,186
<EOL>|187,188
Attending|188,197
:|197,198
_|199,200
_|200,201
_|201,202
.|202,203
<EOL>|203,204
<EOL>|205,206
Abdominal|223,232
pain|233,237
<EOL>|238,239
<EOL>|240,241
Major|241,246
Surgical|247,255
or|256,258
Invasive|259,267
Procedure|268,277
:|277,278
<EOL>|278,279
Colonoscopy|279,290
with|291,295
biopsy|296,302
_|303,304
_|304,305
_|305,306
<EOL>|306,307
<EOL>|307,308
<EOL>|309,310
This|338,342
patient|343,350
is|351,353
a|354,355
_|356,357
_|357,358
_|358,359
year|360,364
old|365,368
female|369,375
with|376,380
Hx|381,383
of|384,386
sigmoid|387,394
<EOL>|395,396
diverticulitis|396,410
s|411,412
/|412,413
p|413,414
resection|415,424
in|425,427
_|428,429
_|429,430
_|430,431
,|431,432
who|433,436
complains|437,446
of|447,449
RLQ|450,453
<EOL>|454,455
abdominal|455,464
pain|465,469
.|469,470
The|471,474
patient|475,482
states|483,489
that|490,494
her|495,498
pain|499,503
began|504,509
yesterday|510,519
<EOL>|520,521
afternoon|521,530
,|530,531
worsened|532,540
overnight|541,550
and|551,554
causing|555,562
her|563,566
to|567,569
present|570,577
to|578,580
the|581,584
<EOL>|585,586
ED|586,588
around|589,595
3AM|596,599
.|599,600
She|601,604
describes|605,614
it|615,617
as|618,620
a|621,622
"|623,624
gnawing|624,631
"|631,632
pain|633,637
,|637,638
<EOL>|639,640
nonradiating|640,652
,|652,653
constant|654,662
and|663,666
_|667,668
_|668,669
_|669,670
intensity|671,680
.|680,681
She|682,685
states|686,692
this|693,697
<EOL>|698,699
feels|699,704
similar|705,712
to|713,715
her|716,719
episode|720,727
of|728,730
diverticulitis|731,745
several|746,753
years|754,759
<EOL>|760,761
ago|761,764
,|764,765
only|766,770
is|771,773
present|774,781
on|782,784
the|785,788
other|789,794
side|795,799
of|800,802
her|803,806
abdomen|807,814
.|814,815
She|816,819
<EOL>|820,821
denies|821,827
any|828,831
fever|832,837
,|837,838
nausea|839,845
,|845,846
vomiting|847,855
,|855,856
SOB|857,860
,|860,861
Chest|862,867
pain|868,872
,|872,873
BRBPR|874,879
.|879,880
She|881,884
<EOL>|885,886
does|886,890
endorse|891,898
subjective|899,909
feeling|910,917
of|918,920
chills|921,927
.|927,928
<EOL>|930,931
.|931,932
<EOL>|934,935
Prior|935,940
to|941,943
the|944,947
current|948,955
episode|956,963
,|963,964
the|965,968
patient|969,976
reports|977,984
having|985,991
a|992,993
<EOL>|994,995
"|995,996
sinus|996,1001
infection|1002,1011
"|1011,1012
about|1013,1018
3|1019,1020
weeks|1021,1026
ago|1027,1030
that|1031,1035
resolved|1036,1044
over|1045,1049
one|1050,1053
week|1054,1058
<EOL>|1059,1060
ago|1060,1063
.|1063,1064
About|1065,1070
2|1071,1072
weeks|1073,1078
ago|1079,1082
she|1083,1086
also|1087,1091
began|1092,1097
taking|1098,1104
a|1105,1106
low|1107,1110
dose|1111,1115
OCP|1116,1119
in|1120,1122
<EOL>|1123,1124
order|1124,1129
to|1130,1132
treate|1133,1139
perimenopausal|1140,1154
cramping|1155,1163
.|1163,1164
On|1165,1167
the|1168,1171
second|1172,1178
week|1179,1183
she|1184,1187
<EOL>|1188,1189
started|1189,1196
to|1197,1199
have|1200,1204
spotting|1205,1213
,|1213,1214
with|1215,1219
intermittent|1220,1232
bleeding|1233,1241
and|1242,1245
LH|1246,1248
this|1249,1253
<EOL>|1254,1255
past|1255,1259
week|1260,1264
.|1264,1265
She|1266,1269
had|1270,1273
an|1274,1276
episode|1277,1284
of|1285,1287
diarrhea|1288,1296
one|1297,1300
week|1301,1305
ago|1306,1309
_|1310,1311
_|1311,1312
_|1312,1313
<EOL>|1314,1315
morning|1315,1322
)|1322,1323
,|1323,1324
that|1325,1329
was|1330,1333
nonbloody|1334,1343
and|1344,1347
resolved|1348,1356
on|1357,1359
its|1360,1363
own|1364,1367
.|1367,1368
Starting|1369,1377
<EOL>|1378,1379
on|1379,1381
_|1382,1383
_|1383,1384
_|1384,1385
she|1386,1389
has|1390,1393
had|1394,1397
a|1398,1399
feeling|1400,1407
of|1408,1410
"|1411,1412
lightheadedness|1412,1427
"|1427,1428
<EOL>|1429,1430
associated|1430,1440
with|1441,1445
diaphoresis|1446,1457
and|1458,1461
nausea|1462,1468
.|1468,1469
<EOL>|1471,1472
.|1472,1473
<EOL>|1475,1476
In|1476,1478
the|1479,1482
ED|1483,1485
,|1485,1486
initial|1487,1494
VS|1495,1497
were|1498,1502
:|1502,1503
8|1504,1505
97.2|1506,1510
88|1511,1513
117|1514,1517
/|1517,1518
64|1518,1520
18|1521,1523
100|1524,1527
%|1527,1528
.|1528,1529
Patient|1530,1537
<EOL>|1538,1539
was|1539,1542
given|1543,1548
morphine|1549,1557
4|1558,1559
mg|1560,1562
IV|1563,1565
,|1565,1566
dilaudid|1567,1575
0.5|1576,1579
mg|1580,1582
IV|1583,1585
x|1586,1587
6|1588,1589
,|1589,1590
zofran|1591,1597
4|1598,1599
mg|1600,1602
<EOL>|1603,1604
IV|1604,1606
,|1606,1607
and|1608,1611
3|1612,1613
L|1614,1615
NS.|1616,1619
She|1620,1623
underwent|1624,1633
bimanual|1634,1642
exam|1643,1647
that|1648,1652
was|1653,1656
reportedly|1657,1667
<EOL>|1668,1669
without|1669,1676
signs|1677,1682
of|1683,1685
mass|1686,1690
,|1690,1691
CMT|1692,1695
,|1695,1696
or|1697,1699
adnexal|1700,1707
tenderness|1708,1718
.|1718,1719
Labs|1720,1724
were|1725,1729
<EOL>|1730,1731
notable|1731,1738
for|1739,1742
a|1743,1744
leukocytosis|1745,1757
of|1758,1760
11|1761,1763
,|1763,1764
but|1765,1768
were|1769,1773
otherwise|1774,1783
<EOL>|1784,1785
unremarkable|1785,1797
.|1797,1798
CT|1799,1801
abdomen|1802,1809
showed|1810,1816
normal|1817,1823
appendix|1824,1832
but|1833,1836
thick|1837,1842
-|1842,1843
walled|1843,1849
<EOL>|1850,1851
cecum|1851,1856
with|1857,1861
appearance|1862,1872
of|1873,1875
possible|1876,1884
mass|1885,1889
.|1889,1890
Pelvic|1891,1897
ultrasound|1898,1908
did|1909,1912
<EOL>|1913,1914
not|1914,1917
show|1918,1922
any|1923,1926
source|1927,1933
of|1934,1936
her|1937,1940
pain|1941,1945
.|1945,1946
As|1947,1949
she|1950,1953
did|1954,1957
not|1958,1961
have|1962,1966
adequate|1967,1975
<EOL>|1976,1977
relief|1977,1983
with|1984,1988
pain|1989,1993
medications|1994,2005
,|2005,2006
she|2007,2010
was|2011,2014
admitted|2015,2023
to|2024,2026
the|2027,2030
medical|2031,2038
<EOL>|2039,2040
service|2040,2047
for|2048,2051
pain|2052,2056
control|2057,2064
.|2064,2065
<EOL>|2067,2068
.|2068,2069
<EOL>|2071,2072
Vitals|2072,2078
on|2079,2081
transfer|2082,2090
were|2091,2095
97.2|2096,2100
68|2101,2103
98|2104,2106
/|2106,2107
55|2107,2109
18|2110,2112
100|2113,2116
%|2116,2117
RA|2117,2119
<EOL>|2121,2122
.|2122,2123
<EOL>|2125,2126
On|2126,2128
the|2129,2132
floor|2133,2138
,|2138,2139
patient|2140,2147
reported|2148,2156
continued|2157,2166
_|2167,2168
_|2168,2169
_|2169,2170
pain|2171,2175
in|2176,2178
the|2179,2182
RLQ|2183,2186
,|2186,2187
<EOL>|2188,2189
along|2189,2194
with|2195,2199
some|2200,2204
mild|2205,2209
nausea|2210,2216
.|2216,2217
<EOL>|2219,2220
.|2220,2221
<EOL>|2223,2224
Review|2224,2230
of|2231,2233
systems|2234,2241
:|2241,2242
<EOL>|2244,2245
(|2245,2246
+|2246,2247
)|2247,2248
Per|2249,2252
HPI|2253,2256
<EOL>|2258,2259
(|2259,2260
-|2260,2261
)|2261,2262
Denies|2263,2269
fever|2270,2275
,|2275,2276
chills|2277,2283
,|2283,2284
night|2285,2290
sweats|2291,2297
,|2297,2298
recent|2299,2305
weight|2306,2312
loss|2313,2317
or|2318,2320
<EOL>|2321,2322
gain|2322,2326
.|2326,2327
Denies|2328,2334
headache|2335,2343
,|2343,2344
sinus|2345,2350
tenderness|2351,2361
,|2361,2362
rhinorrhea|2363,2373
or|2374,2376
<EOL>|2377,2378
congestion|2378,2388
.|2388,2389
Denied|2390,2396
cough|2397,2402
,|2402,2403
shortness|2404,2413
of|2414,2416
breath|2417,2423
.|2423,2424
Denied|2425,2431
chest|2432,2437
pain|2438,2442
<EOL>|2443,2444
or|2444,2446
tightness|2447,2456
,|2456,2457
palpitations|2458,2470
.|2470,2471
Denied|2472,2478
vomiting|2479,2487
,|2487,2488
diarrhea|2489,2497
,|2497,2498
<EOL>|2499,2500
constipation|2500,2512
or|2513,2515
BRBPR|2516,2521
.|2521,2522
No|2523,2525
dysuria|2526,2533
.|2533,2534
Denied|2535,2541
arthralgias|2542,2553
or|2554,2556
<EOL>|2557,2558
myalgias|2558,2566
.|2566,2567
<EOL>|2569,2570
<EOL>|2570,2571
<EOL>|2572,2573
Hx|2595,2597
diverticulitis|2598,2612
s|2613,2614
/|2614,2615
p|2615,2616
sigmoid|2617,2624
resection|2625,2634
_|2635,2636
_|2636,2637
_|2637,2638
<EOL>|2640,2641
Anxiety|2641,2648
<EOL>|2650,2651
Allergic|2651,2659
rhinitis|2660,2668
<EOL>|2670,2671
GERD|2671,2675
<EOL>|2677,2678
Eczema|2678,2684
<EOL>|2686,2687
Migraine|2687,2695
headaches|2696,2705
<EOL>|2707,2708
Eustacian|2708,2717
tube|2718,2722
dysfunction|2723,2734
<EOL>|2736,2737
<EOL>|2737,2738
<EOL>|2739,2740
:|2754,2755
<EOL>|2755,2756
_|2756,2757
_|2757,2758
_|2758,2759
<EOL>|2759,2760
:|2774,2775
<EOL>|2775,2776
Father|2776,2782
with|2783,2787
hx|2788,2790
of|2791,2793
colitis|2794,2801
,|2801,2802
F|2803,2804
died|2805,2809
lung|2810,2814
Ca|2815,2817
,|2817,2818
Aunt|2819,2823
with|2824,2828
breast|2829,2835
_|2836,2837
_|2837,2838
_|2838,2839
,|2839,2840
<EOL>|2841,2842
Paternal|2842,2850
GM|2851,2853
with|2854,2858
stomach|2859,2866
Ca|2867,2869
,|2869,2870
Mother|2871,2877
with|2878,2882
CHF|2883,2886
and|2887,2890
DM2|2891,2894
<EOL>|2895,2896
<EOL>|2897,2898
Vitals|2913,2919
:|2919,2920
T|2921,2922
:|2922,2923
97.6|2924,2928
BP|2929,2931
:|2931,2932
96|2933,2935
/|2935,2936
62|2936,2938
P|2939,2940
:|2940,2941
68|2942,2944
R|2945,2946
:|2946,2947
18|2947,2949
O2|2950,2952
:|2952,2953
99|2954,2956
%|2956,2957
on|2958,2960
RA|2961,2963
<EOL>|2965,2966
General|2966,2973
:|2973,2974
Alert|2975,2980
,|2980,2981
oriented|2982,2990
,|2990,2991
no|2992,2994
acute|2995,3000
distress|3001,3009
<EOL>|3011,3012
HEENT|3012,3017
:|3017,3018
Sclera|3019,3025
anicteric|3026,3035
,|3035,3036
MMM|3037,3040
,|3040,3041
oropharynx|3042,3052
clear|3053,3058
<EOL>|3060,3061
Neck|3061,3065
:|3065,3066
supple|3067,3073
,|3073,3074
JVP|3075,3078
not|3079,3082
elevated|3083,3091
,|3091,3092
no|3093,3095
LAD|3096,3099
<EOL>|3101,3102
Lungs|3102,3107
:|3107,3108
Clear|3109,3114
to|3115,3117
auscultation|3118,3130
bilaterally|3131,3142
,|3142,3143
no|3144,3146
wheezes|3147,3154
,|3154,3155
rales|3156,3161
,|3161,3162
<EOL>|3163,3164
rhonchi|3164,3171
<EOL>|3173,3174
CV|3174,3176
:|3176,3177
Regular|3178,3185
rate|3186,3190
and|3191,3194
rhythm|3195,3201
,|3201,3202
normal|3203,3209
S1|3210,3212
+|3213,3214
S2|3215,3217
,|3217,3218
no|3219,3221
murmurs|3222,3229
,|3229,3230
rubs|3231,3235
,|3235,3236
<EOL>|3237,3238
gallops|3238,3245
<EOL>|3247,3248
Abdomen|3248,3255
:|3255,3256
soft|3257,3261
,|3261,3262
non-distended|3263,3276
,|3276,3277
bowel|3278,3283
sounds|3284,3290
present|3291,3298
,|3298,3299
TTP|3300,3303
in|3304,3306
RLQ|3307,3310
<EOL>|3311,3312
with|3312,3316
deep|3317,3321
palpation|3322,3331
only|3332,3336
,|3336,3337
no|3338,3340
rebound|3341,3348
tenderness|3349,3359
or|3360,3362
guarding|3363,3371
,|3371,3372
no|3373,3375
<EOL>|3376,3377
organomegaly|3377,3389
<EOL>|3391,3392
Ext|3392,3395
:|3395,3396
Warm|3397,3401
,|3401,3402
well|3403,3407
perfused|3408,3416
,|3416,3417
2|3418,3419
+|3419,3420
pulses|3421,3427
,|3427,3428
no|3429,3431
clubbing|3432,3440
,|3440,3441
cyanosis|3442,3450
or|3451,3453
<EOL>|3454,3455
edema|3455,3460
<EOL>|3462,3463
<EOL>|3463,3464
<EOL>|3465,3466
Pertinent|3466,3475
Results|3476,3483
:|3483,3484
<EOL>|3484,3485
Laboratory|3485,3495
Findings|3496,3504
:|3504,3505
<EOL>|3505,3506
_|3506,3507
_|3507,3508
_|3508,3509
03|3510,3512
:|3512,3513
30AM|3513,3517
BLOOD|3518,3523
WBC|3524,3527
-|3527,3528
11|3528,3530
.|3530,3531
3|3531,3532
*|3532,3533
RBC|3534,3537
-|3537,3538
3|3538,3539
.|3539,3540
93|3540,3542
*|3542,3543
Hgb|3544,3547
-|3547,3548
12.2|3548,3552
Hct|3553,3556
-|3556,3557
34|3557,3559
.|3559,3560
9|3560,3561
*|3561,3562
<EOL>|3563,3564
MCV|3564,3567
-|3567,3568
89|3568,3570
MCH|3571,3574
-|3574,3575
31.0|3575,3579
MCHC|3580,3584
-|3584,3585
34.8|3585,3589
RDW|3590,3593
-|3593,3594
12.8|3594,3598
Plt|3599,3602
_|3603,3604
_|3604,3605
_|3605,3606
<EOL>|3606,3607
_|3607,3608
_|3608,3609
_|3609,3610
03|3611,3613
:|3613,3614
30AM|3614,3618
BLOOD|3619,3624
Neuts|3625,3630
-|3630,3631
76|3631,3633
.|3633,3634
5|3634,3635
*|3635,3636
_|3637,3638
_|3638,3639
_|3639,3640
Monos|3641,3646
-|3646,3647
2.8|3647,3650
Eos|3651,3654
-|3654,3655
1.8|3655,3658
<EOL>|3659,3660
Baso|3660,3664
-|3664,3665
0.4|3665,3668
<EOL>|3668,3669
_|3669,3670
_|3670,3671
_|3671,3672
05|3673,3675
:|3675,3676
26AM|3676,3680
BLOOD|3681,3686
_|3687,3688
_|3688,3689
_|3689,3690
<EOL>|3690,3691
_|3691,3692
_|3692,3693
_|3693,3694
03|3695,3697
:|3697,3698
30AM|3698,3702
BLOOD|3703,3708
Glucose|3709,3716
-|3716,3717
123|3717,3720
*|3720,3721
UreaN|3722,3727
-|3727,3728
16|3728,3730
Creat|3731,3736
-|3736,3737
0.8|3737,3740
Na|3741,3743
-|3743,3744
137|3744,3747
<EOL>|3748,3749
K|3749,3750
-|3750,3751
4.6|3751,3754
Cl|3755,3757
-|3757,3758
101|3758,3761
HCO3|3762,3766
-|3766,3767
25|3767,3769
AnGap|3770,3775
-|3775,3776
16|3776,3778
<EOL>|3778,3779
_|3779,3780
_|3780,3781
_|3781,3782
03|3783,3785
:|3785,3786
30AM|3786,3790
BLOOD|3791,3796
ALT|3797,3800
-|3800,3801
16|3801,3803
AST|3804,3807
-|3807,3808
37|3808,3810
AlkPhos|3811,3818
-|3818,3819
36|3819,3821
TotBili|3822,3829
-|3829,3830
0.5|3830,3833
<EOL>|3833,3834
_|3834,3835
_|3835,3836
_|3836,3837
03|3838,3840
:|3840,3841
30AM|3841,3845
BLOOD|3846,3851
Lipase|3852,3858
-|3858,3859
28|3859,3861
<EOL>|3861,3862
_|3862,3863
_|3863,3864
_|3864,3865
05|3866,3868
:|3868,3869
27AM|3869,3873
BLOOD|3874,3879
Calcium|3880,3887
-|3887,3888
8|3888,3889
.|3889,3890
3|3890,3891
*|3891,3892
Phos|3893,3897
-|3897,3898
2|3898,3899
.|3899,3900
0|3900,3901
*|3901,3902
#|3902,3903
Mg|3904,3906
-|3906,3907
2.0|3907,3910
<EOL>|3910,3911
_|3911,3912
_|3912,3913
_|3913,3914
03|3915,3917
:|3917,3918
39AM|3918,3922
BLOOD|3923,3928
Lactate|3929,3936
-|3936,3937
0.9|3937,3940
<EOL>|3940,3941
_|3941,3942
_|3942,3943
_|3943,3944
05|3945,3947
:|3947,3948
26AM|3948,3952
BLOOD|3953,3958
WBC|3959,3962
-|3962,3963
5.4|3963,3966
RBC|3967,3970
-|3970,3971
3|3971,3972
.|3972,3973
41|3973,3975
*|3975,3976
Hgb|3977,3980
-|3980,3981
10|3981,3983
.|3983,3984
6|3984,3985
*|3985,3986
Hct|3987,3990
-|3990,3991
30|3991,3993
.|3993,3994
6|3994,3995
*|3995,3996
<EOL>|3997,3998
MCV|3998,4001
-|4001,4002
90|4002,4004
MCH|4005,4008
-|4008,4009
31.1|4009,4013
MCHC|4014,4018
-|4018,4019
34.7|4019,4023
RDW|4024,4027
-|4027,4028
12.5|4028,4032
Plt|4033,4036
_|4037,4038
_|4038,4039
_|4039,4040
<EOL>|4040,4041
_|4041,4042
_|4042,4043
_|4043,4044
05|4045,4047
:|4047,4048
26AM|4048,4052
BLOOD|4053,4058
Glucose|4059,4066
-|4066,4067
88|4067,4069
UreaN|4070,4075
-|4075,4076
5|4076,4077
*|4077,4078
Creat|4079,4084
-|4084,4085
0.7|4085,4088
Na|4089,4091
-|4091,4092
144|4092,4095
<EOL>|4096,4097
K|4097,4098
-|4098,4099
4.1|4099,4102
Cl|4103,4105
-|4105,4106
106|4106,4109
HCO3|4110,4114
-|4114,4115
28|4115,4117
AnGap|4118,4123
-|4123,4124
14|4124,4126
<EOL>|4126,4127
_|4127,4128
_|4128,4129
_|4129,4130
03|4131,4133
:|4133,4134
30AM|4134,4138
URINE|4139,4144
Color|4145,4150
-|4150,4151
Straw|4151,4156
Appear|4157,4163
-|4163,4164
Clear|4164,4169
Sp|4170,4172
_|4173,4174
_|4174,4175
_|4175,4176
<EOL>|4176,4177
_|4177,4178
_|4178,4179
_|4179,4180
03|4181,4183
:|4183,4184
30AM|4184,4188
URINE|4189,4194
Blood|4195,4200
-|4200,4201
TR|4201,4203
Nitrite|4204,4211
-|4211,4212
NEG|4212,4215
Protein|4216,4223
-|4223,4224
NEG|4224,4227
<EOL>|4228,4229
Glucose|4229,4236
-|4236,4237
NEG|4237,4240
Ketone|4241,4247
-|4247,4248
NEG|4248,4251
Bilirub|4252,4259
-|4259,4260
NEG|4260,4263
Urobiln|4264,4271
-|4271,4272
NEG|4272,4275
pH|4276,4278
-|4278,4279
6.5|4279,4282
Leuks|4283,4288
-|4288,4289
MOD|4289,4292
<EOL>|4292,4293
_|4293,4294
_|4294,4295
_|4295,4296
03|4297,4299
:|4299,4300
30AM|4300,4304
URINE|4305,4310
RBC|4311,4314
-|4314,4315
<|4315,4316
1|4316,4317
WBC|4318,4321
-|4321,4322
3|4322,4323
Bacteri|4324,4331
-|4331,4332
FEW|4332,4335
Yeast|4336,4341
-|4341,4342
NONE|4342,4346
Epi|4347,4350
-|4350,4351
0|4351,4352
<EOL>|4352,4353
<EOL>|4353,4354
Microbiology|4354,4366
:|4366,4367
<EOL>|4367,4368
URINE|4368,4373
CULTURE|4374,4381
(|4382,4383
Final|4383,4388
_|4389,4390
_|4390,4391
_|4391,4392
:|4392,4393
<|4397,4398
10,000|4398,4404
organisms|4405,4414
/|4414,4415
ml|4415,4417
<EOL>|4417,4418
Blood|4418,4423
Culture|4424,4431
_|4432,4433
_|4433,4434
_|4434,4435
:|4435,4436
No|4437,4439
growth|4440,4446
(|4447,4448
not|4448,4451
final|4452,4457
at|4458,4460
time|4461,4465
of|4466,4468
<EOL>|4469,4470
discharge|4470,4479
)|4479,4480
<EOL>|4480,4481
<EOL>|4481,4482
Imaging|4482,4489
:|4489,4490
<EOL>|4490,4491
Pelvic|4491,4497
U|4498,4499
/|4499,4500
S|4500,4501
_|4502,4503
_|4503,4504
_|4504,4505
:|4505,4506
FINDINGS|4507,4515
:|4515,4516
Transabdominally|4517,4533
the|4534,4537
uterus|4538,4544
measures|4545,4553
<EOL>|4554,4555
8.6|4555,4558
x|4559,4560
4.6|4561,4564
x|4565,4566
5.4|4567,4570
cm|4571,4573
,|4573,4574
and|4575,4578
is|4579,4581
slightly|4582,4590
heterogeneous|4591,4604
in|4605,4607
appearance|4608,4618
<EOL>|4619,4620
with|4620,4624
no|4625,4627
distinct|4628,4636
fibroids|4637,4645
seen|4646,4650
.|4650,4651
Transvaginal|4652,4664
exam|4665,4669
was|4670,4673
performed|4674,4683
<EOL>|4684,4685
for|4685,4688
better|4689,4695
evaluation|4696,4706
of|4707,4709
the|4710,4713
uterus|4714,4720
and|4721,4724
adnexa|4725,4731
.|4731,4732
The|4733,4736
endometrial|4737,4748
<EOL>|4749,4750
stripe|4750,4756
measures|4757,4765
5|4766,4767
mm|4768,4770
.|4770,4771
The|4772,4775
left|4776,4780
ovary|4781,4786
measures|4787,4795
3.5|4796,4799
x|4800,4801
1.6|4802,4805
x|4806,4807
1.8|4808,4811
<EOL>|4812,4813
cm|4813,4815
.|4815,4816
The|4817,4820
right|4821,4826
ovary|4827,4832
measures|4833,4841
2.9|4842,4845
x|4846,4847
1.4|4848,4851
x|4852,4853
1.7|4854,4857
cm|4858,4860
.|4860,4861
There|4862,4867
is|4868,4870
a|4871,4872
<EOL>|4873,4874
small|4874,4879
echogenic|4880,4889
focus|4890,4895
within|4896,4902
the|4903,4906
right|4907,4912
ovary|4913,4918
measuring|4919,4928
5|4929,4930
x|4931,4932
4|4933,4934
x|4935,4936
4|4937,4938
<EOL>|4939,4940
mm|4940,4942
,|4942,4943
likely|4944,4950
a|4951,4952
small|4953,4958
hemorrhagic|4959,4970
cyst|4971,4975
.|4975,4976
Both|4977,4981
ovaries|4982,4989
demonstrate|4990,5001
<EOL>|5002,5003
normal|5003,5009
arterial|5010,5018
and|5019,5022
venous|5023,5029
waveforms|5030,5039
.|5039,5040
<EOL>|5043,5044
1|5058,5059
.|5059,5060
No|5061,5063
evidence|5064,5072
of|5073,5075
ovarian|5076,5083
torsion|5084,5091
.|5091,5092
<EOL>|5094,5095
2.|5095,5097
Small|5098,5103
right|5104,5109
ovarian|5110,5117
hemorrhagic|5118,5129
cyst|5130,5134
.|5134,5135
<EOL>|5136,5137
.|5137,5138
<EOL>|5138,5139
CT|5139,5141
abd|5142,5145
/|5145,5146
pelvis|5146,5152
w|5153,5154
/|5154,5155
o|5155,5156
contrast|5157,5165
_|5166,5167
_|5167,5168
_|5168,5169
:|5169,5170
Scattered|5172,5181
calcified|5182,5191
<EOL>|5192,5193
granulomas|5193,5203
in|5204,5206
<EOL>|5207,5208
the|5208,5211
lung|5212,5216
bases|5217,5222
are|5223,5226
stable|5227,5233
.|5233,5234
There|5235,5240
is|5241,5243
no|5244,5246
new|5247,5250
focal|5251,5256
pulmonary|5257,5266
<EOL>|5267,5268
nodule|5268,5274
,|5274,5275
<EOL>|5276,5277
consolidation|5277,5290
,|5290,5291
or|5292,5294
effusion|5295,5303
.|5303,5304
The|5305,5308
cardiac|5309,5316
apex|5317,5321
is|5322,5324
within|5325,5331
normal|5332,5338
<EOL>|5339,5340
limits|5340,5346
.|5346,5347
<EOL>|5349,5350
Complete|5350,5358
evaluation|5359,5369
of|5370,5372
the|5373,5376
intra-abdominal|5377,5392
viscera|5393,5400
is|5401,5403
limited|5404,5411
by|5412,5414
<EOL>|5415,5416
the|5416,5419
<EOL>|5420,5421
non-contrast|5421,5433
technique|5434,5443
.|5443,5444
However|5445,5452
,|5452,5453
the|5454,5457
liver|5458,5463
appears|5464,5471
homogeneous|5472,5483
<EOL>|5484,5485
without|5485,5492
focal|5493,5498
lesion|5499,5505
.|5505,5506
No|5507,5509
intra|5510,5515
-|5515,5516
or|5517,5519
extra-hepatic|5520,5533
biliary|5534,5541
ductal|5542,5548
<EOL>|5549,5550
dilatation|5550,5560
is|5561,5563
identified|5564,5574
.|5574,5575
The|5577,5580
gallbladder|5581,5592
,|5592,5593
spleen|5594,5600
,|5600,5601
and|5602,5605
pancreas|5606,5614
<EOL>|5615,5616
appear|5616,5622
within|5623,5629
normal|5630,5636
limits|5637,5643
.|5643,5644
The|5645,5648
adrenal|5649,5656
glands|5657,5663
are|5664,5667
symmetric|5668,5677
<EOL>|5678,5679
without|5679,5686
focal|5687,5692
nodule|5693,5699
.|5699,5700
The|5701,5704
kidneys|5705,5712
appear|5713,5719
homogeneous|5720,5731
without|5732,5739
<EOL>|5740,5741
focal|5741,5746
lesion|5747,5753
or|5754,5756
hydronephrosis|5757,5771
.|5771,5772
The|5773,5776
abdominal|5777,5786
aorta|5787,5792
is|5793,5795
<EOL>|5796,5797
non-aneurysmal|5797,5811
throughout|5812,5822
its|5823,5826
visualized|5827,5837
course|5838,5844
.|5844,5845
The|5846,5849
second|5850,5856
and|5857,5860
<EOL>|5861,5862
third|5862,5867
portions|5868,5876
of|5877,5879
the|5880,5883
duodenum|5884,5892
are|5893,5896
equivocally|5897,5908
thickened|5909,5918
which|5919,5924
<EOL>|5925,5926
may|5926,5929
be|5930,5932
due|5933,5936
to|5937,5939
underdistension|5940,5955
.|5955,5956
No|5957,5959
small|5960,5965
bowel|5966,5971
obstruction|5972,5983
is|5984,5986
<EOL>|5987,5988
identified|5988,5998
.|5998,5999
The|6000,6003
appendix|6004,6012
is|6013,6015
well|6016,6020
visualized|6021,6031
and|6032,6035
is|6036,6038
normal|6039,6045
in|6046,6048
<EOL>|6049,6050
appearance|6050,6060
.|6060,6061
There|6062,6067
is|6068,6070
no|6071,6073
free|6074,6078
fluid|6079,6084
or|6085,6087
free|6088,6092
air|6093,6096
.|6096,6097
<EOL>|6098,6099
<EOL>|6101,6102
CT|6102,6104
PELVIS|6105,6111
WITHOUT|6112,6119
INTRAVENOUS|6120,6131
CONTRAST|6132,6140
_|6141,6142
_|6142,6143
_|6143,6144
:|6144,6145
Initial|6146,6153
images|6154,6160
<EOL>|6161,6162
demonstrated|6162,6174
a|6175,6176
solid|6177,6182
mass|6183,6187
like|6188,6192
abnormality|6193,6204
in|6205,6207
the|6208,6211
cecal|6212,6217
tip|6218,6221
<EOL>|6222,6223
measuring|6223,6232
approximately|6233,6246
3|6247,6248
cm|6249,6251
(|6252,6253
2|6253,6254
:|6254,6255
51|6255,6257
)|6257,6258
.|6258,6259
As|6261,6263
this|6264,6268
was|6269,6272
potentially|6273,6284
<EOL>|6285,6286
concerning|6286,6296
for|6297,6300
a|6301,6302
cecal|6303,6308
mass|6309,6313
,|6313,6314
rescanning|6315,6325
of|6326,6328
a|6329,6330
limited|6331,6338
portion|6339,6346
of|6347,6349
<EOL>|6350,6351
pelvis|6351,6357
was|6358,6361
performed|6362,6371
after|6372,6377
passage|6378,6385
of|6386,6388
oral|6389,6393
contrast|6394,6402
,|6402,6403
confirming|6404,6414
<EOL>|6415,6416
the|6416,6419
finding|6420,6427
and|6428,6431
demonstrating|6432,6445
a|6446,6447
3|6448,6449
cm|6450,6452
mass|6453,6457
with|6458,6462
thickening|6463,6473
of|6474,6476
the|6477,6480
<EOL>|6481,6482
adjacent|6482,6490
cecal|6491,6496
wall|6497,6501
(|6502,6503
601|6503,6506
:|6506,6507
15|6507,6509
)|6509,6510
.|6510,6511
The|6512,6515
adjacent|6516,6524
appendix|6525,6533
is|6534,6536
normal|6537,6543
<EOL>|6544,6545
and|6545,6548
there|6549,6554
is|6555,6557
no|6558,6560
pericecal|6561,6570
inflammatory|6571,6583
change|6584,6590
.|6590,6591
<EOL>|6593,6594
The|6594,6597
remainder|6598,6607
of|6608,6610
the|6611,6614
colon|6615,6620
is|6621,6623
normal|6624,6630
without|6631,6638
evidence|6639,6647
of|6648,6650
<EOL>|6651,6652
obstruction|6652,6663
or|6664,6666
<EOL>|6667,6668
inflammation|6668,6680
.|6680,6681
The|6682,6685
surgical|6686,6694
anastomosis|6695,6706
within|6707,6713
the|6714,6717
lower|6718,6723
midline|6724,6731
<EOL>|6732,6733
pelvis|6733,6739
<EOL>|6740,6741
appears|6741,6748
unremarkable|6749,6761
.|6761,6762
There|6763,6768
is|6769,6771
no|6772,6774
pelvic|6775,6781
free|6782,6786
fluid|6787,6792
.|6792,6793
The|6794,6797
uterus|6798,6804
<EOL>|6805,6806
and|6806,6809
adnexa|6810,6816
<EOL>|6817,6818
appear|6818,6824
within|6825,6831
normal|6832,6838
limits|6839,6845
.|6845,6846
The|6847,6850
bladder|6851,6858
is|6859,6861
markedly|6862,6870
distended|6871,6880
<EOL>|6881,6882
but|6882,6885
is|6886,6888
<EOL>|6889,6890
otherwise|6890,6899
unremarkable|6900,6912
.|6912,6913
No|6914,6916
pathologically|6917,6931
enlarged|6932,6940
pelvic|6941,6947
or|6948,6950
<EOL>|6951,6952
inguinal|6952,6960
lymph|6961,6966
nodes|6967,6972
are|6973,6976
identified|6977,6987
.|6987,6988
<EOL>|6989,6990
OSSEOUS|6990,6997
STRUCTURES|6998,7008
:|7008,7009
No|7010,7012
bone|7013,7017
destructive|7018,7029
lesion|7030,7036
or|7037,7039
acute|7040,7045
fracture|7046,7054
<EOL>|7055,7056
is|7056,7058
<EOL>|7059,7060
identified|7060,7070
.|7070,7071
<EOL>|7073,7074
1.|7087,7089
Findings|7090,7098
consistent|7099,7109
with|7110,7114
a|7115,7116
3|7117,7118
cm|7119,7121
cecal|7122,7127
mass|7128,7132
and|7133,7136
thickening|7137,7147
of|7148,7150
<EOL>|7151,7152
the|7152,7155
cecal|7156,7161
tip|7162,7165
concerning|7166,7176
for|7177,7180
neoplasm|7181,7189
.|7189,7190
Atypical|7191,7199
infectious|7200,7210
<EOL>|7211,7212
process|7212,7219
causing|7220,7227
this|7228,7232
appearance|7233,7243
is|7244,7246
felt|7247,7251
less|7252,7256
likely|7257,7263
due|7264,7267
to|7268,7270
lack|7271,7275
<EOL>|7276,7277
of|7277,7279
inflammatory|7280,7292
stranding|7293,7302
.|7302,7303
Recommend|7304,7313
colonoscopy|7314,7325
for|7326,7329
further|7330,7337
<EOL>|7338,7339
evaluation|7339,7349
.|7349,7350
<EOL>|7352,7353
2.|7353,7355
Normal|7356,7362
appendix|7363,7371
,|7371,7372
no|7373,7375
signs|7376,7381
of|7382,7384
inflammation|7385,7397
.|7397,7398
<EOL>|7399,7400
3.|7400,7402
No|7403,7405
small|7406,7411
or|7412,7414
large|7415,7420
bowel|7421,7426
obstruction|7427,7438
.|7438,7439
<EOL>|7440,7441
4.|7441,7443
Equivocal|7444,7453
thickening|7454,7464
of|7465,7467
duodenum|7468,7476
likely|7477,7483
related|7484,7491
to|7492,7494
<EOL>|7495,7496
underdistention|7496,7511
.|7511,7512
<EOL>|7514,7515
<EOL>|7515,7516
Colonoscopy|7516,7527
_|7528,7529
_|7529,7530
_|7530,7531
:|7531,7532
<EOL>|7532,7533
:|7541,7542
<EOL>|7544,7545
Lumen|7546,7551
:|7551,7552
Evidence|7553,7561
of|7562,7564
a|7565,7566
previous|7567,7575
end|7576,7579
to|7580,7582
end|7583,7586
_|7587,7588
_|7588,7589
_|7589,7590
<EOL>|7591,7592
anastomosis|7592,7603
was|7604,7607
seen|7608,7612
at|7613,7615
the|7616,7619
sigmoid|7620,7627
colon|7628,7633
.|7633,7634
<EOL>|7636,7637
Protruding|7638,7648
Lesions|7649,7656
A|7657,7658
ulcerated|7659,7668
3|7669,7670
cm|7671,7673
mass|7674,7678
of|7679,7681
malignant|7682,7691
<EOL>|7692,7693
appearance|7693,7703
was|7704,7707
found|7708,7713
in|7714,7716
the|7717,7720
cecum|7721,7726
.|7726,7727
The|7728,7731
scope|7732,7737
traversed|7738,7747
the|7748,7751
<EOL>|7752,7753
lesion|7753,7759
.|7759,7760
Cold|7761,7765
forceps|7766,7773
biopsies|7774,7782
were|7783,7787
performed|7788,7797
for|7798,7801
histology|7802,7811
at|7812,7814
<EOL>|7815,7816
the|7816,7819
cecum|7820,7825
.|7825,7826
<EOL>|7828,7829
Excavated|7830,7839
Lesions|7840,7847
Multiple|7848,7856
diverticula|7857,7868
with|7869,7873
small|7874,7879
openings|7880,7888
were|7889,7893
<EOL>|7894,7895
seen|7895,7899
in|7900,7902
the|7903,7906
descending|7907,7917
colon|7918,7923
.|7923,7924
<EOL>|7926,7927
Impression|7927,7937
:|7937,7938
Mass|7939,7943
in|7944,7946
the|7947,7950
cecum|7951,7956
(|7957,7958
biopsy|7958,7964
)|7964,7965
<EOL>|7965,7966
Diverticulosis|7966,7980
of|7981,7983
the|7984,7987
descending|7988,7998
colon|7999,8004
<EOL>|8004,8005
Previous|8005,8013
end|8014,8017
to|8018,8020
end|8021,8024
_|8025,8026
_|8026,8027
_|8027,8028
anastomosis|8029,8040
of|8041,8043
the|8044,8047
sigmoid|8048,8055
<EOL>|8056,8057
colon|8057,8062
<EOL>|8062,8063
Otherwise|8063,8072
normal|8073,8079
colonoscopy|8080,8091
to|8092,8094
cecum|8095,8100
and|8101,8104
terminal|8105,8113
ileum|8114,8119
<EOL>|8120,8121
.|8121,8122
<EOL>|8122,8123
PATHOLOGY|8123,8132
:|8132,8133
<EOL>|8133,8134
"|8146,8147
Cecal|8147,8152
mass|8153,8157
"|8157,8158
,|8158,8159
mucosal|8160,8167
biopsies|8168,8176
:|8176,8177
<EOL>|8178,8179
Colonic|8179,8186
mucosa|8187,8193
with|8194,8198
focal|8199,8204
ischemic|8205,8213
change|8214,8220
and|8221,8224
abundant|8225,8233
<EOL>|8234,8235
associated|8235,8245
ulceration|8246,8256
,|8256,8257
exudate|8258,8265
,|8265,8266
and|8267,8270
granulation|8271,8282
tissue|8283,8289
<EOL>|8290,8291
formation|8291,8300
;|8300,8301
no|8302,8304
carcinoma|8305,8314
or|8315,8317
dysplasia|8318,8327
in|8328,8330
these|8331,8336
samples|8337,8344
.|8344,8345
Five|8347,8351
<EOL>|8352,8353
levels|8353,8359
are|8360,8363
examined|8364,8372
.|8372,8373
<EOL>|8373,8374
<EOL>|8374,8375
<EOL>|8376,8377
<EOL>|8377,8378
<EOL>|8379,8380
The|8403,8406
patient|8407,8414
is|8415,8417
a|8418,8419
_|8420,8421
_|8421,8422
_|8422,8423
year|8424,8428
-|8428,8429
old|8429,8432
female|8433,8439
with|8440,8444
history|8445,8452
significant|8453,8464
for|8465,8468
<EOL>|8469,8470
diverticulitis|8470,8484
s|8485,8486
/|8486,8487
p|8487,8488
sigmoid|8489,8496
resection|8497,8506
in|8507,8509
_|8510,8511
_|8511,8512
_|8512,8513
,|8513,8514
who|8515,8518
presented|8519,8528
with|8529,8533
<EOL>|8534,8535
abdominal|8535,8544
pain|8545,8549
and|8550,8553
was|8554,8557
found|8558,8563
to|8564,8566
have|8567,8571
cecal|8572,8577
mass|8578,8582
.|8582,8583
<EOL>|8585,8586
.|8586,8587
<EOL>|8589,8590
#|8590,8591
Abdominal|8592,8601
pain|8602,8606
:|8606,8607
Was|8608,8611
most|8612,8616
likely|8617,8623
related|8624,8631
to|8632,8634
hemorrhagic|8635,8646
ovarian|8647,8654
<EOL>|8655,8656
cyst|8656,8660
.|8660,8661
Initially|8663,8672
,|8672,8673
patient|8674,8681
had|8682,8685
significant|8686,8697
pain|8698,8702
that|8703,8707
was|8708,8711
not|8712,8715
<EOL>|8716,8717
relieved|8717,8725
with|8726,8730
dilaudid|8731,8739
.|8739,8740
However|8742,8749
,|8749,8750
over|8751,8755
the|8756,8759
course|8760,8766
of|8767,8769
several|8770,8777
<EOL>|8778,8779
days|8779,8783
her|8784,8787
pain|8788,8792
resolved|8793,8801
on|8802,8804
its|8805,8808
own|8809,8812
and|8813,8816
she|8817,8820
no|8821,8823
longer|8824,8830
required|8831,8839
any|8840,8843
<EOL>|8844,8845
pain|8845,8849
medications|8850,8861
.|8861,8862
Bloodwork|8864,8873
and|8874,8877
imaging|8878,8885
were|8886,8890
not|8891,8894
suggestive|8895,8905
of|8906,8908
<EOL>|8909,8910
any|8910,8913
intra-abdominal|8914,8929
infection|8930,8939
.|8939,8940
The|8942,8945
patient|8946,8953
was|8954,8957
advised|8958,8965
to|8966,8968
<EOL>|8969,8970
follow|8970,8976
-|8976,8977
up|8977,8979
with|8980,8984
her|8985,8988
gynecologist|8989,9001
regarding|9002,9011
her|9012,9015
ovarian|9016,9023
cyst|9024,9028
,|9028,9029
and|9030,9033
<EOL>|9034,9035
the|9035,9038
need|9039,9043
for|9044,9047
continued|9048,9057
therapy|9058,9065
with|9066,9070
low|9071,9074
dose|9075,9079
oral|9080,9084
contraceptive|9085,9098
.|9098,9099
<EOL>|9100,9101
<EOL>|9103,9104
.|9104,9105
<EOL>|9107,9108
#|9108,9109
Cecal|9110,9115
Mass|9116,9120
:|9120,9121
During|9122,9128
the|9129,9132
workup|9133,9139
of|9140,9142
this|9143,9147
patient|9148,9155
's|9155,9157
abdominal|9158,9167
<EOL>|9168,9169
pain|9169,9173
,|9173,9174
a|9175,9176
CT|9177,9179
of|9180,9182
the|9183,9186
abdomen|9187,9194
and|9195,9198
pelvis|9199,9205
revealed|9206,9214
a|9215,9216
3|9217,9218
cm|9219,9221
cecal|9222,9227
mass|9228,9232
<EOL>|9233,9234
concerning|9234,9244
for|9245,9248
malignancy|9249,9259
.|9259,9260
During|9262,9268
this|9269,9273
hospitalization|9274,9289
she|9290,9293
<EOL>|9294,9295
underwent|9295,9304
colonoscopy|9305,9316
with|9317,9321
biopsy|9322,9328
of|9329,9331
the|9332,9335
mass|9336,9340
.|9340,9341
She|9343,9346
was|9347,9350
<EOL>|9351,9352
instructed|9352,9362
to|9363,9365
follow|9366,9372
-|9372,9373
up|9373,9375
with|9376,9380
her|9381,9384
outpatient|9385,9395
gastroenterologist|9396,9414
<EOL>|9415,9416
regarding|9416,9425
the|9426,9429
results|9430,9437
of|9438,9440
this|9441,9445
biopsy|9446,9452
in|9453,9455
one|9456,9459
week|9460,9464
.|9464,9465
The|9467,9470
biopsy|9471,9477
<EOL>|9478,9479
was|9479,9482
negative|9483,9491
for|9492,9495
malignancy|9496,9506
.|9506,9507
<EOL>|9510,9511
.|9511,9512
<EOL>|9514,9515
#|9515,9516
Anxiety|9517,9524
-|9525,9526
Patient|9527,9534
was|9535,9538
continued|9539,9548
on|9549,9551
home|9552,9556
regimen|9557,9564
of|9565,9567
zoloft|9568,9574
and|9575,9578
<EOL>|9579,9580
ativan|9580,9586
.|9586,9587
<EOL>|9589,9590
.|9590,9591
<EOL>|9593,9594
#|9594,9595
Gerd|9596,9600
-|9601,9602
Patient|9603,9610
continued|9611,9620
on|9621,9623
omeprazole|9624,9634
,|9634,9635
zantac|9636,9642
BID|9643,9646
per|9647,9650
<EOL>|9651,9652
outpatient|9652,9662
regimen|9663,9670
.|9670,9671
<EOL>|9673,9674
<EOL>|9674,9675
<EOL>|9676,9677
Medications|9677,9688
on|9689,9691
Admission|9692,9701
:|9701,9702
<EOL>|9702,9703
-|9703,9704
Fish|9704,9708
Oil|9709,9712
1,000|9713,9718
mg|9719,9721
Cap|9722,9725
<EOL>|9727,9728
-|9728,9729
Axert|9729,9734
12.5|9735,9739
mg|9740,9742
Tab|9743,9746
<EOL>|9748,9749
1|9749,9750
Tablet|9751,9757
(|9757,9758
s|9758,9759
)|9759,9760
by|9761,9763
mouth|9764,9769
at|9770,9772
onset|9773,9778
of|9779,9781
HA|9782,9784
may|9785,9788
repeat|9789,9795
in|9796,9798
2|9799,9800
hour|9801,9805
up|9806,9808
till|9809,9813
<EOL>|9814,9815
2|9815,9816
a|9817,9818
day|9819,9822
<EOL>|9824,9825
-|9825,9826
Lexapro|9826,9833
10|9834,9836
mg|9837,9839
Tab|9840,9843
daily|9844,9849
<EOL>|9851,9852
-|9852,9853
Cholecalciferol|9853,9868
(|9869,9870
Vitamin|9870,9877
D3|9878,9880
)|9880,9881
1,000|9882,9887
unit|9888,9892
Tab|9893,9896
<EOL>|9898,9899
-|9899,9900
lorazepam|9900,9909
0.5|9910,9913
mg|9914,9916
Tab|9917,9920
qd|9921,9923
prn|9924,9927
<EOL>|9929,9930
-|9930,9931
Omeprazole|9931,9941
20|9942,9944
mg|9945,9947
Cap|9948,9951
,|9951,9952
Delayed|9953,9960
Release|9961,9968
BID|9969,9972
<EOL>|9974,9975
-|9975,9976
tramadol|9976,9984
50|9985,9987
mg|9988,9990
Tab|9991,9994
every|9995,10000
six|10001,10004
(|10005,10006
6|10006,10007
)|10007,10008
hours|10009,10014
as|10015,10017
needed|10018,10024
for|10025,10028
pain|10029,10033
<EOL>|10035,10036
-|10036,10037
oxycodone|10037,10046
5|10047,10048
mg|10049,10051
Tab|10052,10055
<EOL>|10057,10058
_|10058,10059
_|10059,10060
_|10060,10061
Tablet|10062,10068
(|10068,10069
s|10069,10070
)|10070,10071
by|10072,10074
mouth|10075,10080
qhs|10081,10084
prn|10085,10088
as|10089,10091
needed|10092,10098
for|10099,10102
pain|10103,10107
<EOL>|10109,10110
-|10110,10111
Multivitamin|10111,10123
Cap|10124,10127
<EOL>|10129,10130
-|10130,10131
Zantac|10131,10137
150|10138,10141
mg|10142,10144
Cap|10145,10148
1|10149,10150
Capsule|10151,10158
(|10158,10159
s|10159,10160
)|10160,10161
by|10162,10164
mouth|10165,10170
twice|10171,10176
a|10177,10178
day|10179,10182
<EOL>|10184,10185
-|10185,10186
Fluticasone|10186,10197
50|10198,10200
mcg|10201,10204
/|10204,10205
Actuation|10205,10214
Nasal|10215,10220
Spray|10221,10226
,|10226,10227
Susp|10228,10232
<EOL>|10234,10235
2|10235,10236
sprays|10237,10243
(|10243,10244
s|10244,10245
)|10245,10246
intranasally|10247,10259
for|10260,10263
7d|10264,10266
,|10266,10267
then|10268,10272
1|10273,10274
spray|10275,10280
qd|10281,10283
<EOL>|10285,10286
-|10286,10287
Calcium|10287,10294
Citrate|10295,10302
1,000|10303,10308
mg|10309,10311
Tab|10312,10315
<EOL>|10317,10318
-|10318,10319
OCPs|10319,10323
-|10324,10325
Camrasce|10326,10334
?|10334,10335
started|10336,10343
2|10344,10345
weeks|10346,10351
ago|10352,10355
<EOL>|10357,10358
<EOL>|10358,10359
<EOL>|10360,10361
Discharge|10361,10370
Medications|10371,10382
:|10382,10383
<EOL>|10383,10384
1.|10384,10386
omega|10387,10392
-|10392,10393
3|10393,10394
fatty|10395,10400
acids|10401,10406
Capsule|10411,10418
Sig|10419,10422
:|10422,10423
One|10424,10427
(|10428,10429
1|10429,10430
)|10430,10431
Capsule|10432,10439
PO|10440,10442
DAILY|10443,10448
<EOL>|10449,10450
(|10450,10451
Daily|10451,10456
)|10456,10457
.|10457,10458
<EOL>|10460,10461
2.|10461,10463
Axert|10464,10469
12.5|10470,10474
mg|10475,10477
Tablet|10478,10484
Sig|10485,10488
:|10488,10489
One|10490,10493
(|10494,10495
1|10495,10496
)|10496,10497
Tablet|10498,10504
PO|10505,10507
once|10508,10512
a|10513,10514
day|10515,10518
as|10519,10521
<EOL>|10522,10523
needed|10523,10529
for|10530,10533
migraine|10534,10542
.|10542,10543
<EOL>|10545,10546
3.|10546,10548
escitalopram|10549,10561
10|10562,10564
mg|10565,10567
Tablet|10568,10574
Sig|10575,10578
:|10578,10579
One|10580,10583
(|10584,10585
1|10585,10586
)|10586,10587
Tablet|10588,10594
PO|10595,10597
DAILY|10598,10603
<EOL>|10604,10605
(|10605,10606
Daily|10606,10611
)|10611,10612
.|10612,10613
<EOL>|10615,10616
4.|10616,10618
cholecalciferol|10619,10634
(|10635,10636
vitamin|10636,10643
D3|10644,10646
)|10646,10647
1,000|10648,10653
unit|10654,10658
Capsule|10659,10666
Sig|10667,10670
:|10670,10671
One|10672,10675
(|10676,10677
1|10677,10678
)|10678,10679
<EOL>|10680,10681
Capsule|10681,10688
PO|10689,10691
once|10692,10696
a|10697,10698
day|10699,10702
.|10702,10703
<EOL>|10705,10706
5.|10706,10708
lorazepam|10709,10718
0.5|10719,10722
mg|10723,10725
Tablet|10726,10732
Sig|10733,10736
:|10736,10737
One|10738,10741
(|10742,10743
1|10743,10744
)|10744,10745
Tablet|10746,10752
PO|10753,10755
HS|10756,10758
(|10759,10760
at|10760,10762
<EOL>|10763,10764
bedtime|10764,10771
)|10771,10772
as|10773,10775
needed|10776,10782
for|10783,10786
anxiety|10787,10794
.|10794,10795
<EOL>|10797,10798
6.|10798,10800
omeprazole|10801,10811
20|10812,10814
mg|10815,10817
Capsule|10818,10825
,|10825,10826
Delayed|10827,10834
Release|10835,10842
(|10842,10843
E.C|10843,10846
.|10846,10847
)|10847,10848
Sig|10849,10852
:|10852,10853
One|10854,10857
(|10858,10859
1|10859,10860
)|10860,10861
<EOL>|10862,10863
Capsule|10863,10870
,|10870,10871
Delayed|10872,10879
Release|10880,10887
(|10887,10888
E.C|10888,10891
.|10891,10892
)|10892,10893
PO|10894,10896
BID|10897,10900
(|10901,10902
2|10902,10903
times|10904,10909
a|10910,10911
day|10912,10915
)|10915,10916
.|10916,10917
<EOL>|10919,10920
7.|10920,10922
multivitamin|10923,10935
Tablet|10940,10946
Sig|10947,10950
:|10950,10951
One|10952,10955
(|10956,10957
1|10957,10958
)|10958,10959
Tablet|10960,10966
PO|10967,10969
DAILY|10970,10975
(|10976,10977
Daily|10977,10982
)|10982,10983
.|10983,10984
<EOL>|10985,10986
<EOL>|10987,10988
8.|10988,10990
ranitidine|10991,11001
HCl|11002,11005
150|11006,11009
mg|11010,11012
Tablet|11013,11019
Sig|11020,11023
:|11023,11024
One|11025,11028
(|11029,11030
1|11030,11031
)|11031,11032
Tablet|11033,11039
PO|11040,11042
BID|11043,11046
(|11047,11048
2|11048,11049
<EOL>|11050,11051
times|11051,11056
a|11057,11058
day|11059,11062
)|11062,11063
.|11063,11064
<EOL>|11066,11067
9.|11067,11069
fluticasone|11070,11081
50|11082,11084
mcg|11085,11088
/|11088,11089
Actuation|11089,11098
Spray|11099,11104
,|11104,11105
Suspension|11106,11116
Sig|11117,11120
:|11120,11121
One|11122,11125
(|11126,11127
1|11127,11128
)|11128,11129
<EOL>|11130,11131
Spray|11131,11136
Nasal|11137,11142
DAILY|11143,11148
(|11149,11150
Daily|11150,11155
)|11155,11156
.|11156,11157
<EOL>|11159,11160
10.|11160,11163
calcium|11164,11171
carbonate|11172,11181
500|11182,11185
mg|11186,11188
calcium|11189,11196
(|11197,11198
1,250|11198,11203
mg|11204,11206
)|11206,11207
Tablet|11208,11214
Sig|11215,11218
:|11218,11219
Two|11220,11223
<EOL>|11224,11225
(|11225,11226
2|11226,11227
)|11227,11228
Tablet|11229,11235
PO|11236,11238
once|11239,11243
a|11244,11245
day|11246,11249
.|11249,11250
<EOL>|11252,11253
<EOL>|11253,11254
<EOL>|11255,11256
Discharge|11256,11265
Disposition|11266,11277
:|11277,11278
<EOL>|11278,11279
Home|11279,11283
<EOL>|11283,11284
<EOL>|11285,11286
Discharge|11286,11295
Diagnosis|11296,11305
:|11305,11306
<EOL>|11306,11307
Cecal|11307,11312
Mass|11313,11317
<EOL>|11317,11318
Hemorrhagic|11318,11329
ovarian|11330,11337
cyst|11338,11342
<EOL>|11342,11343
<EOL>|11343,11344
<EOL>|11345,11346
Mental|11367,11373
Status|11374,11380
:|11380,11381
Clear|11382,11387
and|11388,11391
coherent|11392,11400
.|11400,11401
<EOL>|11401,11402
Level|11402,11407
of|11408,11410
Consciousness|11411,11424
:|11424,11425
Alert|11426,11431
and|11432,11435
interactive|11436,11447
.|11447,11448
<EOL>|11448,11449
Activity|11449,11457
Status|11458,11464
:|11464,11465
Ambulatory|11466,11476
-|11477,11478
Independent|11479,11490
.|11490,11491
<EOL>|11491,11492
<EOL>|11492,11493
<EOL>|11494,11495
Dear|11519,11523
Ms.|11524,11527
_|11528,11529
_|11529,11530
_|11530,11531
,|11531,11532
<EOL>|11532,11533
<EOL>|11533,11534
You|11534,11537
were|11538,11542
admitted|11543,11551
to|11552,11554
the|11555,11558
hospital|11559,11567
for|11568,11571
abdominal|11572,11581
pain|11582,11586
,|11586,11587
which|11588,11593
we|11594,11596
<EOL>|11597,11598
think|11598,11603
was|11604,11607
related|11608,11615
to|11616,11618
a|11619,11620
hemorrhagic|11621,11632
ovarian|11633,11640
cyst|11641,11645
.|11645,11646
You|11648,11651
were|11652,11656
<EOL>|11657,11658
treated|11658,11665
with|11666,11670
analgesics|11671,11681
,|11681,11682
and|11683,11686
your|11687,11691
pain|11692,11696
resolved|11697,11705
.|11705,11706
You|11708,11711
also|11712,11716
had|11717,11720
a|11721,11722
<EOL>|11723,11724
CAT|11724,11727
scan|11728,11732
showing|11733,11740
a|11741,11742
mass|11743,11747
in|11748,11750
the|11751,11754
cecum|11755,11760
.|11760,11761
You|11763,11766
underwent|11767,11776
a|11777,11778
<EOL>|11779,11780
colonoscopy|11780,11791
to|11792,11794
biopsy|11795,11801
this|11802,11806
mass|11807,11811
,|11811,11812
and|11813,11816
you|11817,11820
should|11821,11827
follow|11828,11834
-|11834,11835
up|11835,11837
with|11838,11842
<EOL>|11843,11844
your|11844,11848
gastroenterologist|11849,11867
.|11867,11868
<EOL>|11869,11870
<EOL>|11870,11871
You|11871,11874
should|11875,11881
also|11882,11886
see|11887,11890
your|11891,11895
gynecologist|11896,11908
regarding|11909,11918
the|11919,11922
need|11923,11927
to|11928,11930
<EOL>|11931,11932
restart|11932,11939
your|11940,11944
oral|11945,11949
contraceptive|11950,11963
.|11963,11964
<EOL>|11964,11965
<EOL>|11965,11966
We|11966,11968
did|11969,11972
not|11973,11976
make|11977,11981
any|11982,11985
changes|11986,11993
to|11994,11996
your|11997,12001
home|12002,12006
medications|12007,12018
.|12018,12019
<EOL>|12020,12021
<EOL>|12022,12023
Followup|12023,12031
Instructions|12032,12044
:|12044,12045
<EOL>|12045,12046
_|12046,12047
_|12047,12048
_|12048,12049
<EOL>|12049,12050

