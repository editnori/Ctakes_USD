CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|Known|Modifier|false|false||Knownnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Adverse reaction to drug|Finding|true|false||Adverse Drug Reactionsnull|Adverse reaction to drug|Finding|true|false||Drug Reactionsnull|Pharmaceutical Preparations|Drug|false|false||Drug
null|Pharmacologic Substance|Drug|false|false||Drugnull|Drug problem|Finding|false|false||Drugnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Fever|Finding|false|false||Feversnull|Chills|Finding|false|false||chillsnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|null|Device|false|false||stentnull|degree of relationship - exchange|Finding|false|false||exchangenull|Exchange (clinical)|Attribute|false|false||exchangenull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|Medical History|Finding|false|false||medical historynull|Medical referral type|Finding|false|false||medical
null|Medical|Finding|false|false||medical
null|Medical school type|Finding|false|false||medicalnull|Medical service|Procedure|false|false||medicalnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Malignant neoplasm of urinary bladder|Disorder|true|false|C0005682|bladder cancer
null|Carcinoma of bladder|Disorder|true|false|C0005682|bladder cancer
null|Bladder Neoplasm|Disorder|true|false|C0005682|bladder cancernull|Neoplasm of uncertain or unknown behavior of bladder|Disorder|false|false|C0005682|bladder
null|Benign neoplasm of bladder|Disorder|false|false|C0005682|bladder
null|Carcinoma in situ of bladder|Disorder|false|false|C0005682|bladdernull|Procedures on bladder|Procedure|false|false|C0005682|bladdernull|Urinary Bladder|Anatomy|false|false|C0872388;C0496930;C0154017;C0154091;C0006826;C0699885;C0005684;C0005695|bladdernull|Malignant Neoplasms|Disorder|false|false|C0005682|cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|SLC35G1 gene|Finding|false|false||post
null|DESI1 gene|Finding|false|false||postnull|Post Device|Device|false|false||postnull|Post|Time|false|false||postnull|Robotics|Subject|false|false||roboticnull|Total abdominal hysterectomy|Procedure|false|false||TAHnull|Tahitian language|Entity|false|false||TAHnull|Buthionine Sulfoximine|Drug|false|false||BSO
null|Buthionine Sulfoximine|Drug|false|false||BSO
null|Buthionine Sulfoximine|Drug|false|false||BSOnull|ACP2 protein, human|Drug|false|false||lap
null|ACP2 protein, human|Drug|false|false||lapnull|Congenital laryngeal adductor palsy|Disorder|false|false||lapnull|Left atrial pressure|Finding|false|false||lap
null|ACP2 gene|Finding|false|false||lap
null|PICALM wt Allele|Finding|false|false||lap
null|LAP3 wt Allele|Finding|false|false||lap
null|ACP2 wt Allele|Finding|false|false||lap
null|LAP3 gene|Finding|false|false||lap
null|CENPJ gene|Finding|false|false||lap
null|CEBPB wt Allele|Finding|false|false||lap
null|PICALM gene|Finding|false|false||lap
null|CEBPB gene|Finding|false|false||lapnull|Laparoscopy|Procedure|false|false||lapnull|Lap - unit|LabModifier|false|false||lapnull|Complete cystectomy|Procedure|false|false||radical cystectomynull|Radicals (chemistry)|Drug|false|false||radicalnull|Radical (qualifier value)|Modifier|false|false||radicalnull|Cystectomy|Procedure|false|false||cystectomynull|Ileal Loop|Anatomy|false|false||ileal loopnull|ileum|Anatomy|false|false||ilealnull|Loop|Modifier|false|false||loopnull|null|Finding|false|false||diversion
null|Diversion|Finding|false|false||diversionnull|Diversion procedure|Procedure|false|false||diversionnull|Adenohypophyseal Diseases|Disorder|false|false||anteriornull|Anterior|Modifier|false|false||anteriornull|Vaginectomy|Procedure|false|false||vaginectomynull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Clinical act of insertion|Procedure|false|false||placement
null|Implantation procedure|Procedure|false|false||placement
null|null|Procedure|false|false||placementnull|Placement|Modifier|false|false||placementnull|null|Device|false|false||drainage cathetersnull|Body Fluid Discharge|Finding|false|false||drainage
null|Body Substance Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|catheter device|Device|false|false||cathetersnull|Further|Modifier|false|false||furthernull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Bilateral hydronephrosis|Disorder|false|false||bilateral hydronephrosisnull|Bilateral|Modifier|false|false||bilateralnull|Hydronephrosis|Disorder|false|false||hydronephrosisnull|Bilateral|Modifier|false|false||bilateralnull|Urostomy procedure|Procedure|false|false|C0559495|urostomynull|Urological stoma|Anatomy|false|false|C1533810;C0441587;C0021107;C0856443;C0883304;C1427122;C1719071|urostomynull|placement of tube|Procedure|false|false|C0559495|tube placementnull|Unspecified tube|Finding|false|false|C0559495|tube
null|TUBE1 gene|Finding|false|false|C0559495|tubenull|biomedical tube device|Device|false|false||tube
null|Packaging Tube|Device|false|false||tubenull|tube|Modifier|false|false||tubenull|Tube (unit of presentation)|LabModifier|false|false||tube
null|Tube Dosing Unit|LabModifier|false|false||tubenull|null|Procedure|false|false|C0559495|placement
null|Implantation procedure|Procedure|false|false|C0559495|placement
null|Clinical act of insertion|Procedure|false|false|C0559495|placementnull|Placement|Modifier|false|false||placementnull|Then - dosing instruction fragment|Finding|false|false|C0041951|thennull|Then|Time|false|false||thennull|Ureteral Route of Administration|Finding|false|false|C0041951|ureteralnull|Ureter|Anatomy|false|false|C1720594;C1522613|ureteralnull|null|Device|false|false||stentnull|Clinical act of insertion|Procedure|false|false||placementsnull|Improvement|Finding|false|false||improvementnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Extended Priority Codes - Routine|Finding|false|false||routine
null|Report priority - Routine|Finding|false|false||routine
null|Admission Type - Routine|Finding|false|false||routine
null|Level of Care - Routine|Finding|false|false||routine
null|Processing priority - Routine|Finding|false|false||routine
null|Referral priority - Routine|Finding|false|false||routinenull|Routine coag|Procedure|false|false||routinenull|Priority - Routine|Time|false|false||routinenull|Routine|Modifier|false|false||routinenull|null|Device|false|false||stentnull|degree of relationship - exchange|Finding|false|false||exchangenull|Exchange (clinical)|Attribute|false|false||exchangenull|Cystoscopy|Procedure|false|false||cystoscopynull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Uncomplicated|Modifier|false|false||uncomplicatednull|Procedure (set of actions)|Finding|false|false||procedurenull|Interventional procedure|Procedure|false|false||procedurenull|null|Attribute|false|false||procedurenull|Act Class - procedure|Event|false|false||procedurenull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Recovery Room|Device|false|false||PACUnull|Recovery Room|Entity|false|false||PACUnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Patient need for (contextual qualifier)|Finding|false|false||neednull|Needs|Modifier|false|false||neednull|Admission for treatment|Procedure|false|false||admission for treatmentnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|Sepsis|Disorder|false|false||sepsis
null|Septicemia|Disorder|false|false||sepsisnull|Sepsis <Sepsidae>|Entity|false|false||sepsisnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|ampicillin|Drug|false|false||ampicillin
null|ampicillins|Drug|false|false||ampicillin
null|ampicillins|Drug|false|false||ampicillin
null|ampicillin|Drug|false|false||ampicillinnull|gentamicin|Drug|false|false||gentamicin
null|gentamicin|Drug|false|false||gentamicinnull|Gentamicin measurement|Procedure|false|false||gentamicinnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Pharmaceutical Preparations|Drug|false|false||drug
null|Pharmacologic Substance|Drug|false|false||drugnull|Drug problem|Finding|false|false||drugnull|resistant - Observation Interpretation Susceptibility|Finding|false|false||resistant
null|Resistant (qualifier value)|Finding|false|false||resistantnull|Antimicrobial Resistance Result|Lab|false|false||resistantnull|Organism|Entity|false|false||organismsnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Feeling feverish|Finding|false|false||feeling feverishnull|Fever|Finding|false|false||feverishnull|Chills|Finding|false|false||chillsnull|Nausea and vomiting|Finding|false|false||nausea and vomitingnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Vomiting|Finding|false|false||vomitingnull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Medical service|Procedure|false|false||medical service
null|Physician service|Procedure|false|false||medical servicenull|Hospital Service - Medical Service|Entity|false|false||medical servicenull|Medical referral type|Finding|false|false||medical
null|Medical|Finding|false|false||medical
null|Medical school type|Finding|false|false||medicalnull|Medical service|Procedure|false|false||medicalnull|ActInformationPrivacyReason - service|Finding|false|false||servicenull|Software Service|Device|false|false||servicenull|Services|Event|false|false||servicenull|Further|Modifier|false|false||furthernull|Evaluation and management note|Finding|false|false||evaluation and managementnull|Evaluation and Management|Procedure|false|false||evaluation and managementnull|Processing type - Evaluation|Finding|false|false||evaluationnull|Evaluation procedure|Procedure|false|false||evaluation
null|Evaluation|Procedure|false|false||evaluationnull|Disease Management|Procedure|false|false||managementnull|Management Occupations|Subject|false|false||managementnull|Management procedure|Event|false|false||management
null|Administration occupational activities|Event|false|false||managementnull|Floor (anatomic)|Anatomy|false|false|C1578483;C1550655;C1578481;C1578486;C1578484;C1578485|floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Relationship modifier - Patient|Finding|false|false|C3714591|patient
null|Specimen Type - Patient|Finding|false|false|C3714591|patient
null|Mail Claim Party - Patient|Finding|false|false|C3714591|patient
null|Report source - Patient|Finding|false|false|C3714591|patient
null|null|Finding|false|false|C3714591|patient
null|Disabled Person Code - Patient|Finding|false|false|C3714591|patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Persistent|Time|false|false||persistentnull|Chills|Finding|false|false||chillsnull|Slightly (qualifier value)|Modifier|false|false||slightly
null|Slight (qualifier value)|Modifier|false|false||slightlynull|Nausea|Finding|false|false||nauseousnull|Abdominal Pain|Finding|false|false|C0000726|abdominal painnull|Abdomen|Anatomy|false|false|C0000737;C1549543;C0030193|abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Administration Method - Pain|Finding|false|false|C0000726|pain
null|Pain|Finding|false|false|C0000726|painnull|null|Attribute|false|false||painnull|Feelings|Finding|false|false||feelingnull|Observation Interpretation - better|Finding|false|false||betternull|Better|Modifier|false|false||betternull|Stat (do immediately)|Time|false|false||immediatelynull|Still|Disorder|false|false||stillnull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Medical History|Finding|false|false|C0042027;C1508753|history ofnull|History of present illness (finding)|Finding|false|false|C0042027;C0042027;C1508753;C1185740|history
null|History of previous events|Finding|false|false|C0042027;C0042027;C1508753;C1185740|history
null|Historical aspects qualifier|Finding|false|false|C0042027;C0042027;C1508753;C1185740|history
null|Medical History|Finding|false|false|C0042027;C0042027;C1508753;C1185740|history
null|Concept History|Finding|false|false|C0042027;C0042027;C1508753;C1185740|historynull|History|Subject|false|false||historynull|Recurrent urinary tract infection|Disorder|false|false|C0042027;C0042027;C1508753;C1185740|urinary tract infections
null|Urinary tract infection|Disorder|false|false|C0042027;C0042027;C1508753;C1185740|urinary tract infectionsnull|Urinary tract|Anatomy|false|false|C0042029;C0262655;C3714514;C0851162;C0262926;C1705255;C0019665;C0262512;C2004062;C0262926|urinary tract
null|Urinary system|Anatomy|false|false|C0042029;C0262655;C3714514;C0851162;C0262926;C1705255;C0019665;C0262512;C2004062;C0262926|urinary tractnull|Urinary tract|Anatomy|false|false|C0042029;C0262655;C0851162;C0262926;C1705255;C0019665;C0262512;C2004062|urinarynull|urinary|Modifier|false|false||urinarynull|Tract|Anatomy|false|false|C3714514;C0851162;C0262926;C1705255;C0019665;C0262512;C2004062;C0042029;C0262655|tractnull|Infection of musculoskeletal system|Disorder|false|false|C0042027;C0042027;C1508753;C1185740|infectionsnull|Infection|Finding|false|false|C1185740;C0042027;C1508753|infectionsnull|Recent|Time|false|false||recentlynull|ciprofloxacin|Drug|false|false||ciprofloxacin
null|ciprofloxacin|Drug|false|false||ciprofloxacinnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Course|Time|false|false||coursenull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Complaint (finding)|Finding|false|false||complaintsnull|Hypertensive disease|Disorder|false|false||Hypertensionnull|ACP2 protein, human|Drug|false|false||lap
null|ACP2 protein, human|Drug|false|false||lapnull|Congenital laryngeal adductor palsy|Disorder|false|false||lapnull|Left atrial pressure|Finding|false|false||lap
null|ACP2 gene|Finding|false|false||lap
null|PICALM wt Allele|Finding|false|false||lap
null|LAP3 wt Allele|Finding|false|false||lap
null|ACP2 wt Allele|Finding|false|false||lap
null|LAP3 gene|Finding|false|false||lap
null|CENPJ gene|Finding|false|false||lap
null|CEBPB wt Allele|Finding|false|false||lap
null|PICALM gene|Finding|false|false||lap
null|CEBPB gene|Finding|false|false||lapnull|Laparoscopy|Procedure|false|false||lapnull|Lap - unit|LabModifier|false|false||lapnull|Structure of left knee region|Anatomy|false|false|C1555302;C0035139;C0559956;C1552822;C0086511;C0562271|left knee
null|Structure of left knee|Anatomy|false|false|C1555302;C0035139;C0559956;C1552822;C0086511;C0562271|left kneenull|Table Cell Horizontal Align - left|Finding|false|false|C0230432;C4281599|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Knee Replacement Arthroplasty|Procedure|false|false|C0230432;C4281599;C1963703;C0022742;C4299094;C0022745|knee replacementnull|null|Attribute|false|false|C1963703;C0022742;C4299094;C0022745|knee replacementnull|Examination of knee joint|Procedure|false|false|C1963703;C0022742;C4299094;C0022745;C0230432;C4281599|kneenull|Knee region structure|Anatomy|false|false|C5575606;C0086511;C0562271|knee
null|Knee|Anatomy|false|false|C5575606;C0086511;C0562271|knee
null|Lower extremity>Knee|Anatomy|false|false|C5575606;C0086511;C0562271|knee
null|Knee joint|Anatomy|false|false|C5575606;C0086511;C0562271|kneenull|Replacement|Finding|false|false|C0230432;C4281599|replacementnull|Replacement - supply|Procedure|false|false|C0230432;C4281599|replacement
null|Surgical Replantation|Procedure|false|false|C0230432;C4281599|replacementnull|Laminectomy|Procedure|false|false||laminectomynull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|Malignant neoplasm of urinary bladder|Disorder|false|false|C0005682|Bladder Cancer
null|Carcinoma of bladder|Disorder|false|false|C0005682|Bladder Cancer
null|Bladder Neoplasm|Disorder|false|false|C0005682|Bladder Cancernull|Carcinoma in situ of bladder|Disorder|false|false|C0005682|Bladder
null|Benign neoplasm of bladder|Disorder|false|false|C0005682|Bladder
null|Neoplasm of uncertain or unknown behavior of bladder|Disorder|false|false|C0005682|Bladdernull|Procedures on bladder|Procedure|false|false|C0005682|Bladdernull|Urinary Bladder|Anatomy|false|false|C0699885;C0005684;C0005695;C0006826;C3887512;C5200928;C1561958;C4522209;C5202936;C0872388;C1861305;C0919553;C3244287;C0441800;C0496930;C0154017;C0154091;C4554016;C0205082|Bladdernull|Malignant Neoplasms|Disorder|false|false|C0005682|Cancernull|Specialty Type - cancer|Title|false|false||Cancernull|Cancer <Cancridae>|Entity|false|false||Cancernull|Enneking High Surgical Grade|Finding|false|false|C1167383;C0005682|high grade
null|Severe (severity modifier)|Finding|false|false|C1167383;C0005682|high gradenull|Message Waiting Priority - High|Finding|false|false|C0005682;C1167383|high
null|high - ActExposureLevelCode|Finding|false|false|C0005682;C1167383|high
null|IPSS Risk Category High|Finding|false|false|C0005682;C1167383|high
null|IPSS-R Risk Category High|Finding|false|false|C0005682;C1167383|high
null|High (finding)|Finding|false|false|C0005682;C1167383|highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Histopathologic Grade|Finding|false|false|C0005682;C1167383|grade
null|Grade|Finding|false|false|C0005682;C1167383|grade
null|School Grade|Finding|false|false|C0005682;C1167383|gradenull|Membrane Attack Complex|Drug|false|false|C1167383|TCC
null|triclocarban|Drug|false|false|C1167383|TCC
null|triclocarban|Drug|false|false|C1167383|TCC
null|Membrane Attack Complex|Drug|false|false|C1167383|TCCnull|TARSAL-CARPAL COALITION SYNDROME|Disorder|false|false|C1167383;C0005682|TCCnull|membrane attack complex location|Anatomy|false|false|C1861305;C5552697;C0077072;C4554016;C0205082;C3887512;C5200928;C1561958;C4522209;C5202936;C0919553;C3244287;C0441800|TCCnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Magnetic Resonance Imaging (MRI) of Pelvis|Procedure|false|false|C0030797|pelvic MRInull|Pelvis|Anatomy|false|false|C0024485;C0587658;C1824234;C0203201|pelvicnull|CYREN gene|Finding|false|false|C0030797|MRInull|Magnetic resonance imaging service|Procedure|false|false|C0030797|MRI
null|Magnetic Resonance Imaging|Procedure|false|false|C0030797|MRInull|Maori Language|Entity|false|false||MRInull|Tumor Cell Invasion|Disorder|false|false||invasionnull|Cell Invasion|Finding|false|false||invasionnull|Into urinary bladder|Modifier|false|false||into bladdernull|Wall of bladder|Anatomy|false|false|C0496930;C0154017;C0154091;C0872388|bladder wallnull|Neoplasm of uncertain or unknown behavior of bladder|Disorder|false|false|C0458421;C0005682|bladder
null|Benign neoplasm of bladder|Disorder|false|false|C0458421;C0005682|bladder
null|Carcinoma in situ of bladder|Disorder|false|false|C0458421;C0005682|bladdernull|Procedures on bladder|Procedure|false|false|C0005682;C0458421|bladdernull|Urinary Bladder|Anatomy|false|false|C0872388;C0496930;C0154017;C0154091|bladdernull|Walls of a building|Device|false|false||wallnull|Neck+Chest>Soft tissue|Anatomy|false|false|C0751437;C4521343;C1522570;C1547928;C3542022|soft tissue
null|soft tissue|Anatomy|false|false|C0751437;C4521343;C1522570;C1547928;C3542022|soft tissuenull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false|C0040300;C0225317;C4532079|softnull|Soft|Modifier|false|false||softnull|Tissue Specimen Code|Finding|false|false|C0225317;C4532079;C0040300|tissuenull|Body tissue|Anatomy|false|false|C3542022;C0751437;C1547928;C4521343;C1522570|tissuenull|Adenohypophyseal Diseases|Disorder|false|false|C0225317;C4532079;C0447612;C0040300|anteriornull|Anterior|Modifier|false|false||anteriornull|Vaginal wall|Anatomy|false|false|C0751437;C0332305;C4521343;C1522570|vaginal wallnull|Vaginal Dosage Form|Drug|false|false|C0042232|vaginalnull|Vaginal Route of Administration|Finding|false|false|C0225317;C4532079;C0042232;C0447612;C0040300|vaginal
null|Vaginal (intended site)|Finding|false|false|C0225317;C4532079;C0042232;C0447612;C0040300|vaginalnull|Vagina|Anatomy|false|false|C4521343;C1522570;C1272941|vaginalnull|Vaginal|Modifier|false|false||vaginalnull|Walls of a building|Device|false|false||wallnull|With staging|Finding|false|false|C0447612|stagingnull|Consent Type - Hysterectomy|Finding|false|false||hysterectomynull|Hysterectomy|Procedure|false|false||hysterectomynull|Bilateral oophorectomy|Procedure|false|false|C4266525;C0042149;C1519876|bilateral oophorectomynull|Bilateral|Modifier|false|false||bilateralnull|Ovariectomy|Procedure|false|false|C4266525;C0042149;C1519876|oophorectomynull|Enlarged uterus|Finding|false|false|C4266525;C0042149;C1519876|large uterusnull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|Neoplasm of uncertain or unknown behavior of uterus|Disorder|false|false|C4266525;C0042149;C1519876|uterus
null|Uterine Diseases|Disorder|false|false|C4266525;C0042149;C1519876|uterusnull|examination of uterus|Procedure|false|false|C4266525;C0042149;C1519876|uterusnull|Pelvis>Uterus|Anatomy|false|false|C0151994;C0869889;C0042131;C0496919;C0029936;C0278321|uterus
null|Mouse Uterus|Anatomy|false|false|C0151994;C0869889;C0042131;C0496919;C0029936;C0278321|uterus
null|Uterus|Anatomy|false|false|C0151994;C0869889;C0042131;C0496919;C0029936;C0278321|uterusnull|Fibroid Tumor|Disorder|false|false||fibroidnull|Pelvic lymph node group|Anatomy|false|false|C0015252;C0728940;C0024202|pelvic lymph nodenull|Pelvis|Anatomy|false|false|C0015252;C0728940;C0024202|pelvicnull|lymph nodes|Anatomy|false|false|C0024202;C0015252;C0728940|lymph nodenull|Lymph|Finding|false|false|C0024204;C0030797;C0729595|lymphnull|removal technique|Procedure|false|false|C0729595;C0024204;C0030797|resection
null|Excision|Procedure|false|false|C0729595;C0024204;C0030797|resectionnull|Complete cystectomy|Procedure|false|false||radical cystectomynull|Radicals (chemistry)|Drug|false|false||radicalnull|Radical (qualifier value)|Modifier|false|false||radicalnull|Cystectomy|Procedure|false|false||cystectomynull|Adenohypophyseal Diseases|Disorder|false|false||anteriornull|Anterior|Modifier|false|false||anteriornull|Vaginectomy|Procedure|false|false||vaginectomynull|Vaginal Dosage Form|Drug|false|false|C0042232|vaginalnull|Vaginal Route of Administration|Finding|false|false|C0042232|vaginal
null|Vaginal (intended site)|Finding|false|false|C0042232|vaginalnull|Vagina|Anatomy|false|false|C4521343;C1522570;C1272941|vaginalnull|Vaginal|Modifier|false|false||vaginalnull|Optical Image Reconstruction|Procedure|false|false||reconstruction
null|Reconstructive Surgical Procedures|Procedure|false|false||reconstructionnull|Structure of ileal conduit|Disorder|false|false|C0020885|ileal conduitnull|Ileal conduit procedure|Procedure|false|false|C0020885|ileal conduitnull|ileum|Anatomy|false|false|C0348002;C0441253|ilealnull|Conduit implant|Device|false|false||conduitnull|Surgical construction|Procedure|false|false||creationnull|Creation|Event|false|false||creationnull|Course|Time|false|false||coursenull|Bacteremia|Finding|false|false||bacteremianull|Growth and Development function|Finding|false|false||development
null|development aspects|Finding|false|false||development
null|biological development|Finding|false|false||development
null|Development|Finding|false|false||developmentnull|Intraabdominal Route of Administration|Finding|false|false||intra-abdominalnull|Intra-abdominal|Modifier|false|false||intra-abdominalnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Collection Object - UML Entity|Finding|false|false||collection
null|Item Collection|Finding|false|false||collection
null|Collections (publication)|Finding|false|false||collection
null|Collection (action)|Finding|false|false||collectionnull|Drain placement|Procedure|false|false||drain placementnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|null|Procedure|false|false||placement
null|Implantation procedure|Procedure|false|false||placement
null|Clinical act of insertion|Procedure|false|false||placementnull|Placement|Modifier|false|false||placementnull|Deep thrombophlebitis|Disorder|false|false|C5239664|DVT
null|Deep Vein Thrombosis|Disorder|false|false|C5239664|DVTnull|area DVT|Anatomy|false|false|C2926618;C0149871;C0151950|DVTnull|null|Attribute|false|false|C5239664|DVTnull|Decreased Coagulation Activity [PE]|Finding|true|false||anticoagulation
null|Anticoagulation function|Finding|true|false||anticoagulation
null|ANTICOAGULATION (finding)|Finding|true|false||anticoagulationnull|Anticoagulation Therapy|Procedure|true|false||anticoagulationnull|Negative|Finding|false|false||Negative fornull|Rh Negative Blood Group|Finding|false|false||Negative
null|Negative|Finding|false|false||Negative
null|Negative Finding|Finding|false|false||Negativenull|Expression Negative|Lab|false|false||Negativenull|Negative - qualifier|Modifier|false|false||Negative
null|Negative Charge|Modifier|false|false||Negativenull|Negative Number|LabModifier|false|false||Negativenull|Malignant neoplasm of urinary bladder|Disorder|false|false|C0005682|bladder CAnull|Neoplasm of uncertain or unknown behavior of bladder|Disorder|false|false|C0005682|bladder
null|Benign neoplasm of bladder|Disorder|false|false|C0005682|bladder
null|Carcinoma in situ of bladder|Disorder|false|false|C0005682|bladdernull|Procedures on bladder|Procedure|false|false|C0005682|bladdernull|Urinary Bladder|Anatomy|false|false|C0496930;C0154017;C0154091;C0005684;C0872388|bladdernull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|C1orf210 gene|Finding|false|false||Tempnull|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Procedure|false|false||Tempnull|Temperature|LabModifier|false|false||Tempnull|delivery (history)|Finding|false|false||delivery
null|Transfer Technique|Finding|false|false||delivery
null|null|Finding|false|false||deliverynull|Obstetric Delivery|Procedure|false|false||deliverynull|null|Finding|false|false||Dyspnea
null|Dyspnea|Finding|false|false||Dyspneanull|Richmond Agitation-Sedation Scale Clinical Classification|Finding|false|false||RASSnull|Pain score|Finding|false|false||Pain Scorenull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Score|Finding|false|false||Scorenull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GENERALnull|General medical service|Procedure|false|false||GENERALnull|Generalized|Modifier|false|false||GENERALnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|apparent|Finding|false|false||apparentnull|Emotional distress|Finding|true|false||distress
null|Distress|Finding|true|false||distressnull|Face|Anatomy|false|false|C0231530|facialnull|Facial|Modifier|false|false||facialnull|Muscle twitch|Finding|false|false|C0015450|twitchesnull|Eye|Anatomy|false|false|C5848506|EYESnull|null|Attribute|false|false|C0015392|EYESnull|Anicteric|Finding|false|false||Anictericnull|Pupil|Anatomy|false|false||pupilsnull|Round shape|Modifier|false|false||roundnull|ENT problem|Finding|false|false|C0150934;C0175196|ENT
null|NT5E gene|Finding|false|false|C0150934;C0175196|ENT
null|NT5E wt Allele|Finding|false|false|C0150934;C0175196|ENTnull|Structure of entorhinal cortex|Anatomy|false|false|C0262471;C3889152;C1417861|ENT
null|Ear, nose and throat|Anatomy|false|false|C0262471;C3889152;C1417861|ENTnull|Otolaryngology specialty|Title|false|false||ENTnull|EPRS1 gene|Finding|false|false|C0013443;C0521421|Earsnull|null|Anatomy|false|false|C0041834;C1414437|Ears
null|Ear structure|Anatomy|false|false|C0041834;C1414437|Earsnull|Visible|Modifier|false|false||visiblenull|Erythema|Disorder|false|false|C0013443;C0521421|erythemanull|Physical trauma|Disorder|true|false||trauma
null|Traumatic injury|Disorder|true|false||trauma
null|Trauma|Disorder|true|false||traumanull|Trauma assessment and care|Procedure|true|false||traumanull|Trauma, nursing specialty|Title|false|false||traumanull|trauma qualifier|Modifier|false|false||traumanull|Oropharyngeal|Anatomy|false|false|C0015388;C1546629;C0041834;C0221198;C1546698;C0221198|Oropharynxnull|Lesion|Finding|true|false|C0521367|visible lesionnull|Visible|Modifier|false|false||visiblenull|Lesion|Finding|true|false|C0521367|lesion
null|null|Finding|true|false|C0521367|lesionnull|Erythema|Disorder|true|false|C0521367|erythemanull|null|Finding|false|false|C0521367|exudate
null|Exudate|Finding|false|false|C0521367|exudatenull|Heart regular|Finding|false|false|C4037974;C0018787|Heart regularnull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|Heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|Heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|Heartnull|Chest>Heart|Anatomy|false|false|C0425586;C0153957;C0153500;C0018808;C0795691|Heart
null|Heart|Anatomy|false|false|C0425586;C0153957;C0153500;C0018808;C0795691|Heartnull|Regular|Modifier|false|false||regularnull|Heart murmur|Finding|true|false|C4037974;C0018787|murmurnull|Jugular venous engorgement|Finding|true|false||JVDnull|Respiratory, thoracic and mediastinal disorders|Disorder|false|false||RESPnull|Respiratory rate|Attribute|false|false||RESPnull|Lung|Anatomy|false|false|C1550016|Lungsnull|Remote control command - Clear|Finding|false|false|C0024109|clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Auscultation|Procedure|false|false||auscultationnull|Language Ability Proficiency - Good|Finding|false|false||good
null|Language Proficiency - Good|Finding|false|false||goodnull|Specimen Quality - Good|Modifier|false|false||good
null|Good|Modifier|false|false||goodnull|Air Movements|Phenomenon|false|false||air movementnull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false||air
null|AIRN gene|Finding|false|false||air
null|AI/RHEUM|Finding|false|false||airnull|Movement|Finding|false|false||movementnull|outcomes otolaryngology breathing|Finding|false|false||Breathing
null|Inspiration (function)|Finding|false|false||Breathing
null|Respiration|Finding|false|false||Breathingnull|null|Attribute|false|false||Breathingnull|respiratory system process|Phenomenon|false|false||Breathingnull|Abdomen soft|Finding|false|false|C0230168;C0000726|Abdomen softnull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|Abdomennull|Abdomen problem|Finding|false|false|C0230168;C0000726|Abdomennull|Abdomen|Anatomy|false|false|C0153662;C0426663;C0941288|Abdomen
null|Abdominal Cavity|Anatomy|false|false|C0153662;C0426663;C0941288|Abdomennull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|Palpation|Procedure|false|false||palpationnull|Intestines|Anatomy|false|false||Bowelnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|LRRC4B gene|Finding|true|false||HSMnull|Suprapubic|Anatomy|false|false||suprapubicnull|suprapubic approach|Modifier|false|false||suprapubicnull|Fullness|Modifier|false|false||fullnessnull|Emotional tenderness|Finding|true|false||tenderness
null|Sore to touch|Finding|true|false||tendernessnull|Palpation|Procedure|false|false||palpationnull|null|Finding|false|false||catheternull|catheter device|Device|false|false||catheter
null|XXX>Catheter|Device|false|false||catheternull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Medullary sponge kidney|Disorder|false|false||MSK
null|Medullary sponge kidney|Disorder|false|false||MSKnull|SIK1 gene|Finding|false|false||MSKnull|Supple neck|Finding|false|false|C0027530;C3159206|Neck supplenull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|Neck
null|Neck problem|Finding|false|false|C0027530;C3159206|Necknull|dendritic spine neck|Anatomy|false|false|C2230237;C0812434;C0684335|Neck
null|Neck|Anatomy|false|false|C2230237;C0812434;C0684335|Necknull|Supple|Finding|false|false||supplenull|All extremities|Anatomy|false|false|C0808080|all extremitiesnull|All extremities|Anatomy|false|false|C0808080|extremities
null|Limb structure|Anatomy|false|false|C0808080|extremitiesnull|Strength (attribute)|Finding|false|false|C0278454;C0278454;C0015385|strengthnull|Pharmaceutical Strength|LabModifier|false|false||strength
null|Physical Strength|LabModifier|false|false||strengthnull|Full|Modifier|false|false||fullnull|Symmetric Relationship|Finding|false|false|C0015385;C3687203|symmetric
null|Symmetrical|Finding|false|false|C0015385;C3687203|symmetricnull|All limbs|Anatomy|false|false|C0332516;C2699744|all limbsnull|Limb structure|Anatomy|false|false|C0332516;C2699744|limbsnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765|SKIN
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765|SKINnull|Skin Specimen Source Code|Finding|false|false|C1123023;C4520765|SKIN
null|Skin Specimen|Finding|false|false|C1123023;C4520765|SKINnull|Skin, Human|Anatomy|false|false|C1546781;C0444099;C0178298;C0496955|SKIN
null|Skin|Anatomy|false|false|C1546781;C0444099;C0178298;C0496955|SKINnull|Skin rash|Finding|true|false||rashes
null|Exanthema|Finding|true|false||rashesnull|Ulcer|Finding|true|false||ulcerationsnull|Neurology speciality|Title|false|false||NEUROnull|Neurologic (qualifier value)|Modifier|false|false||NEUROnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|FANCONI ANEMIA, COMPLEMENTATION GROUP E|Disorder|false|false|C0015450;C4266571|facenull|FANCE wt Allele|Finding|false|false|C0015450;C4266571|face
null|FANCE gene|Finding|false|false|C0015450;C4266571|face
null|ELOVL6 gene|Finding|false|false|C0015450;C4266571|facenull|Head>Face|Anatomy|false|false|C3160739;C0332516;C2699744;C1423759;C2828055;C1414531|face
null|Face|Anatomy|false|false|C3160739;C0332516;C2699744;C1423759;C2828055;C1414531|facenull|Face (spatial concept)|Modifier|false|false||facenull|Symmetric Relationship|Finding|false|false|C0015450;C4266571|symmetric
null|Symmetrical|Finding|false|false|C0015450;C4266571|symmetricnull|Gaze|Finding|false|false||gazenull|Immunostimulating conjugate (antigen)|Drug|false|false||conjugatenull|Speech|Finding|false|false||speechnull|Speech assessment|Procedure|false|false||speechnull|All limbs|Anatomy|false|false|C2229507;C0152054;C0036658;C0542538;C3842678;C1306462;C1420817;C4521367;C0702221;C2350522;C0031765|all limbsnull|Limb structure|Anatomy|false|false|C0152054;C3842678;C1306462;C1420817;C4521367;C0031765;C0036658;C0542538;C0702221;C2350522;C2229507|limbsnull|Observation of Sensation|Finding|false|false|C3687203;C0015385|sensation
null|Sensory perception|Finding|false|false|C3687203;C0015385|sensationnull|sensory exam|Procedure|false|false|C3687203;C0015385|sensationnull|Sensation quality|Modifier|false|false||sensationnull|Light touch|Finding|false|false||light touchnull|TNFSF14 protein, human|Drug|false|false||light
null|TNFSF14 protein, human|Drug|false|false||lightnull|Light - subjective measurement|Finding|false|false|C0015385;C3687203|light
null|TNFSF14 wt Allele|Finding|false|false|C0015385;C3687203|light
null|TNFSF14 gene|Finding|false|false|C0015385;C3687203|light
null|Light color|Finding|false|false|C0015385;C3687203|lightnull|Phototherapy|Procedure|false|false|C0015385;C3687203|lightnull|Light|Phenomenon|false|false||lightnull|Light (qualifier)|Modifier|false|false||lightnull|Touch sensation|Finding|false|false|C3687203;C0015385|touch
null|Touch Perception|Finding|false|false|C3687203;C0015385|touchnull|Therapeutic Touch|Procedure|false|false|C0015385;C3687203|touchnull|Tactile|Modifier|false|false||touchnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Psychiatric problem|Disorder|false|false||PSYCH
null|Mental disorders|Disorder|false|false||PSYCHnull|Pleasant|Finding|false|false||pleasantnull|Appropriate affect|Disorder|false|false||appropriate affectnull|Appropriate|Modifier|false|false||appropriatenull|Affect (mental function)|Finding|false|false||affectnull|assessment of affect|Procedure|false|false||affectnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Urostomy bag|Device|false|false||Urostomy bagnull|Urostomy procedure|Procedure|false|false|C0559495|Urostomynull|Urological stoma|Anatomy|false|false|C1704765;C1552710;C0856443|Urostomynull|Bag Data Type|Finding|false|false|C0559495|bagnull|null|Device|false|false||bagnull|Bag (unit of presentation)|LabModifier|false|false||bag
null|Bag Dosing Unit|LabModifier|false|false||bagnull|Place - dosing instruction imperative|Finding|false|false|C0559495|placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Surrounding (qualifier value)|Modifier|false|false||surroundnull|Erythema|Disorder|true|false||erythemanull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Laboratory Results|Lab|false|false||LABORATORY RESULTSnull|Diagnostic Service Section ID - Laboratory|Finding|false|false||LABORATORY
null|Laboratory domain|Finding|false|false||LABORATORY
null|Referral type - Laboratory|Finding|false|false||LABORATORYnull|null|Attribute|false|false||LABORATORYnull|Laboratory|Device|false|false||LABORATORYnull|Laboratory observation|Lab|false|false||LABORATORYnull|Laboratory|Entity|false|false||LABORATORYnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0851353;C0005768;C0229664;C0005767|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C0014792;C1114281|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0005768;C0229664;C0005767;C0851353|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C0014792;C1114281|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0005768;C0229664;C0005767;C0851353|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Microbiology Diagnostic Service Section ID|Finding|false|false||MICROBIOLOGY
null|Microbiological|Finding|false|false||MICROBIOLOGY
null|Microbiology - Laboratory Class|Finding|false|false||MICROBIOLOGYnull|Microbiology procedure|Procedure|false|false||MICROBIOLOGYnull|Science of Microbiology|Title|false|false||MICROBIOLOGYnull|Portion of urine|Finding|false|false|C1515974|URINE
null|null|Finding|false|false|C1515974|URINE
null|Urine|Finding|false|false|C1515974|URINE
null|In Urine|Finding|false|false|C1515974|URINE
null|Urine specimen|Finding|false|false|C1515974|URINEnull|null|Finding|false|false|C1515974|Sitenull|Anatomic Site|Anatomy|false|false|C1546778;C0042036;C2963137;C0042037;C1547942;C1610733|Sitenull|Study Site|Modifier|false|false||Site
null|Site|Modifier|false|false||Sitenull|Cystoscopy|Procedure|false|false|C0227613;C0227665;C0022646|CYSTOSCOPYnull|Right kidney|Anatomy|false|false|C0812426;C1552823;C0496927;C0496892;C0010702;C4554465;C0869841|RIGHT KIDNEYnull|Table Cell Horizontal Align - right|Finding|false|false|C0227613|RIGHTnull|Right sided|Modifier|false|false||RIGHT
null|Right|Modifier|false|false||RIGHTnull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false|C0227613;C0227665;C0022646|KIDNEY
null|Benign neoplasm of kidney|Disorder|false|false|C0227613;C0227665;C0022646|KIDNEYnull|Kidney problem|Finding|false|false|C0227613;C0227665;C0022646|KIDNEYnull|examination of kidney|Procedure|false|false|C0227665;C0022646;C0227613|KIDNEY
null|Procedures on Kidney|Procedure|false|false|C0227665;C0022646;C0227613|KIDNEYnull|Kidney|Anatomy|false|false|C4554465;C0869841;C0010702;C0812426;C0496927;C0496892|KIDNEY
null|Both kidneys|Anatomy|false|false|C4554465;C0869841;C0010702;C0812426;C0496927;C0496892|KIDNEYnull|Wash Dosage Form|Drug|false|false||WASHnull|Wash - dosing instruction imperative|Finding|false|false||WASH
null|Wash - Specimen Source Codes|Finding|false|false||WASH
null|WASHC1 gene|Finding|false|false||WASH
null|Wash - Administration Method|Finding|false|false||WASHnull|Cell Wash|Procedure|false|false||WASHnull|Wash (cleansing action)|Event|false|false||WASHnull|Final report|Finding|false|false||FINAL REPORTnull|Diagnosis Type - Final|Finding|false|false||FINALnull|Final|Time|false|false||FINALnull|End-stage|Modifier|false|false||FINALnull|Report (document)|Finding|false|false||REPORTnull|Reporting|Procedure|false|false||REPORTnull|null|Attribute|false|false||REPORTnull|Urine culture|Procedure|false|false||URINE CULTUREnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Enterococcus faecium|Entity|false|false||ENTEROCOCCUS FAECIUMnull|Enterococcus|Entity|false|false||ENTEROCOCCUSnull|cfu/mL|LabModifier|false|false||CFU/MLnull|Colony-forming unit|LabModifier|false|false||CFUnull|per milliliter|LabModifier|false|false||/MLnull|null|Event|false|false||REQUESTSnull|Microbial susceptibility tests|Procedure|false|false||SUSCEPTIBILITY TESTINGnull|Susceptibility (property) (qualifier value)|Finding|false|false||SUSCEPTIBILITYnull|Disease susceptibility|Attribute|false|false||SUSCEPTIBILITYnull|null|Subject|false|false||SUSCEPTIBILITYnull|Testing|Finding|false|false||TESTING
null|Tests (qualifier value)|Finding|false|false||TESTINGnull|Staphylococcus, coagulase negative (organism)|Entity|false|false||STAPHYLOCOCCUS, COAGULASE NEGATIVEnull|Unspecified Staphylococcus infection in conditions classified elsewhere and of unspecified site|Disorder|false|false||STAPHYLOCOCCUSnull|Genus staphylococcus|Entity|false|false||STAPHYLOCOCCUSnull|Coagulase|Drug|false|false||COAGULASE
null|Coagulase|Drug|false|false||COAGULASEnull|Rh Negative Blood Group|Finding|false|false||NEGATIVE
null|Negative|Finding|false|false||NEGATIVE
null|Negative Finding|Finding|false|false||NEGATIVEnull|Expression Negative|Lab|false|false||NEGATIVEnull|Negative - qualifier|Modifier|false|false||NEGATIVE
null|Negative Charge|Modifier|false|false||NEGATIVEnull|Negative Number|LabModifier|false|false||NEGATIVEnull|cfu/mL|LabModifier|false|false||CFU/MLnull|Colony-forming unit|LabModifier|false|false||CFUnull|per milliliter|LabModifier|false|false||/MLnull|Corynebacterium species|Entity|false|false||CORYNEBACTERIUM SPECIES
null|Corynebacterium|Entity|false|false||CORYNEBACTERIUM SPECIESnull|Corynebacterium|Entity|false|false||CORYNEBACTERIUMnull|Species - Nature of Abnormal Testing|Finding|false|false||SPECIES
null|Species|Finding|false|false||SPECIESnull|Diphtheroids|Entity|false|false||DIPHTHEROIDSnull|cfu/mL|LabModifier|false|false||CFU/MLnull|Colony-forming unit|LabModifier|false|false||CFUnull|per milliliter|LabModifier|false|false||/MLnull|Antimicrobial susceptibility|Finding|false|false||SENSITIVITIESnull|methyl isocyanate|Drug|false|false||MIC
null|methyl isocyanate|Drug|false|false||MICnull|Ductal Carcinoma In Situ with Microinvasion|Disorder|false|false||MICnull|cisplatin/ifosfamide/mitomycin protocol|Procedure|false|false||MIC
null|Minimum Inhibitory Concentration Test|Procedure|false|false||MICnull|Micmac language|Entity|false|false||MICnull|Microgram per Milliliter|LabModifier|false|false||MCG/MLnull|microgram|LabModifier|false|false||MCGnull|per milliliter|LabModifier|false|false||/MLnull|Enterococcus faecium|Entity|false|false||ENTEROCOCCUS FAECIUMnull|Enterococcus|Entity|false|false||ENTEROCOCCUSnull|ampicillin|Drug|false|false||AMPICILLIN
null|ampicillins|Drug|false|false||AMPICILLIN
null|ampicillins|Drug|false|false||AMPICILLIN
null|ampicillin|Drug|false|false||AMPICILLINnull|nitrofurantoin|Drug|false|false||NITROFURANTOIN
null|nitrofurantoin|Drug|false|false||NITROFURANTOINnull|Tetracycline Antibiotics|Drug|false|false||TETRACYCLINE
null|Tetracycline Antibiotics|Drug|false|false||TETRACYCLINE
null|tetracycline|Drug|false|false||TETRACYCLINE
null|tetracycline|Drug|false|false||TETRACYCLINEnull|Tetracyclines causing adverse effects in therapeutic use|Disorder|false|false||TETRACYCLINEnull|vancomycin|Drug|false|false||VANCOMYCIN
null|vancomycin|Drug|false|false||VANCOMYCINnull|Vancomycin measurement|Procedure|false|false||VANCOMYCINnull|Blood culture|Procedure|false|false||Blood culturesnull|Blood and lymphatic system disorders|Disorder|false|false||Bloodnull|peripheral blood|Finding|false|false||Blood
null|Blood|Finding|false|false||Blood
null|In Blood|Finding|false|false||Bloodnull|Culture (Anthropological)|Finding|false|false||culturesnull|Sepsis|Disorder|false|false||sepsis
null|Septicemia|Disorder|false|false||sepsisnull|Sepsis <Sepsidae>|Entity|false|false||sepsisnull|Urinary tract|Anatomy|false|false||urinary tract
null|Urinary system|Anatomy|false|false||urinary tractnull|Urinary tract|Anatomy|false|false||urinarynull|urinary|Modifier|false|false||urinarynull|Tract|Anatomy|false|false||tractnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|null|Device|false|false||stentnull|degree of relationship - exchange|Finding|false|false||exchangenull|Exchange (clinical)|Attribute|false|false||exchangenull|vancomycin|Drug|false|false||vancomycin
null|vancomycin|Drug|false|false||vancomycinnull|Vancomycin measurement|Procedure|false|false||vancomycinnull|cefepime|Drug|false|false||cefepime
null|cefepime|Drug|false|false||cefepimenull|ceftriaxone|Drug|false|false||ceftriaxone
null|ceftriaxone|Drug|false|false||ceftriaxonenull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|resistant - Observation Interpretation Susceptibility|Finding|false|false||resistant
null|Resistant (qualifier value)|Finding|false|false||resistantnull|Antimicrobial Resistance Result|Lab|false|false||resistantnull|Organism|Entity|false|false||organismsnull|Rapid|Modifier|false|false||rapidlynull|Portion of urine|Finding|false|false||urine
null|null|Finding|false|false||urine
null|Urine|Finding|false|false||urine
null|In Urine|Finding|false|false||urine
null|Urine specimen|Finding|false|false||urinenull|Sensitive|Finding|false|false||sensitive tonull|Sensitive|Finding|false|false||sensitivenull|stimulus sensitivity|Modifier|false|false||sensitivenull|ampicillin|Drug|false|false||ampicillin
null|ampicillins|Drug|false|false||ampicillin
null|ampicillins|Drug|false|false||ampicillin
null|ampicillin|Drug|false|false||ampicillinnull|Peripherally inserted central catheter (physical object)|Device|false|false||PICC linenull|Peripherally Inserted Central Catheter Line Insertion|Procedure|false|false||PICCnull|Peripherally inserted central catheter (physical object)|Device|false|false||PICCnull|Line Specimen|Drug|false|false||line
null|Long Interspersed Elements|Drug|false|false||line
null|Long Interspersed Elements|Drug|false|false||linenull|line source specimen code|Finding|false|false||linenull|Intravascular line|Device|false|false||linenull|Linear|Modifier|false|false||linenull|Line Unit of Length|LabModifier|false|false||linenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|Two weeks|Time|false|false||two weeksnull|week|Time|false|false||weeksnull|Total|Modifier|false|false||totalnull|ampicillin|Drug|false|false||ampicillin
null|ampicillins|Drug|false|false||ampicillin
null|ampicillins|Drug|false|false||ampicillin
null|ampicillin|Drug|false|false||ampicillinnull|Complicated|Finding|false|false||complicatednull|Urinary tract|Anatomy|false|false||urinarynull|urinary|Modifier|false|false||urinarynull|Tract|Anatomy|false|false|C3714514;C1561538;C1561539;C1524062;C4534574;C0009450|tractnull|Communicable Diseases|Disorder|false|false|C1185740|infectionnull|Infection|Finding|false|false|C1185740|infectionnull|Additional day|Finding|false|false|C1185740|additional daynull|Additional|Finding|false|false|C1185740|additionalnull|Transaction counts and value totals - day|Finding|false|false|C1185740|day
null|Precision - day|Finding|false|false|C1185740|daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|day|Time|false|false||daysnull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Drugs used in migraine prophylaxis|Drug|false|false||prophylacticnull|Prophylactic behavior|Finding|false|false||prophylacticnull|Condoms, Male|Device|false|false||prophylacticnull|epithelial membrane protein-1|Drug|false|false|C0149552|TMP
null|trimethoprim|Drug|false|false|C0149552|TMP
null|trimethoprim|Drug|false|false|C0149552|TMP
null|EMP1 protein, human|Drug|false|false|C0149552|TMP
null|Thymidine Monophosphate|Drug|false|false|C0149552|TMP
null|Thymidine Monophosphate|Drug|false|false|C0149552|TMPnull|AML Transfusion Medicine Procedures Table|Finding|false|false|C0149552|TMP
null|EMP1 protein, human|Finding|false|false|C0149552|TMP
null|epithelial membrane protein-1|Finding|false|false|C0149552|TMP
null|EMP1 wt Allele, Human|Finding|false|false|C0149552|TMP
null|EMP1 gene|Finding|false|false|C0149552|TMPnull|Structure of temporal pole|Anatomy|false|false|C0812384;C1259382;C1706000;C0384479;C5420102;C1259382;C0040079;C0384479;C0041041|TMPnull|ampicillin|Drug|false|false||ampicillin
null|ampicillins|Drug|false|false||ampicillin
null|ampicillins|Drug|false|false||ampicillin
null|ampicillin|Drug|false|false||ampicillinnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Course|Time|false|false||coursenull|ampicillin|Drug|false|false||ampicillin
null|ampicillins|Drug|false|false||ampicillin
null|ampicillins|Drug|false|false||ampicillin
null|ampicillin|Drug|false|false||ampicillinnull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|Additional|Finding|false|false||additionalnull|day|Time|false|false||daysnull|Restart|Modifier|false|false||restartnull|epithelial membrane protein-1|Drug|false|false|C0149552|TMP
null|trimethoprim|Drug|false|false|C0149552|TMP
null|trimethoprim|Drug|false|false|C0149552|TMP
null|EMP1 protein, human|Drug|false|false|C0149552|TMP
null|Thymidine Monophosphate|Drug|false|false|C0149552|TMP
null|Thymidine Monophosphate|Drug|false|false|C0149552|TMPnull|AML Transfusion Medicine Procedures Table|Finding|false|false|C0149552|TMP
null|EMP1 protein, human|Finding|false|false|C0149552|TMP
null|epithelial membrane protein-1|Finding|false|false|C0149552|TMP
null|EMP1 wt Allele, Human|Finding|false|false|C0149552|TMP
null|EMP1 gene|Finding|false|false|C0149552|TMPnull|Structure of temporal pole|Anatomy|false|false|C0812384;C1259382;C1706000;C0384479;C5420102;C1418850;C1259382;C0040079;C0384479;C0041041|TMPnull|Daily|Time|false|false||dailynull|PPP4C gene|Finding|false|false|C0149552|ppxnull|Antibiotics|Drug|false|false||antibioticnull|Course|Time|false|false||coursenull|Follow-up status|Finding|false|false||follow upnull|follow-up|Procedure|false|false||follow upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|Problems - What subject filter|Finding|false|false||problemsnull|Hospitalization|Procedure|false|false||hospitalizationnull|Initially|Time|false|false||initiallynull|Probable diagnosis|Finding|false|false|C1550297|likely
null|Probably|Finding|false|false|C1550297|likelynull|Prerenal|Anatomy|false|false|C0332148;C0750492|prerenalnull|Sepsis|Disorder|false|false||sepsis
null|Septicemia|Disorder|false|false||sepsisnull|Sepsis <Sepsidae>|Entity|false|false||sepsisnull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|Table Frame - above|Finding|false|false||abovenull|Upper|Modifier|false|false||abovenull|creatinine|Drug|false|false||creatinine
null|creatinine|Drug|false|false||creatininenull|Creatinine metabolic function|Finding|false|false||creatininenull|Creatinine measurement|Procedure|false|false||creatininenull|losartan|Drug|false|false||Losartan
null|losartan|Drug|false|false||Losartannull|Initially|Time|false|false||initiallynull|On discharge|Time|false|false||on dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Hyperlipidemia|Disorder|false|false||Hyperlipidemia
null|Hyperlipoproteinemias|Disorder|false|false||Hyperlipidemianull|Serum lipids high (finding)|Finding|false|false||Hyperlipidemianull|atorvastatin|Drug|false|false||atorvastatin
null|atorvastatin|Drug|false|false||atorvastatinnull|Daily|Time|false|false||dailynull|Hypothyroidism|Disorder|false|false||Hypothyroidismnull|Synthetic Levothyroxine|Drug|false|false||levothyroxine
null|Synthetic Levothyroxine|Drug|false|false||levothyroxine
null|levothyroxine|Drug|false|false||levothyroxine
null|levothyroxine|Drug|false|false||levothyroxine
null|levothyroxine|Drug|false|false||levothyroxinenull|microgram|LabModifier|false|false||mcgnull|Daily|Time|false|false||dailynull|per 30 minutes|Time|false|false||30 minutes
null|30 Minutes|Time|false|false||30 minutesnull|Minute of time|Time|false|false||minutesnull|Minute Unit of Plane Angle|LabModifier|false|false||minutes
null|Minute (diminutive)|LabModifier|false|false||minutes
null|Small|LabModifier|false|false||minutesnull|On discharge|Time|false|false||on dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|activities (history)|Finding|false|false||activitiesnull|Activities|Event|false|false||activitiesnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Accurate (qualifier value)|Modifier|false|false||accuratenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Mild Severity of Illness Code|Finding|false|false||Mildnull|Mild (qualifier value)|Modifier|false|false||Mild
null|Mild Allergy Severity|Modifier|false|false||Mildnull|Fever symptoms (finding)|Finding|false|false||Fever
null|Fever|Finding|false|false||Fevernull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|Cyanocobalamin Drug Class|Drug|false|false||Cyanocobalamin
null|Cyanocobalamin Drug Class|Drug|false|false||Cyanocobalamin
null|vitamin B12|Drug|false|false||Cyanocobalamin
null|vitamin B12|Drug|false|false||Cyanocobalamin
null|vitamin B12|Drug|false|false||Cyanocobalaminnull|microgram|LabModifier|false|false||mcgnull|Daily|Time|false|false||DAILYnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|levothyroxine sodium|Drug|false|false||Levothyroxine Sodium
null|levothyroxine sodium|Drug|false|false||Levothyroxine Sodium
null|levothyroxine sodium|Drug|false|false||Levothyroxine Sodiumnull|Synthetic Levothyroxine|Drug|false|false||Levothyroxine
null|Synthetic Levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxinenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|microgram|LabModifier|false|false||mcgnull|Daily|Time|false|false||DAILYnull|lorazepam|Drug|false|false||LORazepam
null|lorazepam|Drug|false|false||LORazepamnull|Every twelve hours|Time|false|false||Q12Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Anxiety Disorders|Disorder|false|false||anxiety
null|Anxiety|Disorder|false|false||anxietynull|Anxiety symptoms|Finding|false|false||anxietynull|losartan potassium|Drug|false|false||Losartan Potassium
null|losartan potassium|Drug|false|false||Losartan Potassiumnull|losartan|Drug|false|false||Losartan
null|losartan|Drug|false|false||Losartannull|Potassium Drug Class|Drug|false|false||Potassium
null|Dietary Potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassiumnull|Potassium metabolic function|Finding|false|false||Potassiumnull|Potassium measurement|Procedure|false|false||Potassiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitaminsnull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|Daily|Time|false|false||DAILYnull|polyethylene glycols|Drug|false|false||Polyethylene Glycol
null|polyethylene glycols|Drug|false|false||Polyethylene Glycolnull|high-density polyethylene|Drug|false|false||Polyethylene
null|high-density polyethylene|Drug|false|false||Polyethylene
null|polyethylenes|Drug|false|false||Polyethylene
null|polyethylenes|Drug|false|false||Polyethylene
null|Polyethylene|Drug|false|false||Polyethylene
null|Polyethylene|Drug|false|false||Polyethylenenull|ethylene glycol|Drug|false|false||Glycol
null|Glycol|Drug|false|false||Glycol
null|ethylene glycol|Drug|false|false||Glycol
null|Glycols|Drug|false|false||Glycolnull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Constipation|Finding|false|false||Constipationnull|Firstly|Modifier|false|false||Firstnull|First (number)|LabModifier|false|false||Firstnull|Line Specimen|Drug|false|false||Line
null|Long Interspersed Elements|Drug|false|false||Line
null|Long Interspersed Elements|Drug|false|false||Linenull|line source specimen code|Finding|false|false||Linenull|Intravascular line|Device|false|false||Linenull|Linear|Modifier|false|false||Linenull|Line Unit of Length|LabModifier|false|false||Linenull|trimethoprim|Drug|false|false||Trimethoprim
null|trimethoprim|Drug|false|false||Trimethoprimnull|Every twenty four hours|Time|false|false||Q24Hnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|ampicillin|Drug|false|false||Ampicillin
null|ampicillins|Drug|false|false||Ampicillin
null|ampicillins|Drug|false|false||Ampicillin
null|ampicillin|Drug|false|false||Ampicillinnull|Every eight hours|Time|false|false||Q8Hnull|ampicillin sodium|Drug|false|false||ampicillin sodium
null|ampicillin sodium|Drug|false|false||ampicillin sodiumnull|ampicillin|Drug|false|false||ampicillin
null|ampicillins|Drug|false|false||ampicillin
null|ampicillins|Drug|false|false||ampicillin
null|ampicillin|Drug|false|false||ampicillinnull|Sodium supplements|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|Sodium Drug Class|Drug|false|false||sodiumnull|Sodium metabolic function|Finding|false|false||sodiumnull|Sodium measurement|Procedure|false|false||sodiumnull|Every eight hours|Time|false|false||Every eight hoursnull|Every - dosing instruction fragment|Finding|false|false||Everynull|Every (qualifier)|Modifier|false|false||Everynull|Hour|Time|false|false||hoursnull|PRSS30P gene|Finding|false|false||Dispnull|Dispense (activity)|Event|false|false||Dispnull|Vial device|Device|false|false||Vialnull|Vial (unit of presentation)|LabModifier|false|false||Vial
null|Vial Dosing Unit|LabModifier|false|false||Vialnull|refill|Finding|false|false||Refillsnull|ampicillin sodium|Drug|false|false||ampicillin sodium
null|ampicillin sodium|Drug|false|false||ampicillin sodiumnull|ampicillin|Drug|false|false||ampicillin
null|ampicillins|Drug|false|false||ampicillin
null|ampicillins|Drug|false|false||ampicillin
null|ampicillin|Drug|false|false||ampicillinnull|Sodium supplements|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|Sodium Drug Class|Drug|false|false||sodiumnull|Sodium metabolic function|Finding|false|false||sodiumnull|Sodium measurement|Procedure|false|false||sodiumnull|Every eight hours|Time|false|false||Every eight hoursnull|Every - dosing instruction fragment|Finding|false|false||Everynull|Every (qualifier)|Modifier|false|false||Everynull|Hour|Time|false|false||hoursnull|PRSS30P gene|Finding|false|false||Dispnull|Dispense (activity)|Event|false|false||Dispnull|Vial device|Device|false|false||Vialnull|Vial (unit of presentation)|LabModifier|false|false||Vial
null|Vial Dosing Unit|LabModifier|false|false||Vialnull|refill|Finding|false|false||Refillsnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Mild Severity of Illness Code|Finding|false|false||Mildnull|Mild (qualifier value)|Modifier|false|false||Mild
null|Mild Allergy Severity|Modifier|false|false||Mildnull|Fever symptoms (finding)|Finding|false|false||Fever
null|Fever|Finding|false|false||Fevernull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|Cyanocobalamin Drug Class|Drug|false|false||Cyanocobalamin
null|Cyanocobalamin Drug Class|Drug|false|false||Cyanocobalamin
null|vitamin B12|Drug|false|false||Cyanocobalamin
null|vitamin B12|Drug|false|false||Cyanocobalamin
null|vitamin B12|Drug|false|false||Cyanocobalaminnull|microgram|LabModifier|false|false||mcgnull|Daily|Time|false|false||DAILYnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|levothyroxine sodium|Drug|false|false||Levothyroxine Sodium
null|levothyroxine sodium|Drug|false|false||Levothyroxine Sodium
null|levothyroxine sodium|Drug|false|false||Levothyroxine Sodiumnull|Synthetic Levothyroxine|Drug|false|false||Levothyroxine
null|Synthetic Levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxinenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|microgram|LabModifier|false|false||mcgnull|Daily|Time|false|false||DAILYnull|lorazepam|Drug|false|false||LORazepam
null|lorazepam|Drug|false|false||LORazepamnull|Every twelve hours|Time|false|false||Q12Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Anxiety Disorders|Disorder|false|false||anxiety
null|Anxiety|Disorder|false|false||anxietynull|Anxiety symptoms|Finding|false|false||anxietynull|losartan potassium|Drug|false|false||Losartan Potassium
null|losartan potassium|Drug|false|false||Losartan Potassiumnull|losartan|Drug|false|false||Losartan
null|losartan|Drug|false|false||Losartannull|Potassium Drug Class|Drug|false|false||Potassium
null|Dietary Potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassiumnull|Potassium metabolic function|Finding|false|false||Potassiumnull|Potassium measurement|Procedure|false|false||Potassiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitaminsnull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|Daily|Time|false|false||DAILYnull|polyethylene glycols|Drug|false|false||Polyethylene Glycol
null|polyethylene glycols|Drug|false|false||Polyethylene Glycolnull|high-density polyethylene|Drug|false|false||Polyethylene
null|high-density polyethylene|Drug|false|false||Polyethylene
null|polyethylenes|Drug|false|false||Polyethylene
null|polyethylenes|Drug|false|false||Polyethylene
null|Polyethylene|Drug|false|false||Polyethylene
null|Polyethylene|Drug|false|false||Polyethylenenull|ethylene glycol|Drug|false|false||Glycol
null|Glycol|Drug|false|false||Glycol
null|ethylene glycol|Drug|false|false||Glycol
null|Glycols|Drug|false|false||Glycolnull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Constipation|Finding|false|false||Constipationnull|Firstly|Modifier|false|false||Firstnull|First (number)|LabModifier|false|false||Firstnull|Line Specimen|Drug|false|false||Line
null|Long Interspersed Elements|Drug|false|false||Line
null|Long Interspersed Elements|Drug|false|false||Linenull|line source specimen code|Finding|false|false||Linenull|Intravascular line|Device|false|false||Linenull|Linear|Modifier|false|false||Linenull|Line Unit of Length|LabModifier|false|false||Linenull|ARID1A protein, human|Drug|false|false||HELD
null|ARID1A protein, human|Drug|false|false||HELDnull|Held - activity status|Finding|false|false||HELD
null|ARID1A wt Allele|Finding|false|false||HELDnull|trimethoprim|Drug|false|false||Trimethoprim
null|trimethoprim|Drug|false|false||Trimethoprimnull|Every twenty four hours|Time|false|false||Q24Hnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|trimethoprim|Drug|false|false||Trimethoprim
null|trimethoprim|Drug|false|false||Trimethoprimnull|ampicillin|Drug|false|false||ampicillin
null|ampicillins|Drug|false|false||ampicillin
null|ampicillins|Drug|false|false||ampicillin
null|ampicillin|Drug|false|false||ampicillinnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|long-term care|Procedure|false|false||Extended Carenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Complicated|Finding|false|false||Complicatednull|urinastatin|Drug|false|false||UTI
null|urinastatin|Drug|false|false||UTInull|Urinary tract infection|Disorder|false|false||UTInull|AMBP wt Allele|Finding|false|false||UTI
null|AMBP gene|Finding|false|false||UTInull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Fever|Finding|false|false||feversnull|Chills|Finding|false|false||chillsnull|Fever|Finding|false|false||feversnull|Chills|Finding|false|false||chillsnull|null|Device|false|false||stentnull|degree of relationship - exchange|Finding|false|false||exchangenull|Exchange (clinical)|Attribute|false|false||exchangenull|Portion of urine|Finding|false|false||urine
null|null|Finding|false|false||urine
null|Urine|Finding|false|false||urine
null|In Urine|Finding|false|false||urine
null|Urine specimen|Finding|false|false||urinenull|Enterococcus|Entity|false|false||enterococcus speciesnull|Enterococcus|Entity|false|false||enterococcusnull|Species - Nature of Abnormal Testing|Finding|false|false||species
null|Species|Finding|false|false||speciesnull|Source (property) (qualifier value)|Finding|false|false||source
null|Term Source|Finding|false|false||source
null|Source|Finding|false|false||sourcenull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Enterococcus|Entity|false|false||enterococcusnull|Peripherally inserted central catheter (physical object)|Device|false|false||PICC linenull|Peripherally Inserted Central Catheter Line Insertion|Procedure|false|false||PICCnull|Peripherally inserted central catheter (physical object)|Device|false|false||PICCnull|Line Specimen|Drug|false|false||line
null|Long Interspersed Elements|Drug|false|false||line
null|Long Interspersed Elements|Drug|false|false||linenull|line source specimen code|Finding|false|false||linenull|Intravascular line|Device|false|false||linenull|Linear|Modifier|false|false||linenull|Line Unit of Length|LabModifier|false|false||linenull|Total|Modifier|false|false||totalnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Course|Time|false|false||coursenull|ampicillin|Drug|false|false||ampicillin
null|ampicillins|Drug|false|false||ampicillin
null|ampicillins|Drug|false|false||ampicillin
null|ampicillin|Drug|false|false||ampicillinnull|Injury of kidney|Disorder|false|false|C0227665;C0022646|kidney injurynull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false|C0227665;C0022646|kidney
null|Benign neoplasm of kidney|Disorder|false|false|C0227665;C0022646|kidneynull|Kidney problem|Finding|false|false|C0227665;C0022646|kidneynull|examination of kidney|Procedure|false|false|C0227665;C0022646|kidney
null|Procedures on Kidney|Procedure|false|false|C0227665;C0022646|kidneynull|Kidney|Anatomy|false|false|C4554465;C0869841;C0812426;C0496927;C0496892;C0160420|kidney
null|Both kidneys|Anatomy|false|false|C4554465;C0869841;C0812426;C0496927;C0496892;C0160420|kidneynull|Traumatic AND/OR non-traumatic injury|Disorder|false|false||injury
null|Traumatic injury|Disorder|false|false||injurynull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|Production Class Code - Pleasure|Finding|false|false||pleasure
null|pleasurable emotion|Finding|false|false||pleasurenull|Pleasure - Animals raised for recreation|Entity|false|false||pleasurenull|care of - AddressPartType|Finding|false|false||care ofnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions