 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|43,52|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|43,52|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|43,57|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|77,86|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|77,86|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|77,91|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|133,136|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|144,151|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|144,151|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|153,161|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|164,173|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|164,173|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|164,173|false|false|false|C0020517|Hypersensitivity|Allergies
Drug|Antibiotic|SIMPLE_SEGMENT|176,185|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|meropenem
Drug|Clinical Drug|SIMPLE_SEGMENT|176,185|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|meropenem
Drug|Organic Chemical|SIMPLE_SEGMENT|176,185|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|meropenem
Event|Event|SIMPLE_SEGMENT|176,185|false|false|false|||meropenem
Event|Event|SIMPLE_SEGMENT|188,197|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|188,197|false|false|false|C1999232|Attending (action)|Attending
Attribute|Clinical Attribute|SIMPLE_SEGMENT|209,218|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|209,218|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|209,218|false|false|false|C5441521|Complaint (finding)|Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|232,243|false|false|false|C0231832|Respiratory rate|Respiratory
Finding|Body Substance|SIMPLE_SEGMENT|232,243|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|Respiratory
Finding|Functional Concept|SIMPLE_SEGMENT|232,243|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|Respiratory
Finding|Intellectual Product|SIMPLE_SEGMENT|232,243|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|Respiratory
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|232,251|false|false|false|C1145670|Respiratory Failure|Respiratory Failure
Event|Event|SIMPLE_SEGMENT|244,251|false|false|false|||Failure
Finding|Functional Concept|SIMPLE_SEGMENT|244,251|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|Failure
Finding|Idea or Concept|SIMPLE_SEGMENT|244,251|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|Failure
Finding|Individual Behavior|SIMPLE_SEGMENT|244,251|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|Failure
Finding|Classification|SIMPLE_SEGMENT|254,259|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|260,268|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|260,268|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|272,290|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|281,290|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|281,290|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|281,290|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|281,290|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|281,290|false|false|false|C0184661|Interventional procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|292,302|false|false|false|C0443254|mechanical method|Mechanical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|292,302|false|false|false|C0699886|Mechanical Treatments|Mechanical
Event|Event|SIMPLE_SEGMENT|303,313|false|false|false|||Intubation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|303,313|false|false|false|C0021925|Intubation (procedure)|Intubation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|315,323|false|false|false|C0003842|Arteries|Arterial
Drug|Biologically Active Substance|SIMPLE_SEGMENT|325,329|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|325,329|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Drug|Substance|SIMPLE_SEGMENT|325,329|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Event|Event|SIMPLE_SEGMENT|325,329|false|false|false|||Line
Finding|Intellectual Product|SIMPLE_SEGMENT|325,329|false|false|false|C1546701|line source specimen code|Line
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|331,338|false|false|false|C0719205|Central brand of multivitamin with minerals|Central
Drug|Vitamin|SIMPLE_SEGMENT|331,338|false|false|false|C0719205|Central brand of multivitamin with minerals|Central
Event|Event|SIMPLE_SEGMENT|331,338|false|false|false|||Central
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|331,338|false|false|false|C1879652|Central Minus|Central
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|339,345|false|false|false|C0042449|Veins|Venous
Event|Event|SIMPLE_SEGMENT|346,352|false|false|false|||Access
Finding|Functional Concept|SIMPLE_SEGMENT|346,352|false|false|false|C1554204|Role Class - access|Access
Drug|Biologically Active Substance|SIMPLE_SEGMENT|354,358|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|354,358|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Drug|Substance|SIMPLE_SEGMENT|354,358|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Finding|Intellectual Product|SIMPLE_SEGMENT|354,358|false|false|false|C1546701|line source specimen code|Line
Event|Event|SIMPLE_SEGMENT|361,368|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|361,368|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|361,368|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|361,368|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|361,371|false|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|361,387|false|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|361,387|false|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|372,379|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|372,379|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|372,387|false|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|380,387|false|false|false|C0221423|Illness (finding)|Illness
Finding|Idea or Concept|SIMPLE_SEGMENT|404,408|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|SIMPLE_SEGMENT|404,408|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|SIMPLE_SEGMENT|413,418|false|false|false|||woman
Event|Event|SIMPLE_SEGMENT|429,441|false|false|false|||hospitalized
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|460,466|false|false|false|C0036690;C0243026|Sepsis;Septicemia|sepsis
Event|Event|SIMPLE_SEGMENT|460,466|false|false|false|||sepsis
Event|Event|SIMPLE_SEGMENT|471,476|false|false|false|||shock
Finding|Pathologic Function|SIMPLE_SEGMENT|471,476|false|false|false|C0036974|Shock|shock
Event|Event|SIMPLE_SEGMENT|478,489|false|false|false|||complicated
Event|Event|SIMPLE_SEGMENT|493,504|false|false|false|||readmission
Procedure|Health Care Activity|SIMPLE_SEGMENT|493,504|false|false|false|C4489276|Readmission|readmission
Event|Event|SIMPLE_SEGMENT|506,513|false|false|false|||hypoxia
Finding|Finding|SIMPLE_SEGMENT|506,513|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|hypoxia
Finding|Pathologic Function|SIMPLE_SEGMENT|506,513|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|hypoxia
Event|Event|SIMPLE_SEGMENT|514,525|false|false|false|||hypercarbia
Finding|Finding|SIMPLE_SEGMENT|514,525|false|false|false|C0020440|Hypercapnia|hypercarbia
Event|Event|SIMPLE_SEGMENT|536,544|false|false|false|||presents
Attribute|Clinical Attribute|SIMPLE_SEGMENT|550,561|false|false|false|C0231832|Respiratory rate|respiratory
Event|Event|SIMPLE_SEGMENT|550,561|false|false|false|||respiratory
Finding|Body Substance|SIMPLE_SEGMENT|550,561|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|SIMPLE_SEGMENT|550,561|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|SIMPLE_SEGMENT|550,561|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Event|Event|SIMPLE_SEGMENT|563,571|false|false|false|||distress
Finding|Finding|SIMPLE_SEGMENT|563,571|false|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|SIMPLE_SEGMENT|563,571|false|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Attribute|Clinical Attribute|SIMPLE_SEGMENT|576,587|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|SIMPLE_SEGMENT|576,587|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|SIMPLE_SEGMENT|576,587|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|SIMPLE_SEGMENT|576,587|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|576,595|false|false|false|C1145670|Respiratory Failure|respiratory failure
Event|Event|SIMPLE_SEGMENT|588,595|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|588,595|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|588,595|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|588,595|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Body Substance|SIMPLE_SEGMENT|603,610|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|603,610|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|603,610|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|637,641|false|false|false|||well
Finding|Finding|SIMPLE_SEGMENT|637,641|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|646,651|false|false|false|||rehab
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|646,651|false|false|false|C0034991|Rehabilitation therapy|rehab
Event|Event|SIMPLE_SEGMENT|678,683|false|false|false|||noted
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|704,713|false|false|false|C0344315|Depressed mood|depressed
Finding|Mental Process|SIMPLE_SEGMENT|715,721|false|false|false|C0229992|Psyche structure|mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|715,728|false|false|false|C0488568;C0488569||mental status
Finding|Finding|SIMPLE_SEGMENT|715,728|false|false|false|C0278060|Mental state|mental status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|722,728|false|false|false|C5889824||status
Event|Event|SIMPLE_SEGMENT|722,728|false|false|false|||status
Finding|Idea or Concept|SIMPLE_SEGMENT|722,728|false|false|false|C1546481|What subject filter - Status|status
Event|Event|SIMPLE_SEGMENT|731,740|false|false|false|||tachypnea
Finding|Finding|SIMPLE_SEGMENT|731,740|false|false|false|C0231835|Tachypnea|tachypnea
Event|Event|SIMPLE_SEGMENT|746,753|false|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|746,753|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|746,753|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|756,759|false|false|false|C0015063|Ethyl Methanesulfonate|EMS
Drug|Organic Chemical|SIMPLE_SEGMENT|756,759|false|false|false|C0015063|Ethyl Methanesulfonate|EMS
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|756,759|false|false|false|C0015063|Ethyl Methanesulfonate|EMS
Event|Event|SIMPLE_SEGMENT|756,759|false|false|false|||EMS
Finding|Gene or Genome|SIMPLE_SEGMENT|756,759|false|false|false|C5203240|EMSLR gene|EMS
Procedure|Health Care Activity|SIMPLE_SEGMENT|756,759|false|false|false|C0013961|Emergency Medical Services|EMS
Event|Event|SIMPLE_SEGMENT|764,770|false|false|false|||called
Event|Event|SIMPLE_SEGMENT|775,780|false|false|false|||found
Finding|Body Substance|SIMPLE_SEGMENT|785,792|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|785,792|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|785,792|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|798,806|true|false|false|||extremis
Event|Event|SIMPLE_SEGMENT|808,818|true|false|false|||intubation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|808,818|true|false|false|C0021925|Intubation (procedure)|intubation
Event|Event|SIMPLE_SEGMENT|823,832|true|false|false|||attempted
Event|Event|SIMPLE_SEGMENT|840,846|false|false|false|||failed
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|855,861|false|false|false|C0458827;C4071894|Airway structure;Chest>Airway|airway
Event|Event|SIMPLE_SEGMENT|867,873|false|false|false|||placed
Finding|Body Substance|SIMPLE_SEGMENT|882,889|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|882,889|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|882,889|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|894,905|false|false|false|||transported
Event|Event|SIMPLE_SEGMENT|913,922|false|false|false|||emergency
Finding|Finding|SIMPLE_SEGMENT|913,922|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Idea or Concept|SIMPLE_SEGMENT|913,922|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Intellectual Product|SIMPLE_SEGMENT|913,922|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Pathologic Function|SIMPLE_SEGMENT|913,922|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|913,922|false|false|false|C0013956|Emergency Situation|emergency
Procedure|Health Care Activity|SIMPLE_SEGMENT|913,922|false|false|false|C1553500|emergency encounter|emergency
Event|Event|SIMPLE_SEGMENT|924,934|false|false|false|||department
Finding|Idea or Concept|SIMPLE_SEGMENT|924,934|false|false|false|C1547537;C1548283;C1549615|Department - Charge type;Department - No suggested values defined;Organization Unit Type - Department|department
Event|Event|SIMPLE_SEGMENT|951,958|true|false|false|||reports
Finding|Intellectual Product|SIMPLE_SEGMENT|951,958|true|false|false|C0684224|Report (document)|reports
Procedure|Health Care Activity|SIMPLE_SEGMENT|951,958|true|false|false|C0700287|Reporting|reports
Finding|Finding|SIMPLE_SEGMENT|962,971|true|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Functional Concept|SIMPLE_SEGMENT|962,971|true|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Finding|SIMPLE_SEGMENT|962,980|true|false|false|C0574067|Increasing frequency of cough|increased coughing
Event|Event|SIMPLE_SEGMENT|972,980|true|false|false|||coughing
Finding|Sign or Symptom|SIMPLE_SEGMENT|972,980|true|false|false|C0010200|Coughing|coughing
Event|Event|SIMPLE_SEGMENT|985,993|true|false|false|||stooling
Finding|Body Substance|SIMPLE_SEGMENT|1010,1017|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1010,1017|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1010,1017|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|SIMPLE_SEGMENT|1010,1021|false|false|false|C0332310|Has patient|patient has
Finding|Functional Concept|SIMPLE_SEGMENT|1028,1039|false|false|false|C0231242|Complicated|complicated
Finding|Functional Concept|SIMPLE_SEGMENT|1040,1047|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|SIMPLE_SEGMENT|1040,1047|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|SIMPLE_SEGMENT|1040,1047|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1040,1047|false|false|false|C0199168|Medical service|medical
Event|Event|SIMPLE_SEGMENT|1048,1054|false|false|false|||course
Finding|Idea or Concept|SIMPLE_SEGMENT|1069,1074|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|SIMPLE_SEGMENT|1069,1074|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Event|Event|SIMPLE_SEGMENT|1084,1089|false|false|false|||brief
Finding|Intellectual Product|SIMPLE_SEGMENT|1084,1089|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|brief
Finding|Body Substance|SIMPLE_SEGMENT|1095,1102|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1095,1102|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1095,1102|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|1117,1126|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|1117,1126|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|1117,1126|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|1117,1126|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|1117,1126|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|1146,1160|false|false|false|||hosptilazation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1165,1179|false|true|false|C0238106|Clostridium difficile colitis|c.diff colitis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1172,1179|false|true|false|C0009319|Colitis|colitis
Event|Event|SIMPLE_SEGMENT|1172,1179|false|false|false|||colitis
Event|Event|SIMPLE_SEGMENT|1180,1191|false|false|false|||complicated
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1195,1201|false|false|false|C0036690;C0243026|Sepsis;Septicemia|sepsis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1219,1230|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|SIMPLE_SEGMENT|1219,1230|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|SIMPLE_SEGMENT|1219,1230|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|SIMPLE_SEGMENT|1219,1230|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1219,1238|false|false|false|C1145670|Respiratory Failure|respiratory failure
Event|Event|SIMPLE_SEGMENT|1231,1238|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|1231,1238|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|1231,1238|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|1231,1238|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|SIMPLE_SEGMENT|1249,1259|false|false|false|||intubation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1249,1259|false|false|false|C0021925|Intubation (procedure)|intubation
Finding|Idea or Concept|SIMPLE_SEGMENT|1270,1273|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|1270,1273|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|1284,1293|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|1284,1293|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|1284,1293|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|1284,1293|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|1284,1293|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|1304,1313|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|1304,1313|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Body Substance|SIMPLE_SEGMENT|1319,1326|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1319,1326|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1319,1326|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|1332,1337|false|false|false|||noted
Event|Event|SIMPLE_SEGMENT|1344,1355|false|false|false|||complaining
Event|Event|SIMPLE_SEGMENT|1359,1368|false|false|false|||worsening
Event|Event|SIMPLE_SEGMENT|1369,1372|false|false|false|||SOB
Finding|Sign or Symptom|SIMPLE_SEGMENT|1369,1372|false|false|false|C0013404|Dyspnea|SOB
Event|Event|SIMPLE_SEGMENT|1377,1380|false|false|false|||ABG
Finding|Gene or Genome|SIMPLE_SEGMENT|1377,1380|false|false|false|C1412045|A1BG gene|ABG
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1377,1380|false|false|false|C0150411|Analysis of arterial blood gases and pH|ABG
Event|Event|SIMPLE_SEGMENT|1410,1421|false|false|false|||re-admitted
Event|Event|SIMPLE_SEGMENT|1471,1476|false|false|false|||biPAP
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1471,1476|false|false|false|C1956423|Biphasic Continuous Positive Airway Pressure|biPAP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1481,1484|false|false|false|C1334032|HDAC1 protein, human|HD1
Drug|Enzyme|SIMPLE_SEGMENT|1481,1484|false|false|false|C1334032|HDAC1 protein, human|HD1
Finding|Gene or Genome|SIMPLE_SEGMENT|1481,1484|false|false|false|C1333891;C1706171;C4050150|HDAC1 gene;HDAC1 wt Allele;PLEC wt Allele|HD1
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1492,1498|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|1492,1498|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1492,1498|false|false|false|C0030054|oxygen|oxygen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1492,1498|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Event|Event|SIMPLE_SEGMENT|1499,1510|false|false|false|||requirement
Finding|Functional Concept|SIMPLE_SEGMENT|1499,1510|false|false|false|C1514873|Requirement|requirement
Event|Event|SIMPLE_SEGMENT|1523,1525|false|false|false|||2L
Event|Event|SIMPLE_SEGMENT|1536,1544|false|false|false|||etiology
Finding|Conceptual Entity|SIMPLE_SEGMENT|1536,1544|false|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|etiology
Finding|Functional Concept|SIMPLE_SEGMENT|1536,1544|false|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|etiology
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1564,1575|false|false|false|C0231832|Respiratory rate|respiratory
Event|Event|SIMPLE_SEGMENT|1564,1575|false|false|false|||respiratory
Finding|Body Substance|SIMPLE_SEGMENT|1564,1575|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|SIMPLE_SEGMENT|1564,1575|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|SIMPLE_SEGMENT|1564,1575|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Event|Event|SIMPLE_SEGMENT|1577,1584|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|1577,1584|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|1577,1584|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|1577,1584|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|SIMPLE_SEGMENT|1589,1593|false|false|false|||felt
Event|Event|SIMPLE_SEGMENT|1604,1619|false|false|false|||hypoventilation
Finding|Pathologic Function|SIMPLE_SEGMENT|1604,1619|false|false|false|C3203358|Hypoventilation|hypoventilation
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1625,1635|false|false|false|C2830004|Somnolence|somnolence
Event|Event|SIMPLE_SEGMENT|1625,1635|false|false|false|||somnolence
Finding|Finding|SIMPLE_SEGMENT|1625,1635|false|false|false|C0013144|Drowsiness|somnolence
Drug|Organic Chemical|SIMPLE_SEGMENT|1637,1644|false|false|false|C0163712|Relate - vinyl resin|related
Event|Event|SIMPLE_SEGMENT|1637,1644|false|false|false|||related
Finding|Finding|SIMPLE_SEGMENT|1637,1644|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|SIMPLE_SEGMENT|1637,1644|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Event|Event|SIMPLE_SEGMENT|1648,1660|false|false|false|||oversedation
Finding|Finding|SIMPLE_SEGMENT|1648,1660|false|false|false|C0542127|Oversedation|oversedation
Drug|Organic Chemical|SIMPLE_SEGMENT|1666,1673|false|false|false|C0527258|Zyprexa|zyprexa
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1666,1673|false|false|false|C0527258|Zyprexa|zyprexa
Event|Event|SIMPLE_SEGMENT|1684,1688|false|false|false|||held
Event|Event|SIMPLE_SEGMENT|1693,1702|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|1693,1702|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|1693,1702|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|1693,1702|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|1693,1702|false|false|false|C0030685|Patient Discharge|discharge
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1706,1709|true|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|SIMPLE_SEGMENT|1706,1709|true|false|false|||CTA
Finding|Gene or Genome|SIMPLE_SEGMENT|1706,1709|true|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1706,1709|true|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1710,1715|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Event|Event|SIMPLE_SEGMENT|1710,1715|true|false|false|||chest
Finding|Finding|SIMPLE_SEGMENT|1710,1715|true|false|false|C0741025|Chest problem|chest
Event|Event|SIMPLE_SEGMENT|1720,1728|true|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|1720,1728|true|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|1720,1728|true|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1720,1728|true|false|false|C5237010|Expression Negative|negative
Finding|Finding|SIMPLE_SEGMENT|1720,1732|true|false|false|C0205160|Negative|negative for
Event|Event|SIMPLE_SEGMENT|1740,1746|true|false|false|||showed
Event|Event|SIMPLE_SEGMENT|1750,1755|true|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|1750,1755|true|false|false|C1550016|Remote control command - Clear|clear
Event|Event|SIMPLE_SEGMENT|1757,1765|true|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|1757,1765|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|1757,1768|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1769,1778|true|false|false|C0032285|Pneumonia|pneumonia
Event|Event|SIMPLE_SEGMENT|1769,1778|true|false|false|||pneumonia
Event|Event|SIMPLE_SEGMENT|1799,1806|false|false|false|||started
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1810,1814|false|false|false|C0535219|SMC3 protein, human|HCAP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1810,1814|false|false|false|C0535219|SMC3 protein, human|HCAP
Event|Event|SIMPLE_SEGMENT|1810,1814|false|false|false|||HCAP
Finding|Gene or Genome|SIMPLE_SEGMENT|1810,1814|false|false|false|C1419431;C1422826;C1704469;C1822780|DCD gene;RNGTT gene;SMC3 gene;SMC3 wt Allele|HCAP
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1810,1814|false|false|false|C0056451|Cyclophosphamide/Altretamine/Doxorubicin/Cisplatin Regimen|HCAP
Drug|Antibiotic|SIMPLE_SEGMENT|1816,1827|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|SIMPLE_SEGMENT|1816,1827|false|false|false|||antibiotics
Drug|Antibiotic|SIMPLE_SEGMENT|1838,1846|false|false|false|C0055003|cefepime|cefepime
Drug|Organic Chemical|SIMPLE_SEGMENT|1838,1846|false|false|false|C0055003|cefepime|cefepime
Event|Event|SIMPLE_SEGMENT|1838,1846|false|false|false|||cefepime
Event|Event|SIMPLE_SEGMENT|1858,1865|false|false|false|||stopped
Event|Event|SIMPLE_SEGMENT|1884,1893|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|1884,1893|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|1884,1893|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|1884,1893|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|1884,1893|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|1909,1917|true|false|false|||cultures
Finding|Idea or Concept|SIMPLE_SEGMENT|1909,1917|true|false|false|C0010453|Culture (Anthropological)|cultures
Event|Event|SIMPLE_SEGMENT|1923,1931|true|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|1923,1931|true|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|1923,1931|true|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1923,1931|true|false|false|C5237010|Expression Negative|negative
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1950,1963|true|false|false|C0521530|Lung consolidation|consolidation
Event|Event|SIMPLE_SEGMENT|1950,1963|true|false|false|||consolidation
Event|Event|SIMPLE_SEGMENT|1967,1974|true|false|false|||imaging
Finding|Finding|SIMPLE_SEGMENT|1967,1974|true|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1967,1974|true|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Finding|Idea or Concept|SIMPLE_SEGMENT|1991,1998|false|false|false|C1555582|Initial (abbreviation)|initial
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|2022,2030|false|false|false|C0039155|Systole|systolic
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2031,2035|false|false|false|C0231832|Respiratory rate|Resp
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2031,2035|false|false|false|C0851355|Respiratory, thoracic and mediastinal disorders|Resp
Event|Event|SIMPLE_SEGMENT|2031,2035|false|false|false|||Resp
Event|Event|SIMPLE_SEGMENT|2041,2052|true|false|false|||spontaneous
Finding|Finding|SIMPLE_SEGMENT|2041,2065|true|false|false|C0412771|Spontaneous respiration|spontaneous respirations
Event|Event|SIMPLE_SEGMENT|2053,2065|true|false|false|||respirations
Finding|Physiologic Function|SIMPLE_SEGMENT|2053,2065|true|false|false|C0035203|Respiration|respirations
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2070,2073|false|false|false|C2744672|SAT1 protein, human|Sat
Drug|Enzyme|SIMPLE_SEGMENT|2070,2073|false|false|false|C2744672|SAT1 protein, human|Sat
Finding|Gene or Genome|SIMPLE_SEGMENT|2070,2073|false|false|false|C0871290;C1705827;C1822614|College Entrance Examination Board Scholastic Aptitude Test;SAT1 gene;SAT1 wt Allele|Sat
Finding|Intellectual Product|SIMPLE_SEGMENT|2070,2073|false|false|false|C0871290;C1705827;C1822614|College Entrance Examination Board Scholastic Aptitude Test;SAT1 gene;SAT1 wt Allele|Sat
Finding|Idea or Concept|SIMPLE_SEGMENT|2081,2088|false|false|false|C1555582|Initial (abbreviation)|Initial
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2089,2093|false|false|false|C0587081|Laboratory test finding|labs
Event|Event|SIMPLE_SEGMENT|2095,2107|false|false|false|||demonstrated
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2108,2111|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2108,2111|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|hct
Anatomy|Cell|SIMPLE_SEGMENT|2118,2121|false|false|false|C0023516|Leukocytes|wbc
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2128,2138|false|false|false|C0010294|creatinine|creatinine
Drug|Organic Chemical|SIMPLE_SEGMENT|2128,2138|false|false|false|C0010294|creatinine|creatinine
Event|Event|SIMPLE_SEGMENT|2128,2138|false|false|false|||creatinine
Finding|Physiologic Function|SIMPLE_SEGMENT|2128,2138|false|false|false|C4551889|Creatinine metabolic function|creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2128,2138|false|false|false|C0201975|Creatinine measurement|creatinine
Event|Event|SIMPLE_SEGMENT|2144,2147|false|false|false|||BIN
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2152,2158|false|false|false|C0023764|lipase|lipase
Drug|Enzyme|SIMPLE_SEGMENT|2152,2158|false|false|false|C0023764|lipase|lipase
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2152,2158|false|false|false|C0023764|lipase|lipase
Event|Event|SIMPLE_SEGMENT|2152,2158|false|false|false|||lipase
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2152,2158|false|false|false|C0373670|Lipase measurement|lipase
Drug|Organic Chemical|SIMPLE_SEGMENT|2168,2175|false|false|false|C0022924;C0376261|Lactates;lactate|lactate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2168,2175|false|false|false|C0022924;C0376261|Lactates;lactate|lactate
Event|Event|SIMPLE_SEGMENT|2168,2175|false|false|false|||lactate
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2168,2175|false|false|false|C0202115|Lactic acid measurement|lactate
Event|Event|SIMPLE_SEGMENT|2183,2186|false|false|false|||cxr
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2183,2186|false|false|false|C0039985|Plain chest X-ray|cxr
Event|Event|SIMPLE_SEGMENT|2187,2199|false|false|false|||demonstrated
Anatomy|Tissue|SIMPLE_SEGMENT|2210,2217|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2210,2217|false|false|false|C0032226|Pleural Diseases|pleural
Event|Event|SIMPLE_SEGMENT|2219,2228|false|false|false|||effusions
Finding|Pathologic Function|SIMPLE_SEGMENT|2219,2228|false|false|false|C0013687|effusion|effusions
Event|Event|SIMPLE_SEGMENT|2246,2258|false|false|false|||demonstrated
Finding|Gene or Genome|SIMPLE_SEGMENT|2259,2264|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|2272,2280|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Event|Event|SIMPLE_SEGMENT|2272,2280|false|false|false|||positive
Finding|Classification|SIMPLE_SEGMENT|2272,2280|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|SIMPLE_SEGMENT|2272,2280|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2282,2290|false|false|false|C0028137|Nitrites|nitrites
Drug|Inorganic Chemical|SIMPLE_SEGMENT|2282,2290|false|false|false|C0028137|Nitrites|nitrites
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2282,2290|false|false|false|C0028137|Nitrites|nitrites
Event|Event|SIMPLE_SEGMENT|2282,2290|false|false|false|||nitrites
Anatomy|Cell|SIMPLE_SEGMENT|2299,2302|false|false|false|C0023516|Leukocytes|wbc
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2309,2320|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|SIMPLE_SEGMENT|2309,2320|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|SIMPLE_SEGMENT|2309,2320|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|SIMPLE_SEGMENT|2309,2320|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2309,2328|false|false|false|C1145670|Respiratory Failure|respiratory failure
Event|Event|SIMPLE_SEGMENT|2321,2328|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|2321,2328|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|2321,2328|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|2321,2328|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Body Substance|SIMPLE_SEGMENT|2333,2340|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|2333,2340|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|2333,2340|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|2346,2355|false|false|false|||intubated
Finding|Finding|SIMPLE_SEGMENT|2346,2355|false|false|false|C4698386|Intubated|intubated
Finding|Idea or Concept|SIMPLE_SEGMENT|2364,2371|false|false|false|C1555582|Initial (abbreviation)|initial
Event|Event|SIMPLE_SEGMENT|2372,2375|false|false|false|||ABG
Finding|Gene or Genome|SIMPLE_SEGMENT|2372,2375|false|false|false|C1412045|A1BG gene|ABG
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2372,2375|false|false|false|C0150411|Analysis of arterial blood gases and pH|ABG
Finding|Gene or Genome|SIMPLE_SEGMENT|2410,2414|false|false|false|C3469826;C3470073|DESI1 gene;SLC35G1 gene|post
Event|Event|SIMPLE_SEGMENT|2416,2426|false|false|false|||intubation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2416,2426|false|false|false|C0021925|Intubation (procedure)|intubation
Finding|Body Substance|SIMPLE_SEGMENT|2433,2440|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|2433,2440|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|2433,2440|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2451,2461|false|false|false|C0042313|vancomycin|vancomycin
Drug|Antibiotic|SIMPLE_SEGMENT|2451,2461|false|false|false|C0042313|vancomycin|vancomycin
Event|Event|SIMPLE_SEGMENT|2451,2461|false|false|false|||vancomycin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2451,2461|false|false|false|C0489941|Vancomycin measurement|vancomycin
Drug|Antibiotic|SIMPLE_SEGMENT|2466,2474|false|false|false|C0055003|cefepime|cefepime
Drug|Organic Chemical|SIMPLE_SEGMENT|2466,2474|false|false|false|C0055003|cefepime|cefepime
Event|Event|SIMPLE_SEGMENT|2466,2474|false|false|false|||cefepime
Event|Event|SIMPLE_SEGMENT|2480,2488|false|false|false|||coverage
Finding|Functional Concept|SIMPLE_SEGMENT|2480,2488|false|false|false|C1551362;C1999244;C3854012|coverage - HL7PublishingDomain;coverage - financial contract|coverage
Finding|Idea or Concept|SIMPLE_SEGMENT|2480,2488|false|false|false|C1551362;C1999244;C3854012|coverage - HL7PublishingDomain;coverage - financial contract|coverage
Finding|Intellectual Product|SIMPLE_SEGMENT|2480,2488|false|false|false|C1551362;C1999244;C3854012|coverage - HL7PublishingDomain;coverage - financial contract|coverage
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2499,2506|false|false|false|C0042027|Urinary tract|urinary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2511,2520|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2511,2520|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|2511,2520|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Event|Event|SIMPLE_SEGMENT|2521,2527|false|false|false|||source
Finding|Finding|SIMPLE_SEGMENT|2521,2527|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Functional Concept|SIMPLE_SEGMENT|2521,2527|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Intellectual Product|SIMPLE_SEGMENT|2521,2527|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Event|Event|SIMPLE_SEGMENT|2534,2544|false|false|false|||intubation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2534,2544|false|false|false|C0021925|Intubation (procedure)|intubation
Event|Event|SIMPLE_SEGMENT|2553,2560|false|false|false|||dropped
Event|Event|SIMPLE_SEGMENT|2581,2588|false|false|false|||started
Drug|Organic Chemical|SIMPLE_SEGMENT|2592,2600|false|false|false|C0733815|Levophed|levophed
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2592,2600|false|false|false|C0733815|Levophed|levophed
Event|Event|SIMPLE_SEGMENT|2592,2600|false|false|false|||levophed
Drug|Organic Chemical|SIMPLE_SEGMENT|2606,2619|false|false|false|C0031469|phenylephrine|phenylephrine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2606,2619|false|false|false|C0031469|phenylephrine|phenylephrine
Event|Event|SIMPLE_SEGMENT|2606,2619|false|false|false|||phenylephrine
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2641,2645|false|false|false|C2049629|Peripherally Inserted Central Catheter Line Insertion|PICC
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2646,2650|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|2646,2650|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Substance|SIMPLE_SEGMENT|2646,2650|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Event|Event|SIMPLE_SEGMENT|2646,2650|false|false|false|||line
Finding|Intellectual Product|SIMPLE_SEGMENT|2646,2650|false|false|false|C1546701|line source specimen code|line
Event|Event|SIMPLE_SEGMENT|2652,2657|false|false|false|||Given
Event|Event|SIMPLE_SEGMENT|2662,2669|false|false|false|||altered
Finding|Functional Concept|SIMPLE_SEGMENT|2662,2669|false|false|false|C0392747|Changing|altered
Finding|Mental Process|SIMPLE_SEGMENT|2671,2677|false|false|false|C0229992|Psyche structure|mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2671,2684|false|false|false|C0488568;C0488569||mental status
Finding|Finding|SIMPLE_SEGMENT|2671,2684|false|false|false|C0278060|Mental state|mental status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2678,2684|false|false|false|C5889824||status
Event|Event|SIMPLE_SEGMENT|2678,2684|false|false|false|||status
Finding|Idea or Concept|SIMPLE_SEGMENT|2678,2684|false|false|false|C1546481|What subject filter - Status|status
Event|Activity|SIMPLE_SEGMENT|2688,2695|false|false|false|C1706079||arrival
Event|Event|SIMPLE_SEGMENT|2688,2695|false|false|false|||arrival
Finding|Functional Concept|SIMPLE_SEGMENT|2688,2695|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2699,2703|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2699,2703|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2699,2703|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2699,2703|false|false|false|C0876917|Procedure on head|head
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2699,2706|false|false|false|C0202691|CAT scan of head|head CT
Event|Event|SIMPLE_SEGMENT|2704,2706|false|false|false|||CT
Event|Event|SIMPLE_SEGMENT|2727,2733|true|false|false|||showed
Finding|Intellectual Product|SIMPLE_SEGMENT|2738,2743|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2744,2752|true|false|false|C2926606||findings
Event|Event|SIMPLE_SEGMENT|2744,2752|true|false|false|||findings
Finding|Functional Concept|SIMPLE_SEGMENT|2744,2752|true|false|false|C2607943|findings aspects|findings
Event|Event|SIMPLE_SEGMENT|2754,2760|false|false|false|||Vitals
Event|Event|SIMPLE_SEGMENT|2764,2772|false|false|false|||transfer
Finding|Functional Concept|SIMPLE_SEGMENT|2764,2772|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|SIMPLE_SEGMENT|2764,2772|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|SIMPLE_SEGMENT|2764,2772|false|false|false|C4706767|Transfer (immobility management)|transfer
Event|Event|SIMPLE_SEGMENT|2812,2820|false|false|false|||settings
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2827,2831|false|false|false|C3484065||fio2
Event|Event|SIMPLE_SEGMENT|2827,2831|false|false|false|||fio2
Finding|Finding|SIMPLE_SEGMENT|2827,2831|false|false|false|C0428167|Fraction of inspired oxygen|fio2
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2827,2831|false|false|false|C1512797;C2370852|Inspired Oxygen Fraction Test;fraction of inspired oxygen (FiO2) (treatment)|fio2
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2827,2831|false|false|false|C1512797;C2370852|Inspired Oxygen Fraction Test;fraction of inspired oxygen (FiO2) (treatment)|fio2
Event|Event|SIMPLE_SEGMENT|2849,2853|false|false|false|||peep
Finding|Finding|SIMPLE_SEGMENT|2849,2853|false|false|false|C3494516|Positive end expiratory pressure (finding)|peep
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2849,2853|false|false|false|C0032740|Positive End-Expiratory Pressure|peep
Event|Event|SIMPLE_SEGMENT|2857,2865|false|false|false|||Sedation
Finding|Finding|SIMPLE_SEGMENT|2857,2865|false|false|false|C0235195;C5400562|Sedated state;Sedation|Sedation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2857,2865|false|false|false|C0344106|Sedation procedure|Sedation
Drug|Organic Chemical|SIMPLE_SEGMENT|2872,2881|false|false|false|C0026056|midazolam|midazolam
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2872,2881|false|false|false|C0026056|midazolam|midazolam
Event|Event|SIMPLE_SEGMENT|2872,2881|false|false|false|||midazolam
Drug|Organic Chemical|SIMPLE_SEGMENT|2886,2894|false|false|false|C0015846|fentanyl|fentanyl
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2886,2894|false|false|false|C0015846|fentanyl|fentanyl
Event|Event|SIMPLE_SEGMENT|2886,2894|false|false|false|||fentanyl
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2886,2894|false|false|false|C0524136|Fentanyl measurement|fentanyl
Event|Event|SIMPLE_SEGMENT|2904,2915|false|false|false|||transferred
Drug|Organic Chemical|SIMPLE_SEGMENT|2919,2927|false|false|false|C0733815|Levophed|levophed
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2919,2927|false|false|false|C0733815|Levophed|levophed
Event|Event|SIMPLE_SEGMENT|2928,2933|false|false|false|||alone
Finding|Finding|SIMPLE_SEGMENT|2928,2933|false|false|false|C0439044|Living Alone|alone
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2938,2942|false|false|false|C0026045|Microtubule-Associated Proteins|MAPs
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2938,2942|false|false|false|C0026045|Microtubule-Associated Proteins|MAPs
Event|Event|SIMPLE_SEGMENT|2938,2942|false|false|false|||MAPs
Finding|Gene or Genome|SIMPLE_SEGMENT|2938,2942|false|false|false|C0024779;C1824157|C3orf62 gene;Map|MAPs
Finding|Intellectual Product|SIMPLE_SEGMENT|2938,2942|false|false|false|C0024779;C1824157|C3orf62 gene;Map|MAPs
Event|Activity|SIMPLE_SEGMENT|2956,2963|false|false|false|C1706079||arrival
Event|Event|SIMPLE_SEGMENT|2956,2963|false|false|false|||arrival
Finding|Functional Concept|SIMPLE_SEGMENT|2956,2963|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Event|Event|SIMPLE_SEGMENT|2978,2984|false|false|false|||vitals
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3031,3035|false|false|false|C3484065||FiO2
Event|Event|SIMPLE_SEGMENT|3031,3035|false|false|false|||FiO2
Finding|Finding|SIMPLE_SEGMENT|3031,3035|false|false|false|C0428167|Fraction of inspired oxygen|FiO2
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3031,3035|false|false|false|C1512797;C2370852|Inspired Oxygen Fraction Test;fraction of inspired oxygen (FiO2) (treatment)|FiO2
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3031,3035|false|false|false|C1512797;C2370852|Inspired Oxygen Fraction Test;fraction of inspired oxygen (FiO2) (treatment)|FiO2
Finding|Body Substance|SIMPLE_SEGMENT|3042,3049|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|3042,3049|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|3042,3049|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Organic Chemical|SIMPLE_SEGMENT|3059,3067|true|false|false|C0733815|Levophed|levophed
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3059,3067|true|false|false|C0733815|Levophed|levophed
Event|Event|SIMPLE_SEGMENT|3068,3072|true|false|false|||drip
Event|Event|SIMPLE_SEGMENT|3083,3090|true|false|false|||sedated
Finding|Finding|SIMPLE_SEGMENT|3083,3090|true|false|false|C0235195|Sedated state|sedated
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|3096,3108|true|false|false|C0752295|Confusional Arousals|unresponsive
Event|Event|SIMPLE_SEGMENT|3096,3108|true|false|false|||unresponsive
Finding|Finding|SIMPLE_SEGMENT|3096,3108|true|false|false|C0205269;C0237284|Unresponsive to Treatment;unresponsive behavior|unresponsive
Finding|Functional Concept|SIMPLE_SEGMENT|3096,3108|true|false|false|C0205269;C0237284|Unresponsive to Treatment;unresponsive behavior|unresponsive
Event|Event|SIMPLE_SEGMENT|3112,3118|true|false|false|||verbal
Finding|Functional Concept|SIMPLE_SEGMENT|3112,3118|true|false|false|C1548941|Participation Mode - verbal|verbal
Procedure|Health Care Activity|SIMPLE_SEGMENT|3112,3118|true|false|false|C1608381|Consent Mode - Verbal|verbal
Finding|Sign or Symptom|SIMPLE_SEGMENT|3123,3130|false|false|false|C0030193|Pain|painful
Event|Event|SIMPLE_SEGMENT|3131,3138|false|false|false|||stimuli
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|3131,3138|false|false|false|C0234402|Stimulus|stimuli
Event|Event|SIMPLE_SEGMENT|3145,3152|false|false|false|||thought
Finding|Idea or Concept|SIMPLE_SEGMENT|3145,3152|false|false|false|C0039869;C4319827|Thought|thought
Finding|Mental Process|SIMPLE_SEGMENT|3145,3152|false|false|false|C0039869;C4319827|Thought|thought
Finding|Intellectual Product|SIMPLE_SEGMENT|3163,3168|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|brief
Event|Event|SIMPLE_SEGMENT|3169,3176|false|false|false|||episode
Finding|Finding|SIMPLE_SEGMENT|3180,3201|false|false|false|C0011103;C0231474|Decerebrate Posturing;Decerebrate State|decerebrate posturing
Finding|Pathologic Function|SIMPLE_SEGMENT|3180,3201|false|false|false|C0011103;C0231474|Decerebrate Posturing;Decerebrate State|decerebrate posturing
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3192,3201|false|false|false|C0872410|Posturing|posturing
Event|Event|SIMPLE_SEGMENT|3192,3201|false|false|false|||posturing
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3212,3229|false|false|false|C1140618|Upper Extremity|upper extremities
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3218,3229|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Event|Event|SIMPLE_SEGMENT|3234,3240|false|false|false|||Review
Finding|Idea or Concept|SIMPLE_SEGMENT|3234,3240|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|Review
Finding|Intellectual Product|SIMPLE_SEGMENT|3234,3240|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|Review
Finding|Functional Concept|SIMPLE_SEGMENT|3234,3243|false|false|false|C0699752|Review of|Review of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3234,3251|false|false|false|C0488564;C0488565||Review of systems
Procedure|Health Care Activity|SIMPLE_SEGMENT|3234,3251|false|false|false|C0489633|Review of systems (procedure)|Review of systems
Event|Event|SIMPLE_SEGMENT|3244,3251|false|false|false|||systems
Finding|Functional Concept|SIMPLE_SEGMENT|3244,3251|false|false|false|C0449913|System|systems
Event|Event|SIMPLE_SEGMENT|3254,3260|false|false|false|||Unable
Finding|Finding|SIMPLE_SEGMENT|3254,3260|false|false|false|C1299582|Unable|Unable
Event|Activity|SIMPLE_SEGMENT|3264,3270|false|false|false|C1706701|Acquisition (action)|Obtain
Event|Event|SIMPLE_SEGMENT|3264,3270|false|false|false|||Obtain
Finding|Functional Concept|SIMPLE_SEGMENT|3264,3270|false|false|false|C1301820|Obtain|Obtain
Finding|Finding|SIMPLE_SEGMENT|3274,3294|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|3279,3286|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|3279,3286|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|3279,3286|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|3279,3286|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|3279,3286|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|3279,3294|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|3287,3294|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|3287,3294|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|3287,3294|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3296,3302|false|false|false|C0002871|Anemia|Anemia
Event|Event|SIMPLE_SEGMENT|3296,3302|false|false|false|||Anemia
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3305,3327|false|false|false|C0694540|borderline cholesterol|Borderline cholesterol
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3316,3327|false|false|false|C0008377|cholesterol|cholesterol
Drug|Organic Chemical|SIMPLE_SEGMENT|3316,3327|false|false|false|C0008377|cholesterol|cholesterol
Event|Event|SIMPLE_SEGMENT|3316,3327|false|false|false|||cholesterol
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3316,3327|false|false|false|C0201950|Cholesterol measurement|cholesterol
Finding|Sign or Symptom|SIMPLE_SEGMENT|3350,3360|false|false|false|C0016204|Flatulence|Flatulence
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3363,3368|false|false|false|C0018787;C4037974|Chest>Heart;Heart|Heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3363,3368|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|Heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|3363,3368|false|false|false|C0795691|HEART PROBLEM|Heart
Finding|Finding|SIMPLE_SEGMENT|3363,3375|false|false|false|C0018808|Heart murmur|Heart Murmur
Event|Event|SIMPLE_SEGMENT|3369,3375|false|false|false|||Murmur
Finding|Finding|SIMPLE_SEGMENT|3369,3375|false|false|false|C0018808|Heart murmur|Murmur
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3378,3390|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|SIMPLE_SEGMENT|3378,3390|false|false|false|||Hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3393,3407|false|false|false|C0020676|Hypothyroidism|Hypothyroidism
Event|Event|SIMPLE_SEGMENT|3393,3407|false|false|false|||Hypothyroidism
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3410,3430|false|false|false|C0026266|Mitral Valve Insufficiency|Mitral Regurgitation
Event|Event|SIMPLE_SEGMENT|3417,3430|false|false|false|||Regurgitation
Finding|Finding|SIMPLE_SEGMENT|3417,3430|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|Regurgitation
Finding|Sign or Symptom|SIMPLE_SEGMENT|3417,3430|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|Regurgitation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|3417,3430|false|false|false|C0460152|Regurgitation - mechanism|Regurgitation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3433,3445|false|false|false|C0029456|Osteoporosis|Osteoporosis
Event|Event|SIMPLE_SEGMENT|3433,3445|false|false|false|||Osteoporosis
Finding|Finding|SIMPLE_SEGMENT|3433,3445|false|false|false|C2911643|Encounter due to family history of osteoporosis|Osteoporosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3448,3457|false|false|false|C0032285|Pneumonia|Pneumonia
Event|Event|SIMPLE_SEGMENT|3448,3457|false|false|false|||Pneumonia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3460,3469|false|false|false|C0037199|Sinusitis|Sinusitis
Event|Event|SIMPLE_SEGMENT|3460,3469|false|false|false|||Sinusitis
Finding|Functional Concept|SIMPLE_SEGMENT|3484,3490|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|3484,3498|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|3491,3498|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|3491,3498|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|3491,3498|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|3491,3498|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|3504,3510|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|3504,3510|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|3504,3510|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|3504,3510|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|3504,3518|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|3511,3518|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|3511,3518|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|3511,3518|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|3511,3518|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Event|Event|SIMPLE_SEGMENT|3525,3532|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|3525,3532|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|3525,3532|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|3525,3532|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|3525,3535|false|false|false|C0262926|Medical History|history of
Finding|Finding|SIMPLE_SEGMENT|3525,3548|false|false|false|C0455527||history of hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3536,3548|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|SIMPLE_SEGMENT|3536,3548|false|false|false|||hypertension
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3553,3563|false|false|false|C3812393|ErbB Receptors|her family
Drug|Enzyme|SIMPLE_SEGMENT|3553,3563|false|false|false|C3812393|ErbB Receptors|her family
Finding|Receptor|SIMPLE_SEGMENT|3553,3563|false|false|false|C3812393|ErbB Receptors|her family
Event|Event|SIMPLE_SEGMENT|3557,3563|false|false|false|||family
Finding|Classification|SIMPLE_SEGMENT|3557,3563|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|3557,3563|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|3557,3563|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|3557,3563|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|3566,3572|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|SIMPLE_SEGMENT|3566,3572|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Classification|SIMPLE_SEGMENT|3575,3581|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|3575,3581|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|3575,3581|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|3575,3581|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Event|Event|SIMPLE_SEGMENT|3589,3596|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|3589,3596|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|3589,3596|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|3589,3596|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|3589,3599|false|false|false|C0262926|Medical History|history of
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3609,3616|false|false|false|C0006826|Malignant Neoplasms|cancers
Event|Event|SIMPLE_SEGMENT|3609,3616|false|false|false|||cancers
Event|Event|SIMPLE_SEGMENT|3629,3640|false|false|false|||grandfather
Event|Event|SIMPLE_SEGMENT|3649,3656|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|3649,3656|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|3649,3656|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|3649,3656|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|3649,3659|false|false|false|C0262926|Medical History|history of
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3660,3667|false|false|false|C0038351;C3714551;C4266636|Abdomen>Stomach;Stomach;Stomach structure|stomach
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3660,3667|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3660,3667|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Event|Event|SIMPLE_SEGMENT|3660,3667|false|false|false|||stomach
Finding|Finding|SIMPLE_SEGMENT|3660,3667|false|false|false|C0577027|Stomach problem|stomach
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3660,3667|false|false|false|C0872393|Procedure on stomach|stomach
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3660,3674|false|false|false|C0024623;C0699791|Malignant neoplasm of stomach;Stomach Carcinoma|stomach cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3668,3674|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|SIMPLE_SEGMENT|3668,3674|false|false|false|||cancer
Event|Event|SIMPLE_SEGMENT|3695,3702|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|3695,3702|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|3695,3702|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|3695,3702|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|3695,3705|false|false|false|C0262926|Medical History|history of
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3706,3712|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3706,3712|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3706,3712|false|false|false|C1950455|Throat Homeopathic Medication|throat
Event|Event|SIMPLE_SEGMENT|3706,3712|false|false|false|||throat
Finding|Body Substance|SIMPLE_SEGMENT|3706,3712|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Finding|Intellectual Product|SIMPLE_SEGMENT|3706,3712|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3714,3720|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|SIMPLE_SEGMENT|3714,3720|false|false|false|||cancer
Event|Event|SIMPLE_SEGMENT|3726,3733|true|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|3726,3733|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|3726,3733|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|3726,3733|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|3726,3736|true|false|false|C0262926|Medical History|history of
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3737,3742|true|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3737,3742|true|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3737,3742|true|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Finding|Finding|SIMPLE_SEGMENT|3737,3742|true|false|false|C0750873|COLON PROBLEM|colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3737,3750|true|false|false|C0007102|Malignant tumor of colon|colon cancers
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3743,3750|true|false|false|C0006826|Malignant Neoplasms|cancers
Event|Event|SIMPLE_SEGMENT|3743,3750|true|false|false|||cancers
Finding|Conceptual Entity|SIMPLE_SEGMENT|3752,3758|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|SIMPLE_SEGMENT|3752,3758|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3763,3769|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|SIMPLE_SEGMENT|3763,3769|false|false|false|||stroke
Finding|Finding|SIMPLE_SEGMENT|3763,3769|false|false|false|C5977286|Stroke (heart beat)|stroke
Finding|Classification|SIMPLE_SEGMENT|3775,3781|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|3775,3781|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|3775,3781|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|3775,3781|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|3790,3796|false|false|false|C1546508|Relationship - Mother|Mother
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3803,3808|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3803,3808|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|3803,3808|false|false|false|C0795691|HEART PROBLEM|heart
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3803,3814|false|false|false|C0018826;C1305961|Heart Valves|heart valve
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3809,3814|false|false|false|C1186983|Anatomical valve|valve
Event|Event|SIMPLE_SEGMENT|3815,3823|false|false|false|||replaced
Event|Event|SIMPLE_SEGMENT|3828,3836|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|3828,3836|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|3828,3836|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|3828,3836|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|3828,3841|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3828,3841|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|3837,3841|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|3837,3841|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3837,3841|false|false|false|C0582103|Medical Examination|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3843,3852|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|SIMPLE_SEGMENT|3853,3861|false|false|false|||PHYSICAL
Finding|Finding|SIMPLE_SEGMENT|3853,3861|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|SIMPLE_SEGMENT|3853,3861|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|3853,3861|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|SIMPLE_SEGMENT|3853,3866|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|3853,3866|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Event|Event|SIMPLE_SEGMENT|3862,3866|false|false|false|||EXAM
Finding|Functional Concept|SIMPLE_SEGMENT|3862,3866|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|3862,3866|false|false|false|C0582103|Medical Examination|EXAM
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3908,3912|false|false|false|C3484065||FiO2
Event|Event|SIMPLE_SEGMENT|3908,3912|false|false|false|||FiO2
Finding|Finding|SIMPLE_SEGMENT|3908,3912|false|false|false|C0428167|Fraction of inspired oxygen|FiO2
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3908,3912|false|false|false|C1512797;C2370852|Inspired Oxygen Fraction Test;fraction of inspired oxygen (FiO2) (treatment)|FiO2
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3908,3912|false|false|false|C1512797;C2370852|Inspired Oxygen Fraction Test;fraction of inspired oxygen (FiO2) (treatment)|FiO2
Event|Event|SIMPLE_SEGMENT|3915,3922|false|false|false|||General
Finding|Classification|SIMPLE_SEGMENT|3915,3922|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|SIMPLE_SEGMENT|3915,3922|false|false|false|C3812897|General medical service|General
Event|Event|SIMPLE_SEGMENT|3924,3933|false|false|false|||Intubated
Finding|Finding|SIMPLE_SEGMENT|3924,3933|false|false|false|C4698386|Intubated|Intubated
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|3935,3947|false|false|false|C0752295|Confusional Arousals|unresponsive
Event|Event|SIMPLE_SEGMENT|3935,3947|false|false|false|||unresponsive
Finding|Finding|SIMPLE_SEGMENT|3935,3947|false|false|false|C0205269;C0237284|Unresponsive to Treatment;unresponsive behavior|unresponsive
Finding|Functional Concept|SIMPLE_SEGMENT|3935,3947|false|false|false|C0205269;C0237284|Unresponsive to Treatment;unresponsive behavior|unresponsive
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3949,3953|false|false|false|C4750744|Acute limbic encephalitis following transplant|pale
Event|Event|SIMPLE_SEGMENT|3949,3953|false|false|false|||pale
Finding|Finding|SIMPLE_SEGMENT|3949,3953|false|false|false|C0241137;C0678215|Body pale (finding);Pallor of skin|pale
Event|Event|SIMPLE_SEGMENT|3960,3964|false|false|false|||thin
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3967,3972|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3974,3980|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3974,3980|false|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|SIMPLE_SEGMENT|3974,3980|false|false|false|||Sclera
Procedure|Health Care Activity|SIMPLE_SEGMENT|3974,3980|false|false|false|C2228481|examination of sclera|Sclera
Event|Event|SIMPLE_SEGMENT|3981,3990|false|false|false|||anicteric
Finding|Finding|SIMPLE_SEGMENT|3981,3990|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3992,3995|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3992,3995|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3997,4007|false|false|false|C0521367|Oropharyngeal|oropharynx
Event|Event|SIMPLE_SEGMENT|4008,4013|false|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|4008,4013|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4015,4021|false|false|false|C0034121|Pupil|pupils
Event|Event|SIMPLE_SEGMENT|4023,4034|false|false|false|||constricted
Finding|Finding|SIMPLE_SEGMENT|4023,4034|false|false|false|C1444778|Constricting sensation quality|constricted
Finding|Finding|SIMPLE_SEGMENT|4039,4047|false|false|false|C3842079|Sluggish|sluggish
Event|Event|SIMPLE_SEGMENT|4064,4071|false|false|false|||dobhoff
Finding|Finding|SIMPLE_SEGMENT|4084,4091|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|SIMPLE_SEGMENT|4084,4091|false|false|false|C0150312;C0449450|Present;Presentation|present
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4094,4098|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|SIMPLE_SEGMENT|4094,4098|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|SIMPLE_SEGMENT|4094,4098|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|SIMPLE_SEGMENT|4100,4106|true|false|false|||supple
Finding|Functional Concept|SIMPLE_SEGMENT|4100,4106|true|false|false|C0332254|Supple|supple
Event|Event|SIMPLE_SEGMENT|4108,4111|true|false|false|||JVP
Finding|Finding|SIMPLE_SEGMENT|4108,4111|true|false|false|C0428897|Jugular venous pressure|JVP
Event|Event|SIMPLE_SEGMENT|4116,4124|true|false|false|||elevated
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4129,4132|true|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4129,4132|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|SIMPLE_SEGMENT|4129,4132|true|false|false|||LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|4129,4132|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Activity|SIMPLE_SEGMENT|4147,4151|false|false|false|C0871208|Rating (action)|rate
Event|Event|SIMPLE_SEGMENT|4147,4151|false|false|false|||rate
Finding|Idea or Concept|SIMPLE_SEGMENT|4147,4151|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|SIMPLE_SEGMENT|4156,4162|false|false|false|||rhythm
Finding|Finding|SIMPLE_SEGMENT|4156,4162|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|SIMPLE_SEGMENT|4156,4162|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Event|Event|SIMPLE_SEGMENT|4195,4198|false|false|false|||SEM
Finding|Finding|SIMPLE_SEGMENT|4195,4198|false|false|false|C0694547|SYSTOLIC EJECTION MURMUR|SEM
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4200,4204|false|false|false|C0339510|Vitelliform Macular Dystrophy|best
Event|Event|SIMPLE_SEGMENT|4200,4204|false|false|false|||best
Finding|Gene or Genome|SIMPLE_SEGMENT|4200,4204|false|false|false|C1826421;C5781213|BEST1 gene;BEST1 wt Allele|best
Event|Event|SIMPLE_SEGMENT|4205,4210|false|false|false|||heard
Event|Event|SIMPLE_SEGMENT|4220,4223|false|false|false|||LSB
Anatomy|Cell Component|SIMPLE_SEGMENT|4237,4244|false|false|false|C1660780|midline cell component|midline
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4237,4253|false|false|false|C5389501|midline catheter (treatment)|midline catheter
Event|Event|SIMPLE_SEGMENT|4245,4253|false|false|false|||catheter
Finding|Intellectual Product|SIMPLE_SEGMENT|4245,4253|false|false|false|C1546572||catheter
Event|Event|SIMPLE_SEGMENT|4254,4261|false|false|false|||present
Finding|Finding|SIMPLE_SEGMENT|4254,4261|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|SIMPLE_SEGMENT|4254,4261|false|false|false|C0150312;C0449450|Present;Presentation|present
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4271,4276|false|false|false|C4048756|Right arm|R arm
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4273,4276|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|4273,4276|false|false|false|C3495676|Anorectal Malformations|arm
Event|Event|SIMPLE_SEGMENT|4273,4276|false|false|false|||arm
Finding|Gene or Genome|SIMPLE_SEGMENT|4273,4276|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4273,4276|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|SIMPLE_SEGMENT|4273,4276|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4273,4276|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4277,4282|false|false|false|C0024109|Lung|Lungs
Finding|Finding|SIMPLE_SEGMENT|4294,4302|true|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Finding|Functional Concept|SIMPLE_SEGMENT|4313,4324|true|false|false|C0205359|Spontaneous|spontaneous
Finding|Finding|SIMPLE_SEGMENT|4313,4337|true|false|false|C0412771|Spontaneous respiration|spontaneous respirations
Event|Event|SIMPLE_SEGMENT|4325,4337|true|false|false|||respirations
Finding|Physiologic Function|SIMPLE_SEGMENT|4325,4337|true|false|false|C0035203|Respiration|respirations
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4352,4355|false|false|false|C1266159|Trophoblastic tumor, epithelioid|ETT
Event|Event|SIMPLE_SEGMENT|4352,4355|false|false|false|||ETT
Event|Activity|SIMPLE_SEGMENT|4360,4365|false|false|false|C1882509|put - instruction imperative|place
Event|Event|SIMPLE_SEGMENT|4360,4365|false|false|false|||place
Finding|Functional Concept|SIMPLE_SEGMENT|4360,4365|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|SIMPLE_SEGMENT|4360,4365|false|false|false|C1533810||place
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4367,4374|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4367,4374|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Event|Event|SIMPLE_SEGMENT|4367,4374|false|false|false|||Abdomen
Finding|Finding|SIMPLE_SEGMENT|4367,4374|false|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4376,4380|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|SIMPLE_SEGMENT|4376,4380|false|false|false|||soft
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4397,4402|true|false|false|C0021853|Intestines|bowel
Finding|Finding|SIMPLE_SEGMENT|4397,4409|true|false|false|C0232693|Bowel sounds|bowel sounds
Event|Event|SIMPLE_SEGMENT|4403,4409|true|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|4403,4409|true|false|false|C0037709||sounds
Finding|Finding|SIMPLE_SEGMENT|4410,4417|true|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|SIMPLE_SEGMENT|4410,4417|true|false|false|C0150312;C0449450|Present;Presentation|present
Event|Event|SIMPLE_SEGMENT|4423,4435|true|false|false|||organomegaly
Finding|Finding|SIMPLE_SEGMENT|4423,4435|true|false|false|C4054315|Organomegaly|organomegaly
Event|Event|SIMPLE_SEGMENT|4448,4455|false|false|false|||present
Finding|Finding|SIMPLE_SEGMENT|4448,4455|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|SIMPLE_SEGMENT|4448,4455|false|false|false|C0150312;C0449450|Present;Presentation|present
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4477,4481|false|false|false|C5779629|Eruption of skin (disorder)|rash
Event|Event|SIMPLE_SEGMENT|4477,4481|false|false|false|||rash
Finding|Pathologic Function|SIMPLE_SEGMENT|4477,4481|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|SIMPLE_SEGMENT|4477,4481|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4490,4495|false|false|false|C0018246;C0816951;C4266533|Inguinal part of abdomen;Inguinal region;Pelvis>Groin|groin
Event|Governmental or Regulatory Activity|SIMPLE_SEGMENT|4496,4500|false|false|false|C1510751|Academic Research Enhancement Awards|area
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4512,4518|false|false|false|C0032861;C1382110|Powder dose form;powder physical state|powder
Drug|Substance|SIMPLE_SEGMENT|4512,4518|false|false|false|C0032861;C1382110|Powder dose form;powder physical state|powder
Event|Event|SIMPLE_SEGMENT|4512,4518|false|false|false|||powder
Event|Event|SIMPLE_SEGMENT|4520,4521|false|false|false|||/
Drug|Organic Chemical|SIMPLE_SEGMENT|4523,4533|false|false|false|C0025942|miconazole|miconazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4523,4533|false|false|false|C0025942|miconazole|miconazole
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4534,4540|false|false|false|C0032861;C1382110|Powder dose form;powder physical state|powder
Drug|Substance|SIMPLE_SEGMENT|4534,4540|false|false|false|C0032861;C1382110|Powder dose form;powder physical state|powder
Event|Event|SIMPLE_SEGMENT|4534,4540|false|false|false|||powder
Event|Event|SIMPLE_SEGMENT|4541,4548|false|false|false|||present
Finding|Finding|SIMPLE_SEGMENT|4541,4548|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|SIMPLE_SEGMENT|4541,4548|false|false|false|C0150312;C0449450|Present;Presentation|present
Event|Event|SIMPLE_SEGMENT|4564,4576|false|false|false|||distribution
Finding|Cell Function|SIMPLE_SEGMENT|4564,4576|false|false|false|C1704711;C5779816|Distribution;Distribution [PK]|distribution
Finding|Functional Concept|SIMPLE_SEGMENT|4564,4576|false|false|false|C1704711;C5779816|Distribution;Distribution [PK]|distribution
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|4579,4582|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|SIMPLE_SEGMENT|4579,4582|false|false|false|||Ext
Finding|Gene or Genome|SIMPLE_SEGMENT|4579,4582|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|SIMPLE_SEGMENT|4584,4588|false|false|false|||warm
Finding|Finding|SIMPLE_SEGMENT|4584,4588|false|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|4584,4588|false|false|false|C0687712|warming process|warm
Finding|Finding|SIMPLE_SEGMENT|4590,4594|true|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|4595,4603|true|false|false|||perfused
Drug|Food|SIMPLE_SEGMENT|4608,4614|true|false|false|C5890763||pulses
Event|Event|SIMPLE_SEGMENT|4608,4614|true|false|false|||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|4608,4614|true|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|4608,4614|true|false|false|C0034107|Pulse taking|pulses
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|4619,4627|true|false|false|C0149651|Clubbing|clubbing
Event|Event|SIMPLE_SEGMENT|4619,4627|true|false|false|||clubbing
Event|Event|SIMPLE_SEGMENT|4629,4637|true|false|false|||cyanosis
Finding|Sign or Symptom|SIMPLE_SEGMENT|4629,4637|true|false|false|C0010520|Cyanosis|cyanosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4642,4647|true|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|4642,4647|true|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|4642,4647|true|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|4657,4663|false|false|false|||Unable
Finding|Finding|SIMPLE_SEGMENT|4657,4663|false|false|false|C1299582|Unable|Unable
Event|Event|SIMPLE_SEGMENT|4673,4681|false|false|false|||evaluate
Event|Event|SIMPLE_SEGMENT|4689,4705|false|false|false|||unresponsiveness
Finding|Finding|SIMPLE_SEGMENT|4689,4705|false|false|false|C0241526|Unresponsiveness|unresponsiveness
Finding|Body Substance|SIMPLE_SEGMENT|4713,4720|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|4713,4720|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|4713,4720|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|SIMPLE_SEGMENT|4713,4724|false|false|false|C0332310|Has patient|patient has
Event|Event|SIMPLE_SEGMENT|4728,4732|false|false|false|||DTRs
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4749,4764|false|false|false|C0278454|All extremities|all extremities
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4753,4764|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Event|Event|SIMPLE_SEGMENT|4767,4780|false|false|false|||decerebration
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4767,4780|false|false|false|C0178583|Decerebration procedure|decerebration
Event|Event|SIMPLE_SEGMENT|4789,4794|false|false|false|||noted
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4803,4820|false|false|false|C1140618|Upper Extremity|upper extremities
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4809,4820|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Finding|Body Substance|SIMPLE_SEGMENT|4826,4835|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|4826,4835|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|4826,4835|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|4826,4835|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|SIMPLE_SEGMENT|4836,4844|false|false|false|||PHYSICAL
Finding|Finding|SIMPLE_SEGMENT|4836,4844|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|SIMPLE_SEGMENT|4836,4844|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|4836,4844|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|SIMPLE_SEGMENT|4836,4849|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|4836,4849|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Event|Event|SIMPLE_SEGMENT|4845,4849|false|false|false|||EXAM
Finding|Functional Concept|SIMPLE_SEGMENT|4845,4849|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|4845,4849|false|false|false|C0582103|Medical Examination|EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|4877,4886|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|SIMPLE_SEGMENT|4887,4891|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4887,4891|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4906,4911|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4906,4911|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4906,4911|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|4912,4915|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|4922,4925|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4922,4925|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4922,4925|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4932,4935|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4932,4935|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|4932,4935|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4932,4935|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4941,4944|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4941,4944|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|4952,4955|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|4952,4955|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4952,4955|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4952,4955|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4952,4955|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|4961,4964|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4961,4964|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|4961,4964|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|4961,4964|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|4961,4964|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4961,4964|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|4970,4974|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4970,4974|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4991,4994|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5011,5016|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5011,5016|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5011,5016|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5021,5024|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|SIMPLE_SEGMENT|5021,5024|false|false|false|||PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5021,5024|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5047,5052|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5047,5052|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5047,5052|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5065,5070|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5065,5070|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5065,5070|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|5065,5078|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5065,5078|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5065,5078|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5071,5078|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|5071,5078|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5071,5078|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|5071,5078|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5071,5078|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5071,5078|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5123,5127|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5123,5127|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5123,5127|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5151,5156|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5151,5156|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5151,5156|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5160,5163|false|false|false|C0010287|Creatine Kinase|CPK
Drug|Enzyme|SIMPLE_SEGMENT|5160,5163|false|false|false|C0010287|Creatine Kinase|CPK
Event|Event|SIMPLE_SEGMENT|5160,5163|false|false|false|||CPK
Finding|Gene or Genome|SIMPLE_SEGMENT|5160,5163|false|false|false|C1418571|PIK3C2A gene|CPK
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5160,5163|false|false|false|C0201973|Creatine kinase measurement|CPK
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5181,5186|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5181,5186|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5181,5186|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5187,5193|false|false|false|C0023764|lipase|Lipase
Drug|Enzyme|SIMPLE_SEGMENT|5187,5193|false|false|false|C0023764|lipase|Lipase
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5187,5193|false|false|false|C0023764|lipase|Lipase
Event|Event|SIMPLE_SEGMENT|5187,5193|false|false|false|||Lipase
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5187,5193|false|false|false|C0373670|Lipase measurement|Lipase
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5211,5216|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5211,5216|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5211,5216|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5217,5222|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|SIMPLE_SEGMENT|5217,5222|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|SIMPLE_SEGMENT|5217,5222|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5217,5222|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5220,5224|false|false|false|C4722362|MB-6|MB-6
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5251,5256|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5251,5256|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5251,5256|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5251,5264|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5257,5264|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|5257,5264|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5257,5264|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5257,5264|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|5257,5264|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|5257,5264|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|5257,5264|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5257,5264|false|false|false|C0201925|Calcium measurement|Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5286,5290|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|5286,5290|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5286,5290|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Event|Event|SIMPLE_SEGMENT|5286,5290|false|false|false|||Iron
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5286,5290|false|false|false|C0337439|Iron measurement|Iron
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5307,5312|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5307,5312|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5307,5312|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|5337,5343|false|false|false|C0178638|folate|Folate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5337,5343|false|false|false|C0178638|folate|Folate
Drug|Vitamin|SIMPLE_SEGMENT|5337,5343|false|false|false|C0178638|folate|Folate
Event|Event|SIMPLE_SEGMENT|5337,5343|false|false|false|||Folate
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5337,5343|false|false|false|C0523631|Folic acid measurement|Folate
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5362,5365|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5362,5365|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Hormone|SIMPLE_SEGMENT|5362,5365|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5362,5365|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Event|Event|SIMPLE_SEGMENT|5362,5365|false|false|false|||TRF
Finding|Gene or Genome|SIMPLE_SEGMENT|5362,5365|false|false|false|C1334121;C1336604;C1705002|IL5 gene;TERF1 gene;TERF1 wt Allele|TRF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5383,5388|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5383,5388|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5383,5388|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5389,5392|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Enzyme|SIMPLE_SEGMENT|5389,5392|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Organic Chemical|SIMPLE_SEGMENT|5389,5392|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5389,5392|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Event|Event|SIMPLE_SEGMENT|5389,5392|false|false|false|||ASA
Finding|Gene or Genome|SIMPLE_SEGMENT|5389,5392|false|false|false|C1412553|ARSA gene|ASA
Event|Event|SIMPLE_SEGMENT|5393,5396|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|5393,5396|false|false|false|C5848551|Neg - answer|NEG
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|5397,5404|false|false|false|C0161679|Toxic effect of ethyl alcohol|Ethanol
Drug|Organic Chemical|SIMPLE_SEGMENT|5397,5404|false|false|false|C0001962;C3854029;C3854030|CNS depressants ethanol;antiseptics ethanol;ethanol|Ethanol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5397,5404|false|false|false|C0001962;C3854029;C3854030|CNS depressants ethanol;antiseptics ethanol;ethanol|Ethanol
Event|Event|SIMPLE_SEGMENT|5397,5404|false|false|false|||Ethanol
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5397,5404|false|false|false|C0202304|Ethanol measurement|Ethanol
Event|Event|SIMPLE_SEGMENT|5405,5408|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|5405,5408|false|false|false|C5848551|Neg - answer|NEG
Event|Event|SIMPLE_SEGMENT|5417,5420|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|5417,5420|false|false|false|C5848551|Neg - answer|NEG
Event|Event|SIMPLE_SEGMENT|5430,5433|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|5430,5433|false|false|false|C5848551|Neg - answer|NEG
Event|Event|SIMPLE_SEGMENT|5442,5445|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|5442,5445|false|false|false|C5848551|Neg - answer|NEG
Event|Event|SIMPLE_SEGMENT|5454,5457|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|5454,5457|false|false|false|C5848551|Neg - answer|NEG
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5470,5475|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5470,5475|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5470,5475|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Event|SIMPLE_SEGMENT|5476,5479|false|false|false|||pO2
Finding|Classification|SIMPLE_SEGMENT|5476,5479|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|pO2
Finding|Molecular Function|SIMPLE_SEGMENT|5476,5479|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|pO2
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5476,5479|false|false|false|C1283004|PO2 measurement|pO2
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5485,5489|false|false|false|C0391839|Carbon dioxide, partial pressure|pCO2
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5485,5489|false|false|false|C0201931|Carbon dioxide measurement, partial pressure|pCO2
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5515,5519|false|false|false|C2987514|Anatomical base|Base
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5515,5519|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|5515,5519|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|5515,5519|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Finding|Gene or Genome|SIMPLE_SEGMENT|5515,5519|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|Base
Finding|Idea or Concept|SIMPLE_SEGMENT|5515,5519|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|Base
Finding|Intellectual Product|SIMPLE_SEGMENT|5525,5532|false|false|false|C0282411;C0947611|Comment;Published Comment|Comment
Event|Event|SIMPLE_SEGMENT|5539,5542|false|false|false|||TOP
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5555,5560|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5555,5560|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5555,5560|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|5555,5568|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5555,5568|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5555,5568|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5561,5568|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|5561,5568|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5561,5568|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|5561,5568|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5561,5568|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5561,5568|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|5574,5581|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5574,5581|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5574,5581|false|false|false|C0202115|Lactic acid measurement|Lactate
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5619,5624|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5619,5624|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5619,5624|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5625,5628|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5625,5628|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|5625,5628|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5625,5628|false|false|false|C0019029|Hemoglobin concentration|Hgb
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5648,5651|false|false|false|C2744672|SAT1 protein, human|Sat
Drug|Enzyme|SIMPLE_SEGMENT|5648,5651|false|false|false|C2744672|SAT1 protein, human|Sat
Finding|Gene or Genome|SIMPLE_SEGMENT|5648,5651|false|false|false|C0871290;C1705827;C1822614|College Entrance Examination Board Scholastic Aptitude Test;SAT1 gene;SAT1 wt Allele|Sat
Finding|Intellectual Product|SIMPLE_SEGMENT|5648,5651|false|false|false|C0871290;C1705827;C1822614|College Entrance Examination Board Scholastic Aptitude Test;SAT1 gene;SAT1 wt Allele|Sat
Finding|Body Substance|SIMPLE_SEGMENT|5685,5690|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|5685,5690|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|5685,5690|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Finding|SIMPLE_SEGMENT|5685,5696|false|false|false|C0278030|Color of urine|URINE Color
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5691,5696|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|Color
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|5691,5696|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|Color
Event|Event|SIMPLE_SEGMENT|5735,5740|false|false|false|||URINE
Finding|Body Substance|SIMPLE_SEGMENT|5735,5740|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|5735,5740|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|5735,5740|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5735,5746|false|false|false|C0018965|Hematuria|URINE Blood
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5741,5746|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Finding|Body Substance|SIMPLE_SEGMENT|5741,5746|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5747,5750|false|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|MOD
Event|Event|SIMPLE_SEGMENT|5747,5750|false|false|false|||MOD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5751,5758|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5751,5758|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5751,5758|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5759,5762|false|false|false|C1744592|Structure of parieto-occipital fissure|POS
Finding|Intellectual Product|SIMPLE_SEGMENT|5759,5762|false|false|false|C5891108|Health Maintenance Organization Point of Service Plan|POS
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5763,5770|false|false|false|C0033684|Proteins|Protein
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5763,5770|false|false|false|C0033684|Proteins|Protein
Event|Event|SIMPLE_SEGMENT|5763,5770|false|false|false|||Protein
Finding|Conceptual Entity|SIMPLE_SEGMENT|5763,5770|false|false|false|C1521746|Protein Info|Protein
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5763,5770|false|false|false|C0202202|Protein measurement|Protein
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5776,5783|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|5776,5783|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5776,5783|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|5776,5783|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5776,5783|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5776,5783|false|false|false|C0337438|Glucose measurement|Glucose
Event|Event|SIMPLE_SEGMENT|5784,5787|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|5784,5787|false|false|false|C5848551|Neg - answer|NEG
Drug|Organic Chemical|SIMPLE_SEGMENT|5788,5794|false|false|false|C0022634|Ketones|Ketone
Event|Event|SIMPLE_SEGMENT|5795,5798|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|5795,5798|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|SIMPLE_SEGMENT|5807,5810|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|SIMPLE_SEGMENT|5819,5822|false|false|false|C5848551|Neg - answer|NEG
Event|Event|SIMPLE_SEGMENT|5851,5856|false|false|false|||URINE
Finding|Body Substance|SIMPLE_SEGMENT|5851,5856|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|5851,5856|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|5851,5856|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5851,5860|false|false|false|C0221752;C2188659|Red blood cells urine positive|URINE RBC
Anatomy|Cell|SIMPLE_SEGMENT|5857,5860|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5857,5860|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5857,5860|false|false|false|C0014792|Erythrocytes|RBC
Anatomy|Cell|SIMPLE_SEGMENT|5865,5868|false|false|false|C0023516|Leukocytes|WBC
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5882,5885|true|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|MOD
Event|Event|SIMPLE_SEGMENT|5882,5885|true|false|false|||MOD
Drug|Food|SIMPLE_SEGMENT|5886,5891|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Immunologic Factor|SIMPLE_SEGMENT|5886,5891|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|5886,5891|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5886,5891|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Event|Event|SIMPLE_SEGMENT|5892,5896|false|false|false|||NONE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5898,5901|true|false|false|C0267963|Exocrine pancreatic insufficiency|Epi
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5898,5901|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5898,5901|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Hormone|SIMPLE_SEGMENT|5898,5901|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Organic Chemical|SIMPLE_SEGMENT|5898,5901|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5898,5901|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Event|Event|SIMPLE_SEGMENT|5898,5901|true|false|false|||Epi
Finding|Gene or Genome|SIMPLE_SEGMENT|5898,5901|true|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|Epi
Finding|Intellectual Product|SIMPLE_SEGMENT|5898,5901|true|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|Epi
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5898,5901|true|false|false|C0162734;C3641909|Echo-Planar Imaging;Electronic Portal Imaging|Epi
Finding|Body Substance|SIMPLE_SEGMENT|5925,5930|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|5925,5930|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|5925,5930|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Body Substance|SIMPLE_SEGMENT|5953,5958|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|5953,5958|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|5953,5958|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Body Substance|SIMPLE_SEGMENT|5981,5986|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|5981,5986|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|5981,5986|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Finding|SIMPLE_SEGMENT|5981,5993|false|false|false|C0455910|Mucus in urine (finding)|URINE Mucous
Finding|Body Substance|SIMPLE_SEGMENT|5987,5993|false|false|false|C0026727;C2753459|Mucus (substance);mucus layer|Mucous
Event|Event|SIMPLE_SEGMENT|5994,5998|false|false|false|||RARE
Finding|Gene or Genome|SIMPLE_SEGMENT|5994,5998|false|false|false|C1514917|Retinoic Acid Response Element|RARE
Finding|Body Substance|SIMPLE_SEGMENT|6000,6009|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|6000,6009|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|6000,6009|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|6000,6009|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|SIMPLE_SEGMENT|6010,6014|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6010,6014|false|false|false|C0587081|Laboratory test finding|LABS
Event|Event|SIMPLE_SEGMENT|6022,6034|false|false|false|||MICROBIOLOGY
Finding|Functional Concept|SIMPLE_SEGMENT|6022,6034|false|false|false|C0025953;C1571921;C4049106|Microbiological;Microbiology - Laboratory Class;Microbiology Diagnostic Service Section ID|MICROBIOLOGY
Finding|Intellectual Product|SIMPLE_SEGMENT|6022,6034|false|false|false|C0025953;C1571921;C4049106|Microbiological;Microbiology - Laboratory Class;Microbiology Diagnostic Service Section ID|MICROBIOLOGY
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6022,6034|false|false|false|C0085672|Microbiology procedure|MICROBIOLOGY
Finding|Body Substance|SIMPLE_SEGMENT|6039,6044|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Functional Concept|SIMPLE_SEGMENT|6039,6044|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Intellectual Product|SIMPLE_SEGMENT|6039,6044|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6039,6052|false|false|false|C0430404|Urine culture|Urine culture
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6045,6052|false|false|false|C1706355|Culture Dose Form|culture
Event|Event|SIMPLE_SEGMENT|6045,6052|false|false|false|||culture
Finding|Functional Concept|SIMPLE_SEGMENT|6045,6052|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Finding|Idea or Concept|SIMPLE_SEGMENT|6045,6052|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6045,6052|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|culture
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6060,6071|false|false|false|C0033817|Pseudomonas Infections|PSEUDOMONAS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6060,6082|false|false|false|C0854135|Pseudomonas aeruginosa infection|PSEUDOMONAS AERUGINOSA
Event|Event|SIMPLE_SEGMENT|6072,6082|false|false|false|||AERUGINOSA
Event|Event|SIMPLE_SEGMENT|6110,6123|false|false|false|||SENSITIVITIES
Finding|Finding|SIMPLE_SEGMENT|6110,6123|false|false|false|C0427965|Antimicrobial susceptibility|SENSITIVITIES
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6125,6128|false|false|false|C2732473|Ductal Carcinoma In Situ with Microinvasion|MIC
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|6125,6128|false|false|false|C0066256|methyl isocyanate|MIC
Drug|Organic Chemical|SIMPLE_SEGMENT|6125,6128|false|false|false|C0066256|methyl isocyanate|MIC
Event|Event|SIMPLE_SEGMENT|6125,6128|false|false|false|||MIC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6125,6128|false|false|false|C0281162;C0427978|Minimum Inhibitory Concentration Test;cisplatin/ifosfamide/mitomycin protocol|MIC
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6125,6128|false|false|false|C0281162;C0427978|Minimum Inhibitory Concentration Test;cisplatin/ifosfamide/mitomycin protocol|MIC
Event|Event|SIMPLE_SEGMENT|6143,6146|false|false|false|||MCG
Drug|Antibiotic|SIMPLE_SEGMENT|6155,6163|false|false|false|C0002499|amikacin|AMIKACIN
Drug|Organic Chemical|SIMPLE_SEGMENT|6155,6163|false|false|false|C0002499|amikacin|AMIKACIN
Event|Event|SIMPLE_SEGMENT|6155,6163|false|false|false|||AMIKACIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6155,6163|false|false|false|C0002500|Amikacin measurement|AMIKACIN
Drug|Antibiotic|SIMPLE_SEGMENT|6191,6199|false|false|false|C0055003|cefepime|CEFEPIME
Drug|Organic Chemical|SIMPLE_SEGMENT|6191,6199|false|false|false|C0055003|cefepime|CEFEPIME
Drug|Antibiotic|SIMPLE_SEGMENT|6227,6238|false|false|false|C0007559|ceftazidime|CEFTAZIDIME
Drug|Organic Chemical|SIMPLE_SEGMENT|6227,6238|false|false|false|C0007559|ceftazidime|CEFTAZIDIME
Drug|Organic Chemical|SIMPLE_SEGMENT|6263,6276|false|false|false|C0008809|ciprofloxacin|CIPROFLOXACIN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6263,6276|false|false|false|C0008809|ciprofloxacin|CIPROFLOXACIN
Drug|Antibiotic|SIMPLE_SEGMENT|6299,6309|false|false|false|C3854019|gentamicin|GENTAMICIN
Drug|Organic Chemical|SIMPLE_SEGMENT|6299,6309|false|false|false|C3854019|gentamicin|GENTAMICIN
Event|Event|SIMPLE_SEGMENT|6299,6309|false|false|false|||GENTAMICIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6299,6309|false|false|false|C0202391|Gentamicin measurement|GENTAMICIN
Drug|Antibiotic|SIMPLE_SEGMENT|6335,6344|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|MEROPENEM
Drug|Clinical Drug|SIMPLE_SEGMENT|6335,6344|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|MEROPENEM
Drug|Organic Chemical|SIMPLE_SEGMENT|6335,6344|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|MEROPENEM
Drug|Antibiotic|SIMPLE_SEGMENT|6371,6383|false|false|false|C0031955|piperacillin|PIPERACILLIN
Drug|Organic Chemical|SIMPLE_SEGMENT|6371,6383|false|false|false|C0031955|piperacillin|PIPERACILLIN
Drug|Antibiotic|SIMPLE_SEGMENT|6384,6388|false|false|false|C0075870|tazobactam|TAZO
Drug|Organic Chemical|SIMPLE_SEGMENT|6384,6388|false|false|false|C0075870|tazobactam|TAZO
Drug|Antibiotic|SIMPLE_SEGMENT|6407,6417|false|false|false|C0040341|tobramycin|TOBRAMYCIN
Drug|Organic Chemical|SIMPLE_SEGMENT|6407,6417|false|false|false|C0040341|tobramycin|TOBRAMYCIN
Event|Event|SIMPLE_SEGMENT|6407,6417|false|false|false|||TOBRAMYCIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6407,6417|false|false|false|C0202490|Tobramycin measurement|TOBRAMYCIN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6440,6445|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Event|Event|SIMPLE_SEGMENT|6440,6445|false|false|false|||Blood
Finding|Body Substance|SIMPLE_SEGMENT|6440,6445|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6440,6453|false|false|false|C0200949|Blood culture|Blood culture
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6446,6453|false|false|false|C1706355|Culture Dose Form|culture
Event|Event|SIMPLE_SEGMENT|6446,6453|false|false|false|||culture
Finding|Functional Concept|SIMPLE_SEGMENT|6446,6453|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Finding|Idea or Concept|SIMPLE_SEGMENT|6446,6453|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6446,6453|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|culture
Event|Event|SIMPLE_SEGMENT|6475,6482|false|false|false|||SPECIES
Finding|Classification|SIMPLE_SEGMENT|6475,6482|false|false|false|C1548151;C1705920|Species;Species - Nature of Abnormal Testing|SPECIES
Finding|Idea or Concept|SIMPLE_SEGMENT|6475,6482|false|false|false|C1548151;C1705920|Species;Species - Nature of Abnormal Testing|SPECIES
Event|Event|SIMPLE_SEGMENT|6484,6492|false|false|false|||Isolated
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6508,6511|false|false|false|C1137947|SET protein, human|set
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6508,6511|false|false|false|C1137947|SET protein, human|set
Event|Event|SIMPLE_SEGMENT|6508,6511|false|false|false|||set
Finding|Conceptual Entity|SIMPLE_SEGMENT|6508,6511|false|false|false|C0036849;C1366517;C1442518;C1552652;C1705195|Parameterized Data Type - Set;SET gene;Set (Psychology);Set scale;set (group)|set
Finding|Functional Concept|SIMPLE_SEGMENT|6508,6511|false|false|false|C0036849;C1366517;C1442518;C1552652;C1705195|Parameterized Data Type - Set;SET gene;Set (Psychology);Set scale;set (group)|set
Finding|Gene or Genome|SIMPLE_SEGMENT|6508,6511|false|false|false|C0036849;C1366517;C1442518;C1552652;C1705195|Parameterized Data Type - Set;SET gene;Set (Psychology);Set scale;set (group)|set
Finding|Idea or Concept|SIMPLE_SEGMENT|6508,6511|false|false|false|C0036849;C1366517;C1442518;C1552652;C1705195|Parameterized Data Type - Set;SET gene;Set (Psychology);Set scale;set (group)|set
Finding|Mental Process|SIMPLE_SEGMENT|6508,6511|false|false|false|C0036849;C1366517;C1442518;C1552652;C1705195|Parameterized Data Type - Set;SET gene;Set (Psychology);Set scale;set (group)|set
Event|Event|SIMPLE_SEGMENT|6541,6554|false|false|false|||SENSITIVITIES
Finding|Finding|SIMPLE_SEGMENT|6541,6554|false|false|false|C0427965|Antimicrobial susceptibility|SENSITIVITIES
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6556,6559|false|false|false|C2732473|Ductal Carcinoma In Situ with Microinvasion|MIC
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|6556,6559|false|false|false|C0066256|methyl isocyanate|MIC
Drug|Organic Chemical|SIMPLE_SEGMENT|6556,6559|false|false|false|C0066256|methyl isocyanate|MIC
Event|Event|SIMPLE_SEGMENT|6556,6559|false|false|false|||MIC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6556,6559|false|false|false|C0281162;C0427978|Minimum Inhibitory Concentration Test;cisplatin/ifosfamide/mitomycin protocol|MIC
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6556,6559|false|false|false|C0281162;C0427978|Minimum Inhibitory Concentration Test;cisplatin/ifosfamide/mitomycin protocol|MIC
Event|Event|SIMPLE_SEGMENT|6574,6577|false|false|false|||MCG
Drug|Antibiotic|SIMPLE_SEGMENT|6586,6596|false|false|false|C0002680;C2095775|ampicillin;ampicillins|AMPICILLIN
Drug|Organic Chemical|SIMPLE_SEGMENT|6586,6596|false|false|false|C0002680;C2095775|ampicillin;ampicillins|AMPICILLIN
Drug|Antibiotic|SIMPLE_SEGMENT|6622,6632|false|false|false|C3854019|gentamicin|GENTAMICIN
Drug|Organic Chemical|SIMPLE_SEGMENT|6622,6632|false|false|false|C3854019|gentamicin|GENTAMICIN
Event|Event|SIMPLE_SEGMENT|6622,6632|false|false|false|||GENTAMICIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6622,6632|false|false|false|C0202391|Gentamicin measurement|GENTAMICIN
Drug|Antibiotic|SIMPLE_SEGMENT|6658,6668|false|false|false|C0030842|penicillins|PENICILLIN
Drug|Organic Chemical|SIMPLE_SEGMENT|6658,6668|false|false|false|C0030842|penicillins|PENICILLIN
Drug|Antibiotic|SIMPLE_SEGMENT|6658,6670|false|false|false|C0030827|penicillin G|PENICILLIN G
Drug|Organic Chemical|SIMPLE_SEGMENT|6658,6670|false|false|false|C0030827|penicillin G|PENICILLIN G
Finding|Body Substance|SIMPLE_SEGMENT|6691,6697|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|Sputum
Finding|Intellectual Product|SIMPLE_SEGMENT|6691,6697|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|Sputum
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6691,6705|false|false|false|C0523174|Microbial culture of sputum|Sputum culture
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6698,6705|false|false|false|C1706355|Culture Dose Form|culture
Event|Event|SIMPLE_SEGMENT|6698,6705|false|false|false|||culture
Finding|Functional Concept|SIMPLE_SEGMENT|6698,6705|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Finding|Idea or Concept|SIMPLE_SEGMENT|6698,6705|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6698,6705|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|culture
Event|Event|SIMPLE_SEGMENT|6724,6730|false|false|false|||source
Finding|Finding|SIMPLE_SEGMENT|6724,6730|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Functional Concept|SIMPLE_SEGMENT|6724,6730|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Intellectual Product|SIMPLE_SEGMENT|6724,6730|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Event|Event|SIMPLE_SEGMENT|6737,6741|false|false|false|||GRAM
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|6737,6747|false|false|false|C0061856|Gram's stain|GRAM STAIN
Drug|Organic Chemical|SIMPLE_SEGMENT|6737,6747|false|false|false|C0061856|Gram's stain|GRAM STAIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6737,6747|false|false|false|C0200966|Bacterial stain, routine|GRAM STAIN
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|6742,6747|false|false|false|C0038128|Stains|STAIN
Event|Event|SIMPLE_SEGMENT|6742,6747|false|false|false|||STAIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6742,6747|false|false|false|C0487602|Staining method|STAIN
Anatomy|Cell|SIMPLE_SEGMENT|6766,6782|false|false|false|C0014597|Epithelial Cells|epithelial cells
Anatomy|Cell|SIMPLE_SEGMENT|6777,6782|false|false|false|C0007634|Cells|cells
Event|Event|SIMPLE_SEGMENT|6788,6793|false|false|false|||field
Finding|Conceptual Entity|SIMPLE_SEGMENT|6788,6793|false|false|false|C1521738;C2346620;C2349184|Field;Force Field;Knowledge Field|field
Procedure|Health Care Activity|SIMPLE_SEGMENT|6788,6793|false|false|false|C1553496|field - patient encounter|field
Event|Event|SIMPLE_SEGMENT|6821,6826|false|false|false|||FIELD
Finding|Conceptual Entity|SIMPLE_SEGMENT|6821,6826|false|false|false|C1521738;C2346620;C2349184|Field;Force Field;Knowledge Field|FIELD
Procedure|Health Care Activity|SIMPLE_SEGMENT|6821,6826|false|false|false|C1553496|field - patient encounter|FIELD
Event|Event|SIMPLE_SEGMENT|6831,6838|false|false|false|||BUDDING
Finding|Cell Function|SIMPLE_SEGMENT|6831,6838|false|false|false|C1155616|Cell budding|BUDDING
Drug|Food|SIMPLE_SEGMENT|6839,6844|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Immunologic Factor|SIMPLE_SEGMENT|6839,6844|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|6839,6844|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6839,6844|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Event|Event|SIMPLE_SEGMENT|6839,6844|false|false|false|||YEAST
Event|Event|SIMPLE_SEGMENT|6851,6863|false|false|false|||PSEUDOHYPHAE
Event|Event|SIMPLE_SEGMENT|6892,6897|false|false|false|||FIELD
Finding|Conceptual Entity|SIMPLE_SEGMENT|6892,6897|false|false|false|C1521738;C2346620;C2349184|Field;Force Field;Knowledge Field|FIELD
Procedure|Health Care Activity|SIMPLE_SEGMENT|6892,6897|false|false|false|C1553496|field - patient encounter|FIELD
Event|Event|SIMPLE_SEGMENT|6902,6906|false|false|false|||GRAM
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|6907,6915|false|false|false|C4727483|BRAF Gene Rearrangement|POSITIVE
Event|Event|SIMPLE_SEGMENT|6907,6915|false|false|false|||POSITIVE
Finding|Classification|SIMPLE_SEGMENT|6907,6915|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|POSITIVE
Finding|Finding|SIMPLE_SEGMENT|6907,6915|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|POSITIVE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6986,6997|false|false|false|C0231832|Respiratory rate|RESPIRATORY
Finding|Body Substance|SIMPLE_SEGMENT|6986,6997|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|RESPIRATORY
Finding|Functional Concept|SIMPLE_SEGMENT|6986,6997|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|RESPIRATORY
Finding|Intellectual Product|SIMPLE_SEGMENT|6986,6997|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|RESPIRATORY
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6986,7005|false|false|false|C4282127|Respiratory culture|RESPIRATORY CULTURE
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6998,7005|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|SIMPLE_SEGMENT|6998,7005|false|false|false|||CULTURE
Finding|Functional Concept|SIMPLE_SEGMENT|6998,7005|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|6998,7005|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6998,7005|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|7007,7012|false|false|false|C1546485|Diagnosis Type - Final|Final
Finding|Finding|SIMPLE_SEGMENT|7025,7033|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|MODERATE
Finding|Intellectual Product|SIMPLE_SEGMENT|7025,7033|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|MODERATE
Event|Event|SIMPLE_SEGMENT|7034,7040|false|false|false|||GROWTH
Finding|Finding|SIMPLE_SEGMENT|7034,7040|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|7034,7040|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organism Function|SIMPLE_SEGMENT|7034,7040|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Physiologic Function|SIMPLE_SEGMENT|7034,7040|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|7034,7040|false|false|false|C2911660|Growth action|GROWTH
Finding|Functional Concept|SIMPLE_SEGMENT|7041,7050|false|false|false|C0231202|Symbiotic|Commensal
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7051,7062|false|false|false|C0231832|Respiratory rate|Respiratory
Finding|Body Substance|SIMPLE_SEGMENT|7051,7062|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|Respiratory
Finding|Functional Concept|SIMPLE_SEGMENT|7051,7062|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|Respiratory
Finding|Intellectual Product|SIMPLE_SEGMENT|7051,7062|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|Respiratory
Drug|Food|SIMPLE_SEGMENT|7077,7082|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Immunologic Factor|SIMPLE_SEGMENT|7077,7082|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|7077,7082|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7077,7082|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Event|Event|SIMPLE_SEGMENT|7077,7082|false|false|false|||YEAST
Event|Event|SIMPLE_SEGMENT|7091,7097|false|false|false|||GROWTH
Finding|Finding|SIMPLE_SEGMENT|7091,7097|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|7091,7097|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organism Function|SIMPLE_SEGMENT|7091,7097|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Physiologic Function|SIMPLE_SEGMENT|7091,7097|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|7091,7097|false|false|false|C2911660|Growth action|GROWTH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7103,7121|false|false|false|C1294227|Legionella culture|LEGIONELLA CULTURE
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7114,7121|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|SIMPLE_SEGMENT|7114,7121|false|false|false|||CULTURE
Finding|Functional Concept|SIMPLE_SEGMENT|7114,7121|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|7114,7121|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7114,7121|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|SIMPLE_SEGMENT|7143,7153|true|false|false|||LEGIONELLA
Event|Event|SIMPLE_SEGMENT|7154,7162|true|false|false|||ISOLATED
Finding|Body Substance|SIMPLE_SEGMENT|7167,7172|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Functional Concept|SIMPLE_SEGMENT|7167,7172|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Intellectual Product|SIMPLE_SEGMENT|7167,7172|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7167,7180|false|false|false|C0430404|Urine culture|Urine culture
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7173,7180|false|false|false|C1706355|Culture Dose Form|culture
Event|Event|SIMPLE_SEGMENT|7173,7180|false|false|false|||culture
Finding|Functional Concept|SIMPLE_SEGMENT|7173,7180|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Finding|Idea or Concept|SIMPLE_SEGMENT|7173,7180|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7173,7180|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|culture
Drug|Food|SIMPLE_SEGMENT|7194,7199|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Immunologic Factor|SIMPLE_SEGMENT|7194,7199|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|7194,7199|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7194,7199|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Event|Event|SIMPLE_SEGMENT|7194,7199|false|false|false|||YEAST
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7233,7238|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Event|Event|SIMPLE_SEGMENT|7233,7238|false|false|false|||Blood
Finding|Body Substance|SIMPLE_SEGMENT|7233,7238|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7233,7246|false|false|false|C0200949|Blood culture|Blood culture
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7239,7246|false|false|false|C1706355|Culture Dose Form|culture
Event|Event|SIMPLE_SEGMENT|7239,7246|false|false|false|||culture
Finding|Functional Concept|SIMPLE_SEGMENT|7239,7246|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Finding|Idea or Concept|SIMPLE_SEGMENT|7239,7246|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7239,7246|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|culture
Finding|Idea or Concept|SIMPLE_SEGMENT|7252,7257|false|false|false|C1546485|Diagnosis Type - Final|final
Finding|Classification|SIMPLE_SEGMENT|7260,7268|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Finding|Finding|SIMPLE_SEGMENT|7260,7268|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7260,7268|false|false|false|C5237010|Expression Negative|NEGATIVE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7270,7275|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Event|Event|SIMPLE_SEGMENT|7270,7275|false|false|false|||Blood
Finding|Body Substance|SIMPLE_SEGMENT|7270,7275|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7270,7283|false|false|false|C0200949|Blood culture|Blood culture
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7276,7283|false|false|false|C1706355|Culture Dose Form|culture
Event|Event|SIMPLE_SEGMENT|7276,7283|false|false|false|||culture
Finding|Functional Concept|SIMPLE_SEGMENT|7276,7283|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Finding|Idea or Concept|SIMPLE_SEGMENT|7276,7283|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7276,7283|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|culture
Finding|Idea or Concept|SIMPLE_SEGMENT|7289,7294|false|false|false|C1546485|Diagnosis Type - Final|final
Finding|Classification|SIMPLE_SEGMENT|7297,7305|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Finding|Finding|SIMPLE_SEGMENT|7297,7305|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7297,7305|false|false|false|C5237010|Expression Negative|NEGATIVE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7307,7312|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Event|Event|SIMPLE_SEGMENT|7307,7312|false|false|false|||Blood
Finding|Body Substance|SIMPLE_SEGMENT|7307,7312|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7307,7320|false|false|false|C0200949|Blood culture|Blood culture
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7313,7320|false|false|false|C1706355|Culture Dose Form|culture
Event|Event|SIMPLE_SEGMENT|7313,7320|false|false|false|||culture
Finding|Functional Concept|SIMPLE_SEGMENT|7313,7320|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Finding|Idea or Concept|SIMPLE_SEGMENT|7313,7320|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7313,7320|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|culture
Event|Event|SIMPLE_SEGMENT|7326,7333|false|false|false|||pending
Finding|Idea or Concept|SIMPLE_SEGMENT|7326,7333|false|false|false|C1691786;C1704475|Pending - Allergy Clinical Status;Pending - referral status|pending
Event|Event|SIMPLE_SEGMENT|7339,7345|true|false|false|||GROWTH
Finding|Finding|SIMPLE_SEGMENT|7339,7345|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|7339,7345|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organism Function|SIMPLE_SEGMENT|7339,7345|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Physiologic Function|SIMPLE_SEGMENT|7339,7345|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|7339,7345|true|false|false|C2911660|Growth action|GROWTH
Event|Event|SIMPLE_SEGMENT|7349,7353|true|false|false|||DATE
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7359,7364|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|CHEST
Finding|Finding|SIMPLE_SEGMENT|7359,7364|true|false|false|C0741025|Chest problem|CHEST
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7359,7370|true|false|false|C0039985|Plain chest X-ray|CHEST X-RAY
Event|Event|SIMPLE_SEGMENT|7365,7370|false|false|false|||X-RAY
Finding|Functional Concept|SIMPLE_SEGMENT|7365,7370|false|false|false|C0034571;C3244296|ActClaimAttachmentCategoryCode - x-ray;roentgenographic|X-RAY
Finding|Intellectual Product|SIMPLE_SEGMENT|7365,7370|false|false|false|C0034571;C3244296|ActClaimAttachmentCategoryCode - x-ray;roentgenographic|X-RAY
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|7365,7370|false|false|false|C0043309|Roentgen Rays|X-RAY
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7365,7370|false|false|false|C0043299;C1306645;C1962945|Diagnostic radiologic examination;Plain x-ray;Radiographic imaging procedure|X-RAY
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7382,7408|false|false|false|C0747635|Bilateral pleural effusion|Bilateral pleural effusion
Anatomy|Tissue|SIMPLE_SEGMENT|7392,7399|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7392,7399|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Body Substance|SIMPLE_SEGMENT|7392,7408|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Finding|SIMPLE_SEGMENT|7392,7408|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|7392,7408|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Event|Event|SIMPLE_SEGMENT|7400,7408|false|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|7400,7408|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|7400,7408|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|7400,7408|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Event|Event|SIMPLE_SEGMENT|7410,7415|false|false|false|||right
Finding|Functional Concept|SIMPLE_SEGMENT|7410,7415|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Event|Event|SIMPLE_SEGMENT|7429,7433|false|false|false|||left
Finding|Functional Concept|SIMPLE_SEGMENT|7429,7433|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Finding|SIMPLE_SEGMENT|7436,7446|true|false|false|C4722602|Underlying|Underlying
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7448,7461|true|false|false|C0521530|Lung consolidation|consolidation
Event|Event|SIMPLE_SEGMENT|7448,7461|true|false|false|||consolidation
Finding|Intellectual Product|SIMPLE_SEGMENT|7472,7482|true|true|false|C4554154|Completely - dosing instruction fragment|completely
Event|Event|SIMPLE_SEGMENT|7483,7491|true|false|false|||excluded
Event|Event|SIMPLE_SEGMENT|7510,7514|false|false|false|||tube
Finding|Functional Concept|SIMPLE_SEGMENT|7510,7514|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Finding|Gene or Genome|SIMPLE_SEGMENT|7510,7514|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Event|Event|SIMPLE_SEGMENT|7515,7525|false|false|false|||terminates
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7543,7549|false|false|false|C0225594;C4521147|Keel structure;Structure of carina|carina
Event|Event|SIMPLE_SEGMENT|7552,7561|false|false|false|||Recommend
Finding|Idea or Concept|SIMPLE_SEGMENT|7552,7561|false|false|false|C0034866|Recommendation|Recommend
Event|Event|SIMPLE_SEGMENT|7563,7576|false|false|false|||repositioning
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7563,7576|false|false|false|C0556030|Repositioning (procedure)|repositioning
Event|Event|SIMPLE_SEGMENT|7585,7589|false|false|false|||tube
Finding|Functional Concept|SIMPLE_SEGMENT|7585,7589|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Finding|Gene or Genome|SIMPLE_SEGMENT|7585,7589|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Event|Event|SIMPLE_SEGMENT|7590,7600|false|false|false|||terminates
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7605,7612|false|false|false|C0038351;C3714551;C4266636|Abdomen>Stomach;Stomach;Stomach structure|stomach
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7605,7612|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7605,7612|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Event|Event|SIMPLE_SEGMENT|7605,7612|false|false|false|||stomach
Finding|Finding|SIMPLE_SEGMENT|7605,7612|false|false|false|C0577027|Stomach problem|stomach
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7605,7612|false|false|false|C0872393|Procedure on stomach|stomach
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7631,7637|false|false|false|C4522154|Distal Resection Margin|distal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7639,7648|false|false|false|C0014876;C4266613|Chest>Esophagus;Esophagus|esophagus
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7639,7648|false|false|false|C0014852;C0153942;C0154059|Benign neoplasm of esophagus;Carcinoma in situ of esophagus;Esophageal Diseases|esophagus
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7639,7648|false|false|false|C0014852;C0153942;C0154059|Benign neoplasm of esophagus;Carcinoma in situ of esophagus;Esophageal Diseases|esophagus
Event|Event|SIMPLE_SEGMENT|7639,7648|false|false|false|||esophagus
Finding|Finding|SIMPLE_SEGMENT|7639,7648|false|false|false|C0812418|Esophagus problem|esophagus
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7639,7648|false|false|false|C0872395|Procedures on the esophagus|esophagus
Finding|Functional Concept|SIMPLE_SEGMENT|7654,7659|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Event|Event|SIMPLE_SEGMENT|7660,7664|false|false|false|||PICC
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7660,7664|false|false|false|C2049629|Peripherally Inserted Central Catheter Line Insertion|PICC
Event|Event|SIMPLE_SEGMENT|7665,7675|false|false|false|||terminates
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7684,7690|false|false|false|C0004454|Axilla|axilla
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7694,7701|true|false|false|C0881943||CT HEAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7694,7701|true|false|false|C0202691|CAT scan of head|CT HEAD
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7697,7701|true|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|HEAD
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7697,7701|true|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|HEAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7697,7701|true|false|false|C0362076|Problems with head|HEAD
Event|Event|SIMPLE_SEGMENT|7697,7701|true|false|false|||HEAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7697,7701|true|false|false|C0876917|Procedure on head|HEAD
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|7710,7718|true|false|false|C0009924|Contrast Media|CONTRAST
Event|Event|SIMPLE_SEGMENT|7710,7718|true|false|false|||CONTRAST
Event|Event|SIMPLE_SEGMENT|7738,7746|true|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|7738,7746|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|7738,7749|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Event|Event|SIMPLE_SEGMENT|7751,7761|true|false|false|||hemorrhage
Finding|Pathologic Function|SIMPLE_SEGMENT|7751,7761|true|false|false|C0019080|Hemorrhage|hemorrhage
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7763,7768|true|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|7763,7768|true|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|7763,7768|true|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|7770,7780|false|false|false|||infarction
Finding|Pathologic Function|SIMPLE_SEGMENT|7770,7780|false|false|false|C0021308|Infarction|infarction
Event|Event|SIMPLE_SEGMENT|7785,7789|false|false|false|||mass
Finding|Finding|SIMPLE_SEGMENT|7785,7789|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|SIMPLE_SEGMENT|7785,7789|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|SIMPLE_SEGMENT|7785,7789|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Finding|SIMPLE_SEGMENT|7785,7796|false|false|false|C4086564|Mass Effect|mass effect
Event|Event|SIMPLE_SEGMENT|7790,7796|false|false|false|||effect
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7802,7812|false|false|false|C0018827|Heart Ventricle|ventricles
Event|Event|SIMPLE_SEGMENT|7818,7823|false|false|false|||sulci
Event|Event|SIMPLE_SEGMENT|7828,7837|false|false|false|||prominent
Event|Event|SIMPLE_SEGMENT|7839,7849|false|false|false|||suggesting
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7850,7853|false|false|false|C1114365||age
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7850,7853|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|SIMPLE_SEGMENT|7850,7853|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|SIMPLE_SEGMENT|7854,7861|false|false|false|C0163712|Relate - vinyl resin|related
Finding|Finding|SIMPLE_SEGMENT|7854,7861|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|SIMPLE_SEGMENT|7854,7861|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Event|Event|SIMPLE_SEGMENT|7862,7874|false|false|false|||involutional
Event|Event|SIMPLE_SEGMENT|7876,7883|false|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|7876,7883|false|false|false|C0392747|Changing|changes
Event|Event|SIMPLE_SEGMENT|7887,7894|false|false|false|||atrophy
Finding|Pathologic Function|SIMPLE_SEGMENT|7887,7894|false|false|false|C0333641|Atrophic|atrophy
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7896,7924|false|false|false|C0228157|Periventricular white matter|Periventricular white matter
Finding|Finding|SIMPLE_SEGMENT|7896,7938|false|false|false|C4022720|Periventricular white matter hypodensities|Periventricular white matter hypodensities
Anatomy|Tissue|SIMPLE_SEGMENT|7912,7924|false|false|false|C0682708|White matter|white matter
Event|Event|SIMPLE_SEGMENT|7925,7938|false|false|false|||hypodensities
Event|Event|SIMPLE_SEGMENT|7944,7954|false|false|false|||compatible
Finding|Idea or Concept|SIMPLE_SEGMENT|7944,7954|false|false|false|C0332290|Consistent with|compatible
Finding|Idea or Concept|SIMPLE_SEGMENT|7944,7959|false|false|false|C0332290|Consistent with|compatible with
Event|Event|SIMPLE_SEGMENT|7960,7967|false|false|false|||chronic
Finding|Intellectual Product|SIMPLE_SEGMENT|7960,7967|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|7960,7967|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7968,7980|false|false|false|C0225988|Structure of small blood vessel (organ)|small vessel
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7974,7980|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7974,7980|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Finding|Functional Concept|SIMPLE_SEGMENT|7981,7989|false|false|false|C0475224|Ischemic|ischemic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7990,7997|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|7990,7997|false|false|false|||disease
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|8006,8014|false|false|false|C1185718|Cistern|cisterns
Event|Event|SIMPLE_SEGMENT|8022,8028|false|false|false|||patent
Finding|Intellectual Product|SIMPLE_SEGMENT|8022,8028|false|false|false|C0030650|Legal patent|patent
Event|Event|SIMPLE_SEGMENT|8043,8055|false|false|false|||preservation
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8043,8055|false|false|false|C0033085;C1514402|Biologic Preservation;Preservation Technique|preservation
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8078,8093|false|false|false|C1511938|Cellular Differentiation Qualifier|differentiation
Event|Event|SIMPLE_SEGMENT|8078,8093|false|false|false|||differentiation
Finding|Cell Function|SIMPLE_SEGMENT|8078,8093|false|false|false|C0007589;C2945687|Cell Differentiation process;Differentiation|differentiation
Finding|Functional Concept|SIMPLE_SEGMENT|8078,8093|false|false|false|C0007589;C2945687|Cell Differentiation process;Differentiation|differentiation
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|8098,8106|true|false|false|C0016658|Fracture|fracture
Event|Event|SIMPLE_SEGMENT|8098,8106|true|false|false|||fracture
Event|Event|SIMPLE_SEGMENT|8110,8120|true|false|false|||identified
Drug|Substance|SIMPLE_SEGMENT|8132,8137|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|8132,8137|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|8132,8137|false|false|false|C1546638|Fluid Specimen Code|fluid
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8149,8154|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8149,8154|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|SIMPLE_SEGMENT|8149,8154|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8149,8154|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|SIMPLE_SEGMENT|8149,8154|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|SIMPLE_SEGMENT|8149,8154|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|8149,8161|false|false|false|C0027423|Nasal cavity|nasal cavity
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8149,8161|false|false|false|C0728864|Malignant neoplasm of nasal cavity|nasal cavity
Procedure|Health Care Activity|SIMPLE_SEGMENT|8149,8161|false|false|false|C2087464|examination of nasal cavity|nasal cavity
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|8155,8161|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|8155,8161|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8155,8161|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Event|Event|SIMPLE_SEGMENT|8155,8161|false|false|false|||cavity
Finding|Finding|SIMPLE_SEGMENT|8163,8169|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|8163,8169|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8170,8179|false|false|false|C0027627|Neoplasm Metastasis|secondary
Event|Event|SIMPLE_SEGMENT|8170,8179|false|false|false|||secondary
Finding|Functional Concept|SIMPLE_SEGMENT|8170,8179|false|false|false|C1522484|metastatic qualifier|secondary
Event|Event|SIMPLE_SEGMENT|8183,8192|false|false|false|||intubated
Finding|Finding|SIMPLE_SEGMENT|8183,8192|false|false|false|C4698386|Intubated|intubated
Event|Event|SIMPLE_SEGMENT|8194,8199|false|false|false|||state
Finding|Functional Concept|SIMPLE_SEGMENT|8194,8199|false|false|false|C1442792|State|state
Finding|Functional Concept|SIMPLE_SEGMENT|8202,8217|false|false|false|C0333482|atherosclerotic|Atherosclerotic
Event|Event|SIMPLE_SEGMENT|8224,8238|false|false|false|||calcifications
Finding|Finding|SIMPLE_SEGMENT|8224,8238|false|false|false|C0006660;C2242558|Pathologic calcification, calcified structure;Physiologic calcification|calcifications
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|8224,8238|false|false|false|C0006660;C2242558|Pathologic calcification, calcified structure;Physiologic calcification|calcifications
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8256,8263|false|false|false|C0007272|Carotid Arteries|carotid
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8256,8272|false|false|false|C0007272;C4071877|Carotid Arteries;Head+Neck>Carotid artery|carotid arteries
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8264,8272|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Anatomy|Body System|SIMPLE_SEGMENT|8264,8272|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Event|Event|SIMPLE_SEGMENT|8264,8272|false|false|false|||arteries
Procedure|Health Care Activity|SIMPLE_SEGMENT|8264,8272|false|false|false|C0397581|Procedure on artery|arteries
Event|Event|SIMPLE_SEGMENT|8277,8284|false|false|false|||present
Finding|Finding|SIMPLE_SEGMENT|8277,8284|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|SIMPLE_SEGMENT|8277,8284|false|false|false|C0150312;C0449450|Present;Presentation|present
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|8301,8318|false|false|false|C0030471|Nasal sinus|paranasal sinuses
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|8311,8318|false|false|false|C0030471;C4071871|Head>Sinuses;Nasal sinus|sinuses
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|8311,8318|false|false|false|C0016169|pathologic fistula|sinuses
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8321,8328|false|false|false|C0446908;C1521748;C4266570|Head>Mastoid;Mastoid process|mastoid
Procedure|Health Care Activity|SIMPLE_SEGMENT|8321,8328|false|false|false|C2228459|examination of mastoid region|mastoid
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|8321,8338|false|false|false|C0229427|Pneumatic mastoid cell|mastoid air cells
Drug|Inorganic Chemical|SIMPLE_SEGMENT|8329,8332|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8329,8332|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|SIMPLE_SEGMENT|8329,8332|false|false|false|C0001861;C3536832|Air (substance);air|air
Finding|Finding|SIMPLE_SEGMENT|8329,8332|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|SIMPLE_SEGMENT|8329,8332|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|SIMPLE_SEGMENT|8329,8332|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Anatomy|Cell|SIMPLE_SEGMENT|8333,8338|false|false|false|C0007634|Cells|cells
Finding|Intellectual Product|SIMPLE_SEGMENT|8344,8350|false|false|false|C1552826|Table Cell Vertical Align - middle|middle
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|8344,8354|false|false|false|C0013455|middle ear|middle ear
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8344,8354|false|false|false|C0271428;C0496788|Disorder of middle ear;Malignant neoplasm of middle ear|middle ear
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8344,8354|false|false|false|C0271428;C0496788|Disorder of middle ear;Malignant neoplasm of middle ear|middle ear
Procedure|Health Care Activity|SIMPLE_SEGMENT|8344,8354|false|false|false|C2228461|examination of middle ear|middle ear
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8351,8354|false|false|false|C0013443;C0521421|Ear structure|ear
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8351,8354|false|false|false|C0851354|Ear and labyrinth disorders|ear
Finding|Body Substance|SIMPLE_SEGMENT|8351,8354|false|false|false|C1546608;C1550629|SpecimenType - Ear|ear
Finding|Intellectual Product|SIMPLE_SEGMENT|8351,8354|false|false|false|C1546608;C1550629|SpecimenType - Ear|ear
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|8355,8363|false|false|false|C0333343|Body cavities|cavities
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|8355,8363|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavities
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8355,8363|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavities
Event|Event|SIMPLE_SEGMENT|8355,8363|false|false|false|||cavities
Event|Event|SIMPLE_SEGMENT|8378,8383|false|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|8378,8383|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8396,8402|false|false|false|C0015392;C0700042|Eye;Orbital region|ocular
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8396,8402|false|false|false|C0015392;C0700042|Eye;Orbital region|ocular
Finding|Finding|SIMPLE_SEGMENT|8396,8402|false|false|false|C0042789;C1299003;C4521296|Ocular (intended site);Ocular (qualifier);Vision|ocular
Finding|Functional Concept|SIMPLE_SEGMENT|8396,8402|false|false|false|C0042789;C1299003;C4521296|Ocular (intended site);Ocular (qualifier);Vision|ocular
Finding|Organism Function|SIMPLE_SEGMENT|8396,8402|false|false|false|C0042789;C1299003;C4521296|Ocular (intended site);Ocular (qualifier);Vision|ocular
Event|Event|SIMPLE_SEGMENT|8403,8409|false|false|false|||lenses
Event|Event|SIMPLE_SEGMENT|8420,8428|false|false|false|||replaced
Event|Event|SIMPLE_SEGMENT|8430,8440|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|8430,8440|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|8430,8440|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8446,8458|true|false|false|C0524466|Intracranial|intracranial
Finding|Functional Concept|SIMPLE_SEGMENT|8446,8458|true|false|false|C1522213|Intracranial Route of Administration|intracranial
Finding|Pathologic Function|SIMPLE_SEGMENT|8446,8469|true|false|false|C0151699|Intracranial Hemorrhage|intracranial hemorrhage
Event|Event|SIMPLE_SEGMENT|8459,8469|true|false|false|||hemorrhage
Finding|Pathologic Function|SIMPLE_SEGMENT|8459,8469|true|false|false|C0019080|Hemorrhage|hemorrhage
Event|Event|SIMPLE_SEGMENT|8473,8477|true|false|false|||mass
Finding|Finding|SIMPLE_SEGMENT|8473,8477|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|SIMPLE_SEGMENT|8473,8477|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|SIMPLE_SEGMENT|8473,8477|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Finding|SIMPLE_SEGMENT|8473,8484|true|false|false|C4086564|Mass Effect|mass effect
Event|Event|SIMPLE_SEGMENT|8478,8484|true|false|false|||effect
Event|Event|SIMPLE_SEGMENT|8488,8491|false|false|false|||TTE
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8488,8491|false|false|false|C0430462|Transthoracic echocardiography|TTE
Finding|Functional Concept|SIMPLE_SEGMENT|8503,8507|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8503,8514|false|false|false|C0225860|Left atrial structure|left atrium
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8508,8514|false|false|false|C0018792|Heart Atrium|atrium
Event|Event|SIMPLE_SEGMENT|8518,8524|false|false|false|||normal
Finding|Intellectual Product|SIMPLE_SEGMENT|8544,8548|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Pathologic Function|SIMPLE_SEGMENT|8568,8585|false|false|false|C1280751|Focal hypertrophy|focal hypertrophy
Event|Event|SIMPLE_SEGMENT|8574,8585|false|false|false|||hypertrophy
Finding|Pathologic Function|SIMPLE_SEGMENT|8574,8585|false|false|false|C0020564|Hypertrophy|hypertrophy
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|8599,8605|false|false|false|C0936188;C1327729;C2362924|Cell septum;Septum - general anatomical term;Septum of telencephalon|septum
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8599,8605|false|false|false|C0936188;C1327729;C2362924|Cell septum;Septum - general anatomical term;Septum of telencephalon|septum
Anatomy|Cell Component|SIMPLE_SEGMENT|8599,8605|false|false|false|C0936188;C1327729;C2362924|Cell septum;Septum - general anatomical term;Septum of telencephalon|septum
Finding|Functional Concept|SIMPLE_SEGMENT|8612,8616|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|8612,8635|false|false|false|C0503990|Cavity of left ventricle|left ventricular cavity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8612,8640|false|false|false|C0455830|Left ventricular cavity size|left ventricular cavity size
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8617,8628|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|8617,8635|false|false|false|C0507083|Cavity of ventricle|ventricular cavity
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|8629,8635|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|8629,8635|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8629,8635|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Event|Event|SIMPLE_SEGMENT|8636,8640|false|false|false|||size
Event|Event|SIMPLE_SEGMENT|8644,8650|false|false|false|||normal
Finding|Functional Concept|SIMPLE_SEGMENT|8652,8656|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8657,8668|false|false|false|C0018827|Heart Ventricle|ventricular
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|8670,8678|false|false|false|C0039155|Systole|systolic
Event|Event|SIMPLE_SEGMENT|8679,8687|false|false|false|||function
Finding|Finding|SIMPLE_SEGMENT|8679,8687|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|8679,8687|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|8679,8687|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|SIMPLE_SEGMENT|8679,8687|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Event|Event|SIMPLE_SEGMENT|8691,8703|false|false|false|||hyperdynamic
Event|Event|SIMPLE_SEGMENT|8705,8707|false|false|false|||EF
Finding|Functional Concept|SIMPLE_SEGMENT|8716,8721|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8722,8733|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8735,8742|false|false|false|C0935616|chamber [body part]|chamber
Event|Event|SIMPLE_SEGMENT|8752,8756|false|false|false|||free
Finding|Functional Concept|SIMPLE_SEGMENT|8752,8756|false|false|false|C0332296|Free of (attribute)|free
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8757,8768|false|false|false|C1980023|Wall motion|wall motion
Event|Event|SIMPLE_SEGMENT|8762,8768|false|false|false|||motion
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|8762,8768|false|false|false|C0026597|Motion|motion
Event|Event|SIMPLE_SEGMENT|8773,8779|false|false|false|||normal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8785,8791|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8785,8797|false|false|false|C0003501;C4533215|Aortic valve structure;Chest>Aortic valve|aortic valve
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8792,8797|false|false|false|C1186983|Anatomical valve|valve
Event|Event|SIMPLE_SEGMENT|8799,8807|false|false|false|||leaflets
Event|Event|SIMPLE_SEGMENT|8823,8832|false|false|false|||thickened
Finding|Intellectual Product|SIMPLE_SEGMENT|8843,8847|false|false|false|C1547225|Mild Severity of Illness Code|mild
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8848,8854|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8848,8860|false|false|false|C0003501;C4533215|Aortic valve structure;Chest>Aortic valve|aortic valve
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8855,8860|false|false|false|C1186983|Anatomical valve|valve
Event|Event|SIMPLE_SEGMENT|8862,8870|false|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|8862,8870|false|false|false|C1261287|Stenosis|stenosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8872,8877|false|false|false|C1186983|Anatomical valve|valve
Finding|Finding|SIMPLE_SEGMENT|8872,8882|false|false|false|C4687749|Valve Area|valve area
Event|Governmental or Regulatory Activity|SIMPLE_SEGMENT|8878,8882|false|false|false|C1510751|Academic Research Enhancement Awards|area
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|8890,8893|false|false|false|C0555206|Chiari malformation type II|cm2
Event|Event|SIMPLE_SEGMENT|8890,8893|false|false|false|||cm2
Finding|Functional Concept|SIMPLE_SEGMENT|8896,8901|false|false|false|C1883002|Sequence Chromatogram|Trace
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8902,8908|false|false|false|C0003483|Aorta|aortic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8902,8922|false|false|false|C0003504|Aortic Valve Insufficiency|aortic regurgitation
Event|Event|SIMPLE_SEGMENT|8909,8922|false|false|false|||regurgitation
Finding|Finding|SIMPLE_SEGMENT|8909,8922|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|SIMPLE_SEGMENT|8909,8922|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|8909,8922|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Event|Event|SIMPLE_SEGMENT|8927,8931|false|false|false|||seen
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8937,8949|false|false|false|C0026264|Mitral Valve|mitral valve
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8944,8949|false|false|false|C1186983|Anatomical valve|valve
Event|Event|SIMPLE_SEGMENT|8950,8958|false|false|false|||leaflets
Event|Event|SIMPLE_SEGMENT|8970,8979|false|false|false|||thickened
Finding|Finding|SIMPLE_SEGMENT|8991,8997|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|8991,8997|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8998,9026|false|false|false|C0428811|Mitral valve annular calcification|mitral annular calcification
Finding|Finding|SIMPLE_SEGMENT|8998,9026|false|false|false|C1835130|Premature calcification of mitral annulus|mitral annular calcification
Event|Event|SIMPLE_SEGMENT|9013,9026|false|false|false|||calcification
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|9013,9026|false|false|false|C0006660;C0006663;C1533591|Calcification;Calcinosis;Physiologic calcification|calcification
Finding|Pathologic Function|SIMPLE_SEGMENT|9013,9026|false|false|false|C0006660;C0006663;C1533591|Calcification;Calcinosis;Physiologic calcification|calcification
Finding|Finding|SIMPLE_SEGMENT|9028,9036|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|9028,9036|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Event|Event|SIMPLE_SEGMENT|9050,9063|false|false|false|||regurgitation
Finding|Finding|SIMPLE_SEGMENT|9050,9063|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|SIMPLE_SEGMENT|9050,9063|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|9050,9063|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Event|Event|SIMPLE_SEGMENT|9067,9071|false|false|false|||seen
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|9081,9089|false|false|false|C0001166|Acoustics|acoustic
Finding|Finding|SIMPLE_SEGMENT|9081,9099|false|false|false|C1719833|Acoustic shadowing|acoustic shadowing
Event|Event|SIMPLE_SEGMENT|9090,9099|false|false|false|||shadowing
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9090,9099|false|false|false|C0085195;C0600111|Shadowing (Histology);Shadowing (regime/therapy)|shadowing
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9090,9099|false|false|false|C0085195;C0600111|Shadowing (Histology);Shadowing (regime/therapy)|shadowing
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9118,9138|false|false|false|C0026266|Mitral Valve Insufficiency|mitral regurgitation
Event|Event|SIMPLE_SEGMENT|9125,9138|false|false|false|||regurgitation
Finding|Finding|SIMPLE_SEGMENT|9125,9138|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|SIMPLE_SEGMENT|9125,9138|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|9125,9138|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Event|Event|SIMPLE_SEGMENT|9160,9174|false|false|false|||UNDERestimated
Finding|Intellectual Product|SIMPLE_SEGMENT|9187,9191|false|false|false|C1547225|Mild Severity of Illness Code|mild
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9192,9201|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9192,9201|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|9192,9201|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9192,9208|false|false|false|C0034052|Pulmonary artery structure|pulmonary artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9202,9208|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|9202,9208|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|9209,9217|false|false|false|C0039155|Systole|systolic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9209,9230|false|false|false|C0221155|Systolic Hypertension|systolic hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9218,9230|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|SIMPLE_SEGMENT|9218,9230|false|false|false|||hypertension
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9245,9256|true|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9245,9256|true|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9245,9265|true|false|false|C0031039|Pericardial effusion|pericardial effusion
Finding|Body Substance|SIMPLE_SEGMENT|9245,9265|true|false|false|C1253937|Pericardial effusion body substance|pericardial effusion
Event|Event|SIMPLE_SEGMENT|9257,9265|true|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|9257,9265|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|9257,9265|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|9257,9265|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Event|Event|SIMPLE_SEGMENT|9293,9298|false|false|false|||study
Finding|Intellectual Product|SIMPLE_SEGMENT|9293,9298|false|false|false|C1705923|Study Object|study
Procedure|Research Activity|SIMPLE_SEGMENT|9293,9298|false|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|study
Event|Event|SIMPLE_SEGMENT|9317,9325|false|false|false|||reviewed
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9329,9337|false|false|false|C2926606||findings
Event|Event|SIMPLE_SEGMENT|9329,9337|false|false|false|||findings
Finding|Functional Concept|SIMPLE_SEGMENT|9329,9337|false|false|false|C2607943|findings aspects|findings
Event|Event|SIMPLE_SEGMENT|9342,9349|false|false|false|||similar
Finding|Intellectual Product|SIMPLE_SEGMENT|9357,9364|false|false|false|C1550127|Special Handling Code - Upright|UPRIGHT
Phenomenon|Human-caused Phenomenon or Process|SIMPLE_SEGMENT|9357,9364|false|false|false|C1550585|Entity Handling - upright|UPRIGHT
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9365,9370|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|CHEST
Finding|Finding|SIMPLE_SEGMENT|9365,9370|false|false|false|C0741025|Chest problem|CHEST
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9365,9376|false|false|false|C0039985|Plain chest X-ray|CHEST X-RAY
Event|Event|SIMPLE_SEGMENT|9371,9376|false|false|false|||X-RAY
Finding|Functional Concept|SIMPLE_SEGMENT|9371,9376|false|false|false|C0034571;C3244296|ActClaimAttachmentCategoryCode - x-ray;roentgenographic|X-RAY
Finding|Intellectual Product|SIMPLE_SEGMENT|9371,9376|false|false|false|C0034571;C3244296|ActClaimAttachmentCategoryCode - x-ray;roentgenographic|X-RAY
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|9371,9376|false|false|false|C0043309|Roentgen Rays|X-RAY
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9371,9376|false|false|false|C0043299;C1306645;C1962945|Diagnostic radiologic examination;Plain x-ray;Radiographic imaging procedure|X-RAY
Event|Event|SIMPLE_SEGMENT|9384,9392|false|false|false|||Compared
Event|Event|SIMPLE_SEGMENT|9413,9418|false|false|false|||study
Finding|Intellectual Product|SIMPLE_SEGMENT|9413,9418|false|false|false|C1705923|Study Object|study
Procedure|Research Activity|SIMPLE_SEGMENT|9413,9418|false|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|study
Event|Event|SIMPLE_SEGMENT|9429,9440|false|false|false|||improvement
Finding|Conceptual Entity|SIMPLE_SEGMENT|9429,9440|false|false|false|C2986411|Improvement|improvement
Finding|Intellectual Product|SIMPLE_SEGMENT|9449,9453|false|false|false|C1547225|Mild Severity of Illness Code|mild
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9454,9463|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9454,9463|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|9454,9463|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|9454,9469|false|false|false|C0034063|Pulmonary Edema|pulmonary edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9464,9469|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|9464,9469|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|9464,9469|false|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|9475,9483|false|false|false|||decrease
Finding|Finding|SIMPLE_SEGMENT|9475,9483|false|false|false|C0392756|Reduced|decrease
Finding|Functional Concept|SIMPLE_SEGMENT|9498,9502|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Tissue|SIMPLE_SEGMENT|9503,9510|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9503,9510|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Body Substance|SIMPLE_SEGMENT|9503,9519|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Finding|SIMPLE_SEGMENT|9503,9519|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|9503,9519|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Event|Event|SIMPLE_SEGMENT|9511,9519|false|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|9511,9519|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|9511,9519|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|9511,9519|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Finding|SIMPLE_SEGMENT|9521,9529|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|9521,9529|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Functional Concept|SIMPLE_SEGMENT|9530,9535|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Tissue|SIMPLE_SEGMENT|9537,9544|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9537,9544|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Body Substance|SIMPLE_SEGMENT|9537,9553|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Finding|SIMPLE_SEGMENT|9537,9553|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|9537,9553|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Event|Event|SIMPLE_SEGMENT|9545,9553|false|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|9545,9553|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|9545,9553|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|9545,9553|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Event|Event|SIMPLE_SEGMENT|9568,9579|false|false|false|||atelectasis
Finding|Pathologic Function|SIMPLE_SEGMENT|9568,9579|false|false|false|C0004144|Atelectasis|atelectasis
Event|Event|SIMPLE_SEGMENT|9584,9590|false|false|false|||stable
Finding|Intellectual Product|SIMPLE_SEGMENT|9584,9590|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Intellectual Product|SIMPLE_SEGMENT|9597,9604|false|false|false|C1550127|Special Handling Code - Upright|UPRIGHT
Phenomenon|Human-caused Phenomenon or Process|SIMPLE_SEGMENT|9597,9604|false|false|false|C1550585|Entity Handling - upright|UPRIGHT
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9605,9610|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|CHEST
Finding|Finding|SIMPLE_SEGMENT|9605,9610|false|false|false|C0741025|Chest problem|CHEST
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9605,9616|false|false|false|C0039985|Plain chest X-ray|CHEST X-RAY
Event|Event|SIMPLE_SEGMENT|9611,9616|false|false|false|||X-RAY
Finding|Functional Concept|SIMPLE_SEGMENT|9611,9616|false|false|false|C0034571;C3244296|ActClaimAttachmentCategoryCode - x-ray;roentgenographic|X-RAY
Finding|Intellectual Product|SIMPLE_SEGMENT|9611,9616|false|false|false|C0034571;C3244296|ActClaimAttachmentCategoryCode - x-ray;roentgenographic|X-RAY
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|9611,9616|false|false|false|C0043309|Roentgen Rays|X-RAY
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9611,9616|false|false|false|C0043299;C1306645;C1962945|Diagnostic radiologic examination;Plain x-ray;Radiographic imaging procedure|X-RAY
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9624,9631|false|false|false|C0018787|Heart|Cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|9624,9631|false|false|false|C1314974|Cardiac attachment|Cardiac
Event|Event|SIMPLE_SEGMENT|9632,9636|false|false|false|||size
Event|Event|SIMPLE_SEGMENT|9640,9646|false|false|false|||normal
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9648,9653|false|false|false|C1517938|Long Interspersed Elements|Lines
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|9648,9653|false|false|false|C1517938|Long Interspersed Elements|Lines
Event|Event|SIMPLE_SEGMENT|9648,9653|false|false|false|||Lines
Finding|Idea or Concept|SIMPLE_SEGMENT|9648,9653|false|false|false|C1548328|Lines Quantity Limit Request|Lines
Event|Event|SIMPLE_SEGMENT|9659,9664|false|false|false|||tubes
Finding|Intellectual Product|SIMPLE_SEGMENT|9659,9664|false|false|false|C1547937||tubes
Finding|Idea or Concept|SIMPLE_SEGMENT|9677,9685|false|false|false|C1548173;C2828392|Standard (document);Type of Agreement - Standard|standard
Finding|Intellectual Product|SIMPLE_SEGMENT|9677,9685|false|false|false|C1548173;C2828392|Standard (document);Type of Agreement - Standard|standard
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9677,9685|false|false|false|C3873211|Standard base excess calculation technique|standard
Event|Event|SIMPLE_SEGMENT|9686,9694|false|false|false|||position
Finding|Gene or Genome|SIMPLE_SEGMENT|9696,9701|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|Large
Event|Event|SIMPLE_SEGMENT|9702,9707|false|false|false|||right
Finding|Functional Concept|SIMPLE_SEGMENT|9702,9707|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Event|Event|SIMPLE_SEGMENT|9712,9720|false|false|false|||moderate
Finding|Finding|SIMPLE_SEGMENT|9712,9720|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|9712,9720|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Functional Concept|SIMPLE_SEGMENT|9722,9726|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Tissue|SIMPLE_SEGMENT|9727,9734|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9727,9734|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Pathologic Function|SIMPLE_SEGMENT|9727,9744|false|false|false|C0032227|Pleural effusion (disorder)|pleural effusions
Event|Event|SIMPLE_SEGMENT|9735,9744|false|false|false|||effusions
Finding|Pathologic Function|SIMPLE_SEGMENT|9735,9744|false|false|false|C0013687|effusion|effusions
Event|Event|SIMPLE_SEGMENT|9757,9766|false|false|false|||unchanged
Finding|Finding|SIMPLE_SEGMENT|9757,9766|false|false|false|C0442739||unchanged
Event|Event|SIMPLE_SEGMENT|9797,9808|false|false|false|||positioning
Procedure|Health Care Activity|SIMPLE_SEGMENT|9797,9808|false|false|false|C0150305;C1561964|Positioning - therapy;Positioning patient (procedure)|positioning
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9797,9808|false|false|false|C0150305;C1561964|Positioning - therapy;Positioning patient (procedure)|positioning
Finding|Body Substance|SIMPLE_SEGMENT|9816,9823|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|9816,9823|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|9816,9823|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|SIMPLE_SEGMENT|9825,9830|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9825,9841|false|false|false|C1261074|Structure of right upper lobe of lung|Right upper lobe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9831,9841|false|false|false|C0225756|Structure of upper lobe of lung|upper lobe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9837,9841|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|SIMPLE_SEGMENT|9837,9841|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Event|Event|SIMPLE_SEGMENT|9843,9850|false|false|false|||opacity
Finding|Finding|SIMPLE_SEGMENT|9843,9850|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacity
Finding|Pathologic Function|SIMPLE_SEGMENT|9843,9850|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacity
Event|Event|SIMPLE_SEGMENT|9855,9863|false|false|false|||improved
Event|Event|SIMPLE_SEGMENT|9864,9874|false|false|false|||consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|9864,9874|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|9864,9879|false|false|false|C0332290|Consistent with|consistent with
Event|Event|SIMPLE_SEGMENT|9880,9889|false|false|false|||improving
Event|Event|SIMPLE_SEGMENT|9890,9901|false|false|false|||atelectasis
Finding|Pathologic Function|SIMPLE_SEGMENT|9890,9901|false|false|false|C0004144|Atelectasis|atelectasis
Anatomy|Tissue|SIMPLE_SEGMENT|9904,9911|false|false|false|C0032225|Pleura|Pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9904,9911|false|false|false|C0032226|Pleural Diseases|Pleural
Finding|Pathologic Function|SIMPLE_SEGMENT|9904,9921|false|false|false|C0032227|Pleural effusion (disorder)|Pleural effusions
Event|Event|SIMPLE_SEGMENT|9912,9921|false|false|false|||effusions
Finding|Pathologic Function|SIMPLE_SEGMENT|9912,9921|false|false|false|C0013687|effusion|effusions
Event|Event|SIMPLE_SEGMENT|9926,9936|false|false|false|||associated
Event|Event|SIMPLE_SEGMENT|9942,9953|false|false|false|||atelectasis
Finding|Pathologic Function|SIMPLE_SEGMENT|9942,9953|false|false|false|C0004144|Atelectasis|atelectasis
Finding|Functional Concept|SIMPLE_SEGMENT|9970,9975|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Finding|Intellectual Product|SIMPLE_SEGMENT|9991,9995|false|false|false|C1547225|Mild Severity of Illness Code|mild
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9996,10004|false|false|false|C0005847|Blood Vessel|vascular
Event|Event|SIMPLE_SEGMENT|10005,10015|false|false|false|||congestion
Finding|Pathologic Function|SIMPLE_SEGMENT|10005,10015|false|false|false|C0700148|Congestion|congestion
Finding|Intellectual Product|SIMPLE_SEGMENT|10020,10025|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|10026,10034|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10026,10041|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|10026,10041|false|false|false|C0489547|Hospital course|Hospital Course
Finding|Idea or Concept|SIMPLE_SEGMENT|10043,10051|false|false|false|C1547192|Organization unit type - Hospital|HOSPITAL
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10043,10058|false|false|false|C0488549||HOSPITAL COURSE
Finding|Finding|SIMPLE_SEGMENT|10043,10058|false|false|false|C0489547|Hospital course|HOSPITAL COURSE
Event|Event|SIMPLE_SEGMENT|10052,10058|false|false|false|||COURSE
Finding|Idea or Concept|SIMPLE_SEGMENT|10075,10079|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|SIMPLE_SEGMENT|10075,10079|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|SIMPLE_SEGMENT|10084,10089|false|false|false|||woman
Event|Event|SIMPLE_SEGMENT|10100,10112|false|false|false|||hospitalized
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10131,10137|false|false|false|C0036690;C0243026|Sepsis;Septicemia|sepsis
Event|Event|SIMPLE_SEGMENT|10131,10137|false|false|false|||sepsis
Event|Event|SIMPLE_SEGMENT|10142,10147|false|false|false|||shock
Finding|Pathologic Function|SIMPLE_SEGMENT|10142,10147|false|false|false|C0036974|Shock|shock
Event|Event|SIMPLE_SEGMENT|10149,10160|false|false|false|||complicated
Event|Event|SIMPLE_SEGMENT|10164,10175|false|false|false|||readmission
Procedure|Health Care Activity|SIMPLE_SEGMENT|10164,10175|false|false|false|C4489276|Readmission|readmission
Event|Event|SIMPLE_SEGMENT|10177,10184|false|false|false|||hypoxia
Finding|Finding|SIMPLE_SEGMENT|10177,10184|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|hypoxia
Finding|Pathologic Function|SIMPLE_SEGMENT|10177,10184|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|hypoxia
Event|Event|SIMPLE_SEGMENT|10185,10196|false|false|false|||hypercarbia
Finding|Finding|SIMPLE_SEGMENT|10185,10196|false|false|false|C0020440|Hypercapnia|hypercarbia
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10219,10230|false|false|false|C0231832|Respiratory rate|respiratory
Event|Event|SIMPLE_SEGMENT|10219,10230|false|false|false|||respiratory
Finding|Body Substance|SIMPLE_SEGMENT|10219,10230|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|SIMPLE_SEGMENT|10219,10230|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|SIMPLE_SEGMENT|10219,10230|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Event|Event|SIMPLE_SEGMENT|10232,10239|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|10232,10239|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|10232,10239|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|10232,10239|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10244,10251|false|false|false|C0042027|Urinary tract|urinary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10244,10257|false|false|false|C0042027;C1508753|Urinary system;Urinary tract|urinary tract
Anatomy|Body System|SIMPLE_SEGMENT|10244,10257|false|false|false|C0042027;C1508753|Urinary system;Urinary tract|urinary tract
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10244,10267|false|false|false|C0042029|Urinary tract infection|urinary tract infection
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10252,10257|false|false|false|C1185740|Tract|tract
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10258,10267|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|10258,10267|false|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|10258,10267|false|false|false|C3714514|Infection|infection
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10286,10297|false|false|false|C0231832|Respiratory rate|Respiratory
Finding|Body Substance|SIMPLE_SEGMENT|10286,10297|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|Respiratory
Finding|Functional Concept|SIMPLE_SEGMENT|10286,10297|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|Respiratory
Finding|Intellectual Product|SIMPLE_SEGMENT|10286,10297|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|Respiratory
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10286,10305|false|false|false|C1145670|Respiratory Failure|Respiratory Failure
Event|Event|SIMPLE_SEGMENT|10298,10305|false|false|false|||Failure
Finding|Functional Concept|SIMPLE_SEGMENT|10298,10305|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|Failure
Finding|Idea or Concept|SIMPLE_SEGMENT|10298,10305|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|Failure
Finding|Individual Behavior|SIMPLE_SEGMENT|10298,10305|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|Failure
Finding|Conceptual Entity|SIMPLE_SEGMENT|10307,10315|false|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|Etiology
Finding|Functional Concept|SIMPLE_SEGMENT|10307,10315|false|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|Etiology
Finding|Finding|SIMPLE_SEGMENT|10316,10322|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|10316,10322|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|SIMPLE_SEGMENT|10324,10338|false|false|false|||multifactorial
Finding|Finding|SIMPLE_SEGMENT|10324,10338|false|false|false|C1837655|Multifactorial|multifactorial
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10350,10361|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|SIMPLE_SEGMENT|10350,10361|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|SIMPLE_SEGMENT|10350,10361|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|SIMPLE_SEGMENT|10350,10361|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10350,10368|false|false|false|C0035231|Respiratory Muscles|respiratory muscle
Finding|Finding|SIMPLE_SEGMENT|10350,10377|false|false|false|C1836141;C3806467|Respiratory insufficiency due to muscle weakness;Respiratory muscle weakness|respiratory muscle weakness
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10362,10368|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|SIMPLE_SEGMENT|10362,10368|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10362,10377|false|false|false|C0030552|Paresis|muscle weakness
Finding|Sign or Symptom|SIMPLE_SEGMENT|10362,10377|false|false|false|C0151786|Muscle Weakness|muscle weakness
Event|Event|SIMPLE_SEGMENT|10369,10377|false|false|false|||weakness
Finding|Sign or Symptom|SIMPLE_SEGMENT|10369,10377|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Event|Event|SIMPLE_SEGMENT|10382,10386|false|false|false|||pulm
Procedure|Health Care Activity|SIMPLE_SEGMENT|10382,10386|false|false|false|C1315068|Pulmonary ventilator management|pulm
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10388,10393|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|10388,10393|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|10388,10393|false|false|false|C0013604|Edema|edema
Anatomy|Tissue|SIMPLE_SEGMENT|10399,10406|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10399,10406|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Pathologic Function|SIMPLE_SEGMENT|10399,10416|false|false|false|C0032227|Pleural effusion (disorder)|pleural effusions
Event|Event|SIMPLE_SEGMENT|10407,10416|false|false|false|||effusions
Finding|Pathologic Function|SIMPLE_SEGMENT|10407,10416|false|false|false|C0013687|effusion|effusions
Event|Event|SIMPLE_SEGMENT|10420,10425|false|false|false|||noted
Procedure|Health Care Activity|SIMPLE_SEGMENT|10429,10438|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|10439,10444|false|false|false|||x-ray
Finding|Functional Concept|SIMPLE_SEGMENT|10439,10444|false|false|false|C0034571;C3244296|ActClaimAttachmentCategoryCode - x-ray;roentgenographic|x-ray
Finding|Intellectual Product|SIMPLE_SEGMENT|10439,10444|false|false|false|C0034571;C3244296|ActClaimAttachmentCategoryCode - x-ray;roentgenographic|x-ray
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|10439,10444|false|false|false|C0043309|Roentgen Rays|x-ray
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10439,10444|false|false|false|C0043299;C1306645;C1962945|Diagnostic radiologic examination;Plain x-ray;Radiographic imaging procedure|x-ray
Event|Event|SIMPLE_SEGMENT|10451,10458|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|10451,10458|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|10451,10458|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|10451,10458|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|10451,10461|false|false|false|C0262926|Medical History|history of
Event|Event|SIMPLE_SEGMENT|10485,10493|false|false|false|||remained
Event|Event|SIMPLE_SEGMENT|10494,10503|false|false|false|||intubated
Finding|Finding|SIMPLE_SEGMENT|10494,10503|false|false|false|C4698386|Intubated|intubated
Event|Event|SIMPLE_SEGMENT|10526,10530|false|false|false|||stay
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10538,10547|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10538,10547|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|10538,10547|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|10538,10553|false|false|false|C0034063|Pulmonary Edema|pulmonary edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10548,10553|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|10548,10553|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|10548,10553|false|false|false|C0013604|Edema|edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10558,10569|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|SIMPLE_SEGMENT|10558,10569|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|SIMPLE_SEGMENT|10558,10569|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|SIMPLE_SEGMENT|10558,10569|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10558,10576|false|false|false|C0035231|Respiratory Muscles|respiratory muscle
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10570,10576|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|SIMPLE_SEGMENT|10570,10576|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Event|Event|SIMPLE_SEGMENT|10578,10586|false|false|false|||weakness
Finding|Sign or Symptom|SIMPLE_SEGMENT|10578,10586|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Finding|Intellectual Product|SIMPLE_SEGMENT|10594,10598|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Finding|Classification|SIMPLE_SEGMENT|10599,10607|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|10599,10607|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|10599,10607|false|false|false|C5237010|Expression Negative|negative
Event|Event|SIMPLE_SEGMENT|10608,10619|false|false|false|||inspiratory
Finding|Organism Function|SIMPLE_SEGMENT|10608,10619|false|false|false|C0004048|Inspiration (function)|inspiratory
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|10608,10625|false|false|false|C0231823|Inspiratory force|inspiratory force
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|10620,10625|false|false|false|C0441722;C0563538|Force;Mechanical force|force
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10627,10630|false|false|false|C4281719;C4281724|Protein S100-A8;Protein S100-A9|NIF
Drug|Immunologic Factor|SIMPLE_SEGMENT|10627,10630|false|false|false|C4281719;C4281724|Protein S100-A8;Protein S100-A9|NIF
Event|Event|SIMPLE_SEGMENT|10627,10630|false|false|false|||NIF
Finding|Gene or Genome|SIMPLE_SEGMENT|10627,10630|false|false|false|C1335798;C1704874;C1704875|S100A8 wt Allele;S100A9 gene;S100A9 wt Allele|NIF
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10637,10640|false|false|false|C4281719;C4281724|Protein S100-A8;Protein S100-A9|NIF
Drug|Immunologic Factor|SIMPLE_SEGMENT|10637,10640|false|false|false|C4281719;C4281724|Protein S100-A8;Protein S100-A9|NIF
Event|Event|SIMPLE_SEGMENT|10637,10640|false|false|false|||NIF
Finding|Gene or Genome|SIMPLE_SEGMENT|10637,10640|false|false|false|C1335798;C1704874;C1704875|S100A8 wt Allele;S100A9 gene;S100A9 wt Allele|NIF
Event|Event|SIMPLE_SEGMENT|10652,10660|false|false|false|||improved
Event|Activity|SIMPLE_SEGMENT|10666,10678|false|false|false|C2698650|Optimization|optimization
Event|Event|SIMPLE_SEGMENT|10666,10678|false|false|false|||optimization
Event|Event|SIMPLE_SEGMENT|10686,10695|false|false|false|||nutrition
Finding|Finding|SIMPLE_SEGMENT|10686,10695|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|nutrition
Finding|Intellectual Product|SIMPLE_SEGMENT|10686,10695|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|nutrition
Finding|Organism Function|SIMPLE_SEGMENT|10686,10695|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|nutrition
Procedure|Research Activity|SIMPLE_SEGMENT|10686,10695|false|false|false|C0600072;C1521729|Feeding and dietary regimes;Nutritional Study|nutrition
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10686,10695|false|false|false|C0600072;C1521729|Feeding and dietary regimes;Nutritional Study|nutrition
Finding|Conceptual Entity|SIMPLE_SEGMENT|10701,10711|false|false|false|C1521721|Supportive assistance|supportive
Procedure|Health Care Activity|SIMPLE_SEGMENT|10701,10716|false|false|false|C0030231;C0344211|Palliative Care;Supportive care|supportive care
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10701,10716|false|false|false|C0030231;C0344211|Palliative Care;Supportive care|supportive care
Event|Activity|SIMPLE_SEGMENT|10712,10716|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|10712,10716|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|10712,10716|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|10712,10716|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10722,10731|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10722,10731|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|10722,10731|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|10722,10737|false|false|false|C0034063|Pulmonary Edema|pulmonary edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10732,10737|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|10732,10737|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|10732,10737|false|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|10742,10751|false|false|false|||addressed
Finding|Individual Behavior|SIMPLE_SEGMENT|10758,10768|false|false|false|C0001807;C1547300;C1548760|Aggressive behavior;Precaution Code - Aggressive;Risk Codes - Aggressive|aggressive
Finding|Intellectual Product|SIMPLE_SEGMENT|10758,10768|false|false|false|C0001807;C1547300;C1548760|Aggressive behavior;Precaution Code - Aggressive;Risk Codes - Aggressive|aggressive
Event|Event|SIMPLE_SEGMENT|10769,10777|false|false|false|||diuresis
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|10769,10777|false|false|false|C0012797|Diuresis|diuresis
Drug|Organic Chemical|SIMPLE_SEGMENT|10793,10798|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10793,10798|false|false|false|C0699992|Lasix|Lasix
Event|Event|SIMPLE_SEGMENT|10799,10806|false|false|false|||boluses
Finding|Finding|SIMPLE_SEGMENT|10817,10821|false|false|false|C5575035|Well (answer to question)|well
Drug|Organic Chemical|SIMPLE_SEGMENT|10826,10831|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10826,10831|false|false|false|C0699992|Lasix|Lasix
Event|Event|SIMPLE_SEGMENT|10847,10856|false|false|false|||treatment
Finding|Conceptual Entity|SIMPLE_SEGMENT|10847,10856|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|SIMPLE_SEGMENT|10847,10856|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|SIMPLE_SEGMENT|10847,10856|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10847,10856|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Event|Event|SIMPLE_SEGMENT|10866,10872|false|false|false|||issues
Event|Event|SIMPLE_SEGMENT|10882,10886|false|false|false|||able
Finding|Finding|SIMPLE_SEGMENT|10882,10886|false|false|false|C1299581|Able (qualifier value)|able
Event|Event|SIMPLE_SEGMENT|10907,10916|false|false|false|||extubated
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10920,10925|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10920,10925|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|SIMPLE_SEGMENT|10920,10925|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10920,10925|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|SIMPLE_SEGMENT|10920,10925|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|SIMPLE_SEGMENT|10920,10925|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10926,10933|false|false|false|C1550232|Body Parts - Cannula|cannula
Finding|Body Substance|SIMPLE_SEGMENT|10926,10933|false|false|false|C1546577;C1550622|Specimen Type - Cannula|cannula
Finding|Intellectual Product|SIMPLE_SEGMENT|10926,10933|false|false|false|C1546577;C1550622|Specimen Type - Cannula|cannula
Event|Event|SIMPLE_SEGMENT|10951,10958|false|false|false|||started
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10962,10972|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10962,10972|false|false|false|C0065374|lisinopril|Lisinopril
Event|Event|SIMPLE_SEGMENT|10973,10976|false|false|false|||5mg
Event|Event|SIMPLE_SEGMENT|10997,11006|false|false|false|||reduction
Finding|Finding|SIMPLE_SEGMENT|10997,11006|false|false|false|C0392756|Reduced|reduction
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|10997,11006|false|false|false|C0301630|Reduction (chemical)|reduction
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10997,11006|false|false|false|C1293152;C4551656|Reduction procedure;Surgical reduction|reduction
Event|Event|SIMPLE_SEGMENT|11012,11019|false|false|false|||setting
Finding|Mental Process|SIMPLE_SEGMENT|11012,11019|false|false|false|C0542559|contextual factors|setting
Event|Event|SIMPLE_SEGMENT|11053,11060|false|false|false|||causing
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11065,11074|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11065,11074|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|11065,11074|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11076,11081|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|11076,11081|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|11076,11081|false|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|11091,11098|false|false|false|||require
Event|Event|SIMPLE_SEGMENT|11107,11110|false|false|false|||PRN
Finding|Gene or Genome|SIMPLE_SEGMENT|11107,11110|false|true|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|11111,11116|false|false|false|||doses
Drug|Organic Chemical|SIMPLE_SEGMENT|11120,11125|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11120,11125|false|false|false|C0699992|Lasix|Lasix
Event|Event|SIMPLE_SEGMENT|11120,11125|false|false|false|||Lasix
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11129,11134|false|false|false|C0034991|Rehabilitation therapy|rehab
Drug|Organic Chemical|SIMPLE_SEGMENT|11153,11158|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11153,11158|false|false|false|C0699992|Lasix|Lasix
Event|Event|SIMPLE_SEGMENT|11167,11170|false|false|false|||PRN
Finding|Gene or Genome|SIMPLE_SEGMENT|11167,11170|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|11172,11180|false|false|false|||Consider
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11192,11202|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11192,11202|false|false|false|C0065374|lisinopril|lisinopril
Event|Event|SIMPLE_SEGMENT|11192,11202|false|false|false|||lisinopril
Finding|Idea or Concept|SIMPLE_SEGMENT|11216,11222|false|false|false|C1550462|Observation Interpretation - better|better
Event|Event|SIMPLE_SEGMENT|11233,11242|false|false|false|||reduction
Finding|Finding|SIMPLE_SEGMENT|11233,11242|false|false|false|C0392756|Reduced|reduction
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|11233,11242|false|false|false|C0301630|Reduction (chemical)|reduction
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11233,11242|false|false|false|C1293152;C4551656|Reduction procedure;Surgical reduction|reduction
Finding|Finding|SIMPLE_SEGMENT|11243,11251|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|11243,11251|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|11243,11251|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|11243,11251|false|false|false|C0033095||pressure
Event|Event|SIMPLE_SEGMENT|11252,11262|false|false|false|||tolerating
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11268,11279|false|false|false|C0033817|Pseudomonas Infections|Pseudomonas
Event|Event|SIMPLE_SEGMENT|11268,11279|false|false|false|||Pseudomonas
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11280,11283|false|false|false|C0042029|Urinary tract infection|UTI
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11280,11283|false|false|false|C0077906|urinastatin|UTI
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11280,11283|false|false|false|C0077906|urinastatin|UTI
Event|Event|SIMPLE_SEGMENT|11280,11283|false|false|false|||UTI
Finding|Gene or Genome|SIMPLE_SEGMENT|11280,11283|false|false|false|C1412376;C5780748|AMBP gene;AMBP wt Allele|UTI
Finding|Body Substance|SIMPLE_SEGMENT|11285,11292|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|11285,11292|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|11285,11292|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|11293,11297|false|false|false|||grew
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11302,11313|false|false|false|C0033817|Pseudomonas Infections|Pseudomonas
Event|Event|SIMPLE_SEGMENT|11302,11313|false|false|false|||Pseudomonas
Event|Event|SIMPLE_SEGMENT|11314,11323|false|false|false|||sensitive
Finding|Functional Concept|SIMPLE_SEGMENT|11314,11323|false|false|false|C0332324|Sensitive|sensitive
Finding|Functional Concept|SIMPLE_SEGMENT|11314,11326|false|false|false|C0332324|Sensitive|sensitive to
Drug|Antibiotic|SIMPLE_SEGMENT|11343,11353|false|false|false|C3854019|gentamicin|Gentamicin
Drug|Organic Chemical|SIMPLE_SEGMENT|11343,11353|false|false|false|C3854019|gentamicin|Gentamicin
Event|Event|SIMPLE_SEGMENT|11343,11353|false|false|false|||Gentamicin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11343,11353|false|false|false|C0202391|Gentamicin measurement|Gentamicin
Finding|Body Substance|SIMPLE_SEGMENT|11361,11366|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|SIMPLE_SEGMENT|11361,11366|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|SIMPLE_SEGMENT|11361,11366|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11361,11374|false|false|false|C0430404|Urine culture|urine culture
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11367,11374|false|false|false|C1706355|Culture Dose Form|culture
Event|Event|SIMPLE_SEGMENT|11367,11374|false|false|false|||culture
Finding|Functional Concept|SIMPLE_SEGMENT|11367,11374|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Finding|Idea or Concept|SIMPLE_SEGMENT|11367,11374|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11367,11374|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|culture
Event|Event|SIMPLE_SEGMENT|11395,11402|false|false|false|||started
Event|Activity|SIMPLE_SEGMENT|11406,11412|false|false|false|C1705764|Doubling|double
Finding|Functional Concept|SIMPLE_SEGMENT|11406,11412|false|false|false|C0205173|Double (qualifier value)|double
Event|Event|SIMPLE_SEGMENT|11413,11421|false|false|false|||coverage
Finding|Functional Concept|SIMPLE_SEGMENT|11413,11421|false|false|false|C1551362;C1999244;C3854012|coverage - HL7PublishingDomain;coverage - financial contract|coverage
Finding|Idea or Concept|SIMPLE_SEGMENT|11413,11421|false|false|false|C1551362;C1999244;C3854012|coverage - HL7PublishingDomain;coverage - financial contract|coverage
Finding|Intellectual Product|SIMPLE_SEGMENT|11413,11421|false|false|false|C1551362;C1999244;C3854012|coverage - HL7PublishingDomain;coverage - financial contract|coverage
Drug|Organic Chemical|SIMPLE_SEGMENT|11427,11432|false|false|false|C0701042|Cipro|Cipro
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11427,11432|false|false|false|C0701042|Cipro|Cipro
Drug|Antibiotic|SIMPLE_SEGMENT|11433,11441|false|false|false|C0055003|cefepime|Cefepime
Drug|Organic Chemical|SIMPLE_SEGMENT|11433,11441|false|false|false|C0055003|cefepime|Cefepime
Event|Event|SIMPLE_SEGMENT|11449,11457|false|false|false|||cultures
Finding|Idea or Concept|SIMPLE_SEGMENT|11449,11457|false|false|false|C0010453|Culture (Anthropological)|cultures
Event|Event|SIMPLE_SEGMENT|11458,11465|false|false|false|||pending
Finding|Idea or Concept|SIMPLE_SEGMENT|11458,11465|false|false|false|C1691786;C1704475|Pending - Allergy Clinical Status;Pending - referral status|pending
Finding|Intellectual Product|SIMPLE_SEGMENT|11467,11471|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|SIMPLE_SEGMENT|11472,11480|false|false|false|||narrowed
Drug|Antibiotic|SIMPLE_SEGMENT|11484,11492|false|false|false|C0055003|cefepime|Cefepime
Drug|Organic Chemical|SIMPLE_SEGMENT|11484,11492|false|false|false|C0055003|cefepime|Cefepime
Finding|Finding|SIMPLE_SEGMENT|11493,11498|false|false|false|C0439044|Living Alone|alone
Finding|Intellectual Product|SIMPLE_SEGMENT|11500,11504|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|SIMPLE_SEGMENT|11506,11515|false|false|false|||broadened
Event|Event|SIMPLE_SEGMENT|11536,11540|false|false|false|||recs
Event|Event|SIMPLE_SEGMENT|11552,11559|false|false|false|||concern
Finding|Idea or Concept|SIMPLE_SEGMENT|11552,11559|false|false|false|C2699424|Concern|concern
Event|Event|SIMPLE_SEGMENT|11576,11582|false|false|false|||caused
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11585,11589|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|drug
Finding|Finding|SIMPLE_SEGMENT|11585,11589|false|false|false|C0740721|Drug problem|drug
Finding|Pathologic Function|SIMPLE_SEGMENT|11585,11594|false|false|false|C0011609|Drug Eruptions|drug rash
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11590,11594|false|false|false|C5779629|Eruption of skin (disorder)|rash
Event|Event|SIMPLE_SEGMENT|11590,11594|false|false|false|||rash
Finding|Pathologic Function|SIMPLE_SEGMENT|11590,11594|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|SIMPLE_SEGMENT|11590,11594|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Intellectual Product|SIMPLE_SEGMENT|11606,11610|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|SIMPLE_SEGMENT|11611,11619|false|false|false|||switched
Drug|Antibiotic|SIMPLE_SEGMENT|11627,11632|false|false|false|C0250482|Zosyn|Zosyn
Drug|Organic Chemical|SIMPLE_SEGMENT|11627,11632|false|false|false|C0250482|Zosyn|Zosyn
Event|Event|SIMPLE_SEGMENT|11638,11647|false|false|false|||completed
Drug|Antibiotic|SIMPLE_SEGMENT|11648,11653|false|false|false|C0250482|Zosyn|Zosyn
Drug|Organic Chemical|SIMPLE_SEGMENT|11648,11653|false|false|false|C0250482|Zosyn|Zosyn
Drug|Antibiotic|SIMPLE_SEGMENT|11696,11707|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|SIMPLE_SEGMENT|11696,11707|false|false|false|||antibiotics
Finding|Functional Concept|SIMPLE_SEGMENT|11712,11723|false|false|false|C0231242|Complicated|complicated
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11724,11727|false|false|false|C0042029|Urinary tract infection|UTI
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11724,11727|false|false|false|C0077906|urinastatin|UTI
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11724,11727|false|false|false|C0077906|urinastatin|UTI
Event|Event|SIMPLE_SEGMENT|11724,11727|false|false|false|||UTI
Finding|Gene or Genome|SIMPLE_SEGMENT|11724,11727|false|false|false|C1412376;C5780748|AMBP gene;AMBP wt Allele|UTI
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11734,11738|false|false|false|C5779629|Eruption of skin (disorder)|RASH
Event|Event|SIMPLE_SEGMENT|11734,11738|false|false|false|||RASH
Finding|Pathologic Function|SIMPLE_SEGMENT|11734,11738|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|RASH
Finding|Sign or Symptom|SIMPLE_SEGMENT|11734,11738|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|RASH
Event|Event|SIMPLE_SEGMENT|11743,11748|false|false|false|||noted
Finding|Finding|SIMPLE_SEGMENT|11757,11760|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Finding|Gene or Genome|SIMPLE_SEGMENT|11757,11760|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Finding|Sign or Symptom|SIMPLE_SEGMENT|11761,11773|false|false|false|C0221201|Macular rash|macular rash
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11769,11773|false|false|false|C5779629|Eruption of skin (disorder)|rash
Event|Event|SIMPLE_SEGMENT|11769,11773|false|false|false|||rash
Finding|Pathologic Function|SIMPLE_SEGMENT|11769,11773|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|SIMPLE_SEGMENT|11769,11773|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11777,11788|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Event|Event|SIMPLE_SEGMENT|11805,11814|false|false|false|||meropenam
Event|Event|SIMPLE_SEGMENT|11826,11834|false|false|false|||presumed
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11851,11855|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|drug
Finding|Finding|SIMPLE_SEGMENT|11851,11855|false|false|false|C0740721|Drug problem|drug
Finding|Pathologic Function|SIMPLE_SEGMENT|11851,11860|false|true|false|C0011609|Drug Eruptions|drug rash
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11856,11860|false|true|false|C5779629|Eruption of skin (disorder)|rash
Event|Event|SIMPLE_SEGMENT|11856,11860|false|false|false|||rash
Finding|Pathologic Function|SIMPLE_SEGMENT|11856,11860|false|true|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|SIMPLE_SEGMENT|11856,11860|false|true|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Event|Event|SIMPLE_SEGMENT|11865,11874|false|false|false|||meropenam
Event|Event|SIMPLE_SEGMENT|11879,11886|false|false|false|||stopped
Event|Event|SIMPLE_SEGMENT|11911,11919|false|false|false|||believed
Event|Event|SIMPLE_SEGMENT|11932,11942|false|false|false|||consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|11932,11942|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|11932,11947|false|false|false|C0332290|Consistent with|consistent with
Event|Activity|SIMPLE_SEGMENT|11948,11955|false|true|false|C3812666|Personal Contact|contact
Finding|Functional Concept|SIMPLE_SEGMENT|11948,11955|false|true|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|contact
Finding|Idea or Concept|SIMPLE_SEGMENT|11948,11955|false|true|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|contact
Finding|Intellectual Product|SIMPLE_SEGMENT|11948,11955|false|true|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|contact
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|11948,11955|false|true|false|C0392367|Physical contact|contact
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11948,11966|false|true|false|C0011616|Contact Dermatitis|contact dermatitis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11956,11966|false|true|false|C0011603|Dermatitis|dermatitis
Event|Event|SIMPLE_SEGMENT|11956,11966|false|false|false|||dermatitis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11971,11977|false|false|false|C0013595|Eczema|eczema
Event|Event|SIMPLE_SEGMENT|11971,11977|false|false|false|||eczema
Drug|Organic Chemical|SIMPLE_SEGMENT|11980,11993|false|false|false|C0040864|triamcinolone|Triamcinolone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11980,11993|false|false|false|C0040864|triamcinolone|Triamcinolone
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11994,11999|false|false|false|C0700385;C0705539;C1378128|Cream;Dairy Cream;Emollient Cream|cream
Drug|Food|SIMPLE_SEGMENT|11994,11999|false|false|false|C0700385;C0705539;C1378128|Cream;Dairy Cream;Emollient Cream|cream
Event|Event|SIMPLE_SEGMENT|11994,11999|false|false|false|||cream
Event|Event|SIMPLE_SEGMENT|12004,12011|false|false|false|||started
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12016,12020|false|false|false|C5779629|Eruption of skin (disorder)|rash
Event|Event|SIMPLE_SEGMENT|12016,12020|false|false|false|||rash
Finding|Pathologic Function|SIMPLE_SEGMENT|12016,12020|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|SIMPLE_SEGMENT|12016,12020|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Event|Event|SIMPLE_SEGMENT|12021,12029|false|false|false|||improved
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12043,12050|false|false|false|C0009319|Colitis|Colitis
Event|Event|SIMPLE_SEGMENT|12043,12050|false|false|false|||Colitis
Finding|Body Substance|SIMPLE_SEGMENT|12052,12059|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|12052,12059|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|12052,12059|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|12073,12081|false|false|false|||admitted
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12095,12102|false|true|false|C0009319|Colitis|colitis
Event|Event|SIMPLE_SEGMENT|12095,12102|false|false|false|||colitis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12108,12114|false|false|false|C0036690;C0243026|Sepsis;Septicemia|sepsis
Event|Event|SIMPLE_SEGMENT|12108,12114|false|false|false|||sepsis
Finding|Functional Concept|SIMPLE_SEGMENT|12116,12122|false|false|false|C0205341;C1705914|Repeat;Repeat Object|Repeat
Event|Event|SIMPLE_SEGMENT|12130,12133|false|false|false|||PCR
Finding|Finding|SIMPLE_SEGMENT|12130,12133|false|false|false|C4050242;C5202919|Pathologic Complete Response;Residual Cancer Burden Class 0|PCR
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12130,12133|false|false|false|C0032520;C3853643|Polymerase Chain Reaction;Probe with target amplification technique|PCR
Procedure|Molecular Biology Research Technique|SIMPLE_SEGMENT|12130,12133|false|false|false|C0032520;C3853643|Polymerase Chain Reaction;Probe with target amplification technique|PCR
Event|Event|SIMPLE_SEGMENT|12138,12146|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|12138,12146|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|12138,12146|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|12138,12146|false|false|false|C5237010|Expression Negative|negative
Event|Event|SIMPLE_SEGMENT|12154,12158|false|false|false|||last
Event|Event|SIMPLE_SEGMENT|12160,12175|false|false|false|||hospitalization
Procedure|Health Care Activity|SIMPLE_SEGMENT|12160,12175|false|false|false|C0019993|Hospitalization|hospitalization
Event|Event|SIMPLE_SEGMENT|12181,12190|false|false|false|||completed
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12198,12208|false|false|false|C0042313|vancomycin|vancomycin
Drug|Antibiotic|SIMPLE_SEGMENT|12198,12208|false|false|false|C0042313|vancomycin|vancomycin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12198,12208|false|false|false|C0489941|Vancomycin measurement|vancomycin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12232,12242|false|false|false|C0042313|vancomycin|vancomycin
Drug|Antibiotic|SIMPLE_SEGMENT|12232,12242|false|false|false|C0042313|vancomycin|vancomycin
Event|Event|SIMPLE_SEGMENT|12232,12242|false|false|false|||vancomycin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12232,12242|false|false|false|C0489941|Vancomycin measurement|vancomycin
Event|Event|SIMPLE_SEGMENT|12247,12256|false|false|false|||continued
Event|Event|SIMPLE_SEGMENT|12264,12279|false|false|false|||hospitalization
Procedure|Health Care Activity|SIMPLE_SEGMENT|12264,12279|false|false|false|C0019993|Hospitalization|hospitalization
Event|Event|SIMPLE_SEGMENT|12303,12312|false|false|false|||treatment
Finding|Conceptual Entity|SIMPLE_SEGMENT|12303,12312|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|SIMPLE_SEGMENT|12303,12312|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|SIMPLE_SEGMENT|12303,12312|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12303,12312|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Finding|Conceptual Entity|SIMPLE_SEGMENT|12324,12332|false|false|false|C2827424|Spectrum|spectrum
Drug|Antibiotic|SIMPLE_SEGMENT|12333,12344|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|SIMPLE_SEGMENT|12333,12344|false|false|false|||antibiotics
Drug|Antibiotic|SIMPLE_SEGMENT|12347,12352|false|false|false|C0250482|Zosyn|zosyn
Drug|Organic Chemical|SIMPLE_SEGMENT|12347,12352|false|false|false|C0250482|Zosyn|zosyn
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12358,12369|false|false|false|C0033817|Pseudomonas Infections|pseudomonas
Event|Event|SIMPLE_SEGMENT|12358,12369|false|false|false|||pseudomonas
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12370,12373|false|false|false|C0042029|Urinary tract infection|UTI
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12370,12373|false|false|false|C0077906|urinastatin|UTI
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12370,12373|false|false|false|C0077906|urinastatin|UTI
Event|Event|SIMPLE_SEGMENT|12370,12373|false|false|false|||UTI
Finding|Gene or Genome|SIMPLE_SEGMENT|12370,12373|false|false|false|C1412376;C5780748|AMBP gene;AMBP wt Allele|UTI
Drug|Antibiotic|SIMPLE_SEGMENT|12379,12384|false|false|false|C0250482|Zosyn|zosyn
Drug|Organic Chemical|SIMPLE_SEGMENT|12379,12384|false|false|false|C0250482|Zosyn|zosyn
Event|Event|SIMPLE_SEGMENT|12389,12398|false|false|false|||completed
Event|Event|SIMPLE_SEGMENT|12415,12424|false|false|false|||continued
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12428,12433|false|false|false|C0042313|vancomycin|vanco
Drug|Antibiotic|SIMPLE_SEGMENT|12428,12433|false|false|false|C0042313|vancomycin|vanco
Event|Event|SIMPLE_SEGMENT|12428,12433|false|false|false|||vanco
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12450,12456|false|false|false|C0002871|Anemia|Anemia
Event|Event|SIMPLE_SEGMENT|12450,12456|false|false|false|||Anemia
Event|Event|SIMPLE_SEGMENT|12458,12465|false|false|false|||Patient
Finding|Body Substance|SIMPLE_SEGMENT|12458,12465|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|12458,12465|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|12458,12465|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|12471,12477|false|false|false|C0018302|guaiac|guaiac
Drug|Organic Chemical|SIMPLE_SEGMENT|12471,12477|false|false|false|C0018302|guaiac|guaiac
Event|Event|SIMPLE_SEGMENT|12471,12477|false|false|false|||guaiac
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|12471,12486|false|false|false|C0744492|guaiac positive|guaiac positive
Finding|Finding|SIMPLE_SEGMENT|12471,12493|false|false|false|C0266813||guaiac positive stools
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|12478,12486|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Event|Event|SIMPLE_SEGMENT|12478,12486|false|false|false|||positive
Finding|Classification|SIMPLE_SEGMENT|12478,12486|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|SIMPLE_SEGMENT|12478,12486|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12487,12493|false|false|false|C0489144||stools
Event|Event|SIMPLE_SEGMENT|12487,12493|false|false|false|||stools
Finding|Body Substance|SIMPLE_SEGMENT|12487,12493|false|false|false|C0015733|Feces|stools
Event|Event|SIMPLE_SEGMENT|12507,12516|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|12507,12516|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|12518,12521|false|false|false|||new
Finding|Finding|SIMPLE_SEGMENT|12518,12521|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|12518,12521|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Event|Event|SIMPLE_SEGMENT|12532,12541|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|12532,12541|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12543,12546|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12543,12546|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Event|Event|SIMPLE_SEGMENT|12547,12553|false|false|false|||stable
Finding|Intellectual Product|SIMPLE_SEGMENT|12547,12553|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|SIMPLE_SEGMENT|12558,12562|false|false|false|||high
Finding|Finding|SIMPLE_SEGMENT|12558,12562|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|SIMPLE_SEGMENT|12558,12562|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|SIMPLE_SEGMENT|12558,12562|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Event|Event|SIMPLE_SEGMENT|12579,12594|false|false|false|||hospitalization
Procedure|Health Care Activity|SIMPLE_SEGMENT|12579,12594|false|false|false|C0019993|Hospitalization|hospitalization
Event|Event|SIMPLE_SEGMENT|12604,12611|false|false|false|||receive
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|12631,12638|false|false|false|C0009361|Colloids|colloid
Event|Event|SIMPLE_SEGMENT|12631,12638|false|false|false|||colloid
Finding|Body Substance|SIMPLE_SEGMENT|12631,12638|false|false|false|C1527250|Colloid, body substance|colloid
Event|Event|SIMPLE_SEGMENT|12639,12647|false|false|false|||pressure
Finding|Finding|SIMPLE_SEGMENT|12639,12647|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|12639,12647|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|12639,12647|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|12639,12647|false|false|false|C0033095||pressure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12639,12655|false|false|false|C0419008|pressure support|pressure support
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12648,12655|false|false|false|C1317973|Support - dental|support
Drug|Organic Chemical|SIMPLE_SEGMENT|12648,12655|false|false|false|C1171411|Support brand of multivitamin|support
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12648,12655|false|false|false|C1171411|Support brand of multivitamin|support
Drug|Vitamin|SIMPLE_SEGMENT|12648,12655|false|false|false|C1171411|Support brand of multivitamin|support
Event|Event|SIMPLE_SEGMENT|12648,12655|false|false|false|||support
Finding|Conceptual Entity|SIMPLE_SEGMENT|12648,12655|false|false|false|C1521721|Supportive assistance|support
Procedure|Health Care Activity|SIMPLE_SEGMENT|12648,12655|false|false|false|C0344211|Supportive care|support
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12661,12675|false|false|false|C0020676|Hypothyroidism|Hypothyroidism
Event|Event|SIMPLE_SEGMENT|12661,12675|false|false|false|||Hypothyroidism
Event|Event|SIMPLE_SEGMENT|12677,12686|false|false|false|||Continued
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12690,12703|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Hormone|SIMPLE_SEGMENT|12690,12703|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Organic Chemical|SIMPLE_SEGMENT|12690,12703|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12690,12703|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Event|Event|SIMPLE_SEGMENT|12690,12703|false|false|false|||levothyroxine
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12722,12726|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|SIMPLE_SEGMENT|12722,12726|false|false|false|||GERD
Finding|Body Substance|SIMPLE_SEGMENT|12728,12735|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|12728,12735|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|12728,12735|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Organic Chemical|SIMPLE_SEGMENT|12750,12760|false|false|false|C0028978|omeprazole|omeprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12750,12760|false|false|false|C0028978|omeprazole|omeprazole
Event|Event|SIMPLE_SEGMENT|12766,12781|false|false|false|||hospitalization
Procedure|Health Care Activity|SIMPLE_SEGMENT|12766,12781|false|false|false|C0019993|Hospitalization|hospitalization
Event|Event|SIMPLE_SEGMENT|12794,12801|false|false|false|||stopped
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|12826,12834|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Event|Event|SIMPLE_SEGMENT|12826,12834|false|false|false|||positive
Finding|Classification|SIMPLE_SEGMENT|12826,12834|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|SIMPLE_SEGMENT|12826,12834|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Event|Event|SIMPLE_SEGMENT|12849,12861|false|false|false|||transitioned
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12865,12875|false|false|false|C0019593|Histamine H2 Antagonists|H2 blocker
Event|Event|SIMPLE_SEGMENT|12868,12875|false|false|false|||blocker
Event|Event|SIMPLE_SEGMENT|12883,12894|false|false|false|||prophylaxis
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12883,12894|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Event|Event|SIMPLE_SEGMENT|12905,12909|false|false|false|||held
Event|Event|SIMPLE_SEGMENT|12915,12922|false|false|false|||setting
Finding|Mental Process|SIMPLE_SEGMENT|12915,12922|false|false|false|C0542559|contextual factors|setting
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|12926,12934|false|false|false|C0011206|Delirium|delirium
Event|Event|SIMPLE_SEGMENT|12926,12934|false|false|false|||delirium
Drug|Organic Chemical|SIMPLE_SEGMENT|12936,12946|false|false|false|C0015620|famotidine|Famotidine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12936,12946|false|false|false|C0015620|famotidine|Famotidine
Event|Event|SIMPLE_SEGMENT|12936,12946|false|false|false|||Famotidine
Event|Event|SIMPLE_SEGMENT|12951,12960|false|false|false|||restarted
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|12969,12972|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12969,12972|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12969,12972|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|12969,12972|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|12969,12972|false|false|false|C1332410|BID gene|BID
Finding|Intellectual Product|SIMPLE_SEGMENT|12973,12977|false|false|false|C1720092|Once - dosing instruction fragment|once
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|12997,13006|true|false|false|C0011206|Delirium|delirious
Event|Event|SIMPLE_SEGMENT|12997,13006|true|false|false|||delirious
Event|Event|SIMPLE_SEGMENT|13012,13015|false|false|false|||EKG
Finding|Intellectual Product|SIMPLE_SEGMENT|13012,13015|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|13012,13015|false|false|false|C1623258|Electrocardiography|EKG
Event|Event|SIMPLE_SEGMENT|13016,13023|false|false|false|||Changes
Finding|Functional Concept|SIMPLE_SEGMENT|13016,13023|false|false|false|C0392747|Changing|Changes
Finding|Body Substance|SIMPLE_SEGMENT|13025,13032|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|13025,13032|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|13025,13032|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|13045,13048|false|false|false|||STE
Finding|Gene or Genome|SIMPLE_SEGMENT|13045,13048|false|false|false|C1420459;C3811127|SULT1E1 gene;SULT1E1 wt Allele|STE
Event|Event|SIMPLE_SEGMENT|13060,13068|false|false|false|||elevated
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13070,13078|false|false|false|C0041199|Troponin|troponin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|13070,13078|false|false|false|C0041199|Troponin|troponin
Event|Event|SIMPLE_SEGMENT|13070,13078|false|false|false|||troponin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|13070,13078|false|false|false|C0523952|Troponin measurement|troponin
Event|Event|SIMPLE_SEGMENT|13097,13106|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|13097,13106|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|13108,13112|false|false|false|||felt
Finding|Finding|SIMPLE_SEGMENT|13113,13119|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|13113,13119|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|13134,13140|false|false|false|C3263722;C3263723|Traumatic AND/OR non-traumatic injury;Traumatic injury|injury
Event|Event|SIMPLE_SEGMENT|13134,13140|false|false|false|||injury
Event|Event|SIMPLE_SEGMENT|13145,13157|false|false|false|||compressions
Finding|Functional Concept|SIMPLE_SEGMENT|13145,13157|false|false|false|C0332459|Compressed structure|compressions
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|13145,13157|false|false|false|C0728907|Compression|compressions
Event|Event|SIMPLE_SEGMENT|13162,13164|false|false|false|||ED
Event|Event|SIMPLE_SEGMENT|13169,13175|false|false|false|||demand
Finding|Idea or Concept|SIMPLE_SEGMENT|13169,13175|false|false|false|C0699784|Economic demand|demand
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|13169,13175|false|false|false|C0441516|Demand (clinical)|demand
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13169,13184|false|false|false|C4049375|Ischemia co-occurrent and due to increased oxygen demand|demand ischemia
Event|Event|SIMPLE_SEGMENT|13176,13184|false|false|false|||ischemia
Finding|Pathologic Function|SIMPLE_SEGMENT|13176,13184|false|false|false|C0022116|Ischemia|ischemia
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|13176,13184|false|false|false|C4321499|Ischemia Procedure|ischemia
Finding|Body Substance|SIMPLE_SEGMENT|13199,13206|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|13199,13206|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|13199,13206|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|13211,13218|false|false|false|C0015811|Femur|femoral
Event|Event|SIMPLE_SEGMENT|13226,13232|false|false|false|||placed
Event|Event|SIMPLE_SEGMENT|13244,13251|false|false|false|||setting
Finding|Mental Process|SIMPLE_SEGMENT|13244,13251|false|false|false|C0542559|contextual factors|setting
Event|Event|SIMPLE_SEGMENT|13260,13271|false|false|false|||hypotension
Finding|Finding|SIMPLE_SEGMENT|13260,13271|false|false|false|C0020649|Hypotension|hypotension
Event|Event|SIMPLE_SEGMENT|13282,13294|false|false|false|||discontinued
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|13299,13302|false|false|false|C0228479|Structure of intraculminate fissure|ICU
Finding|Intellectual Product|SIMPLE_SEGMENT|13299,13302|false|false|false|C4554035|Inventory of Callous-Unemotional Traits|ICU
Event|Event|SIMPLE_SEGMENT|13307,13315|false|false|false|||replaced
Event|Event|SIMPLE_SEGMENT|13322,13326|false|false|false|||PICC
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|13322,13326|false|false|false|C2049629|Peripherally Inserted Central Catheter Line Insertion|PICC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13340,13343|false|false|false|C1137947|SET protein, human|set
Drug|Biologically Active Substance|SIMPLE_SEGMENT|13340,13343|false|false|false|C1137947|SET protein, human|set
Event|Event|SIMPLE_SEGMENT|13340,13343|false|false|false|||set
Finding|Conceptual Entity|SIMPLE_SEGMENT|13340,13343|false|false|false|C0036849;C1366517;C1442518;C1552652;C1705195|Parameterized Data Type - Set;SET gene;Set (Psychology);Set scale;set (group)|set
Finding|Functional Concept|SIMPLE_SEGMENT|13340,13343|false|false|false|C0036849;C1366517;C1442518;C1552652;C1705195|Parameterized Data Type - Set;SET gene;Set (Psychology);Set scale;set (group)|set
Finding|Gene or Genome|SIMPLE_SEGMENT|13340,13343|false|false|false|C0036849;C1366517;C1442518;C1552652;C1705195|Parameterized Data Type - Set;SET gene;Set (Psychology);Set scale;set (group)|set
Finding|Idea or Concept|SIMPLE_SEGMENT|13340,13343|false|false|false|C0036849;C1366517;C1442518;C1552652;C1705195|Parameterized Data Type - Set;SET gene;Set (Psychology);Set scale;set (group)|set
Finding|Mental Process|SIMPLE_SEGMENT|13340,13343|false|false|false|C0036849;C1366517;C1442518;C1552652;C1705195|Parameterized Data Type - Set;SET gene;Set (Psychology);Set scale;set (group)|set
Event|Event|SIMPLE_SEGMENT|13357,13361|false|false|false|||grew
Finding|Finding|SIMPLE_SEGMENT|13377,13383|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|13377,13383|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Anatomy|Body System|SIMPLE_SEGMENT|13385,13389|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13385,13389|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|13385,13389|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Finding|Body Substance|SIMPLE_SEGMENT|13385,13389|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|SIMPLE_SEGMENT|13385,13389|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Drug|Substance|SIMPLE_SEGMENT|13390,13401|false|false|false|C2827365|Contaminant|contaminant
Event|Event|SIMPLE_SEGMENT|13390,13401|false|false|false|||contaminant
Event|Event|SIMPLE_SEGMENT|13409,13421|false|false|false|||surveillance
Event|Occupational Activity|SIMPLE_SEGMENT|13409,13421|false|false|false|C0684245|legal surveillance|surveillance
Finding|Functional Concept|SIMPLE_SEGMENT|13409,13421|false|false|false|C0220920|surveillance aspects|surveillance
Procedure|Health Care Activity|SIMPLE_SEGMENT|13409,13421|false|false|false|C0733511|Medical Surveillance|surveillance
Event|Event|SIMPLE_SEGMENT|13425,13433|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|13425,13433|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|13425,13433|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|13425,13433|false|false|false|C5237010|Expression Negative|negative
Finding|Idea or Concept|SIMPLE_SEGMENT|13438,13450|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Event|Event|SIMPLE_SEGMENT|13451,13457|false|false|false|||ISSUES
Event|Event|SIMPLE_SEGMENT|13461,13465|false|false|false|||Code
Event|Occupational Activity|SIMPLE_SEGMENT|13461,13465|false|false|false|C0009219|Coding|Code
Finding|Intellectual Product|SIMPLE_SEGMENT|13461,13465|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|Code
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|13474,13478|false|false|false|C0587081|Laboratory test finding|Labs
Event|Event|SIMPLE_SEGMENT|13504,13508|false|false|false|||chem
Finding|Functional Concept|SIMPLE_SEGMENT|13504,13508|false|false|false|C0079107|chemical aspects|chem
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|13504,13508|false|false|false|C0201682|Chemical procedure|chem
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|13504,13510|false|false|false|C2237045|Basic metabolic panel|chem 7
Event|Event|SIMPLE_SEGMENT|13548,13556|false|false|false|||diuresed
Event|Event|SIMPLE_SEGMENT|13559,13568|false|false|false|||Nutrition
Finding|Finding|SIMPLE_SEGMENT|13559,13568|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|Nutrition
Finding|Intellectual Product|SIMPLE_SEGMENT|13559,13568|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|Nutrition
Finding|Organism Function|SIMPLE_SEGMENT|13559,13568|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|Nutrition
Procedure|Research Activity|SIMPLE_SEGMENT|13559,13568|false|false|false|C0600072;C1521729|Feeding and dietary regimes;Nutritional Study|Nutrition
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|13559,13568|false|false|false|C0600072;C1521729|Feeding and dietary regimes;Nutritional Study|Nutrition
Finding|Functional Concept|SIMPLE_SEGMENT|13570,13574|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|Tube
Finding|Gene or Genome|SIMPLE_SEGMENT|13570,13574|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|Tube
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13583,13587|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|13583,13592|false|false|false|C0301569|Soft diet|soft diet
Drug|Food|SIMPLE_SEGMENT|13588,13592|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|SIMPLE_SEGMENT|13588,13592|false|false|false|||diet
Finding|Functional Concept|SIMPLE_SEGMENT|13588,13592|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|SIMPLE_SEGMENT|13588,13592|false|false|false|C0012159|Diet therapy|diet
Event|Event|SIMPLE_SEGMENT|13602,13609|false|false|false|||liqiuds
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13612,13623|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13612,13623|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|13612,13623|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|13612,13623|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|13612,13636|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|SIMPLE_SEGMENT|13627,13636|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|13627,13636|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Organic Chemical|SIMPLE_SEGMENT|13641,13652|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13641,13652|false|false|false|C0082607|fluticasone|fluticasone
Event|Event|SIMPLE_SEGMENT|13641,13652|false|false|false|||fluticasone
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13670,13675|false|false|false|C1154182|Spray Dosage Form|Spray
Event|Activity|SIMPLE_SEGMENT|13670,13675|false|false|false|C2003858|Spray (action)|Spray
Event|Event|SIMPLE_SEGMENT|13670,13675|false|false|false|||Spray
Finding|Functional Concept|SIMPLE_SEGMENT|13670,13675|false|false|false|C4521772|Spray (administration method)|Spray
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13670,13687|false|false|false|C1710170|SPRAY, SUSPENSION|Spray, Suspension
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13677,13687|false|false|false|C0038960;C1382107|Suspension substance;Suspensions|Suspension
Drug|Substance|SIMPLE_SEGMENT|13677,13687|false|false|false|C0038960;C1382107|Suspension substance;Suspensions|Suspension
Event|Event|SIMPLE_SEGMENT|13677,13687|false|false|false|||Suspension
Finding|Functional Concept|SIMPLE_SEGMENT|13677,13687|false|false|false|C1705537|Suspension (action)|Suspension
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|13698,13701|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13698,13701|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|13698,13701|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|13698,13701|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|13698,13701|false|false|false|C1332410|BID gene|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13706,13719|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Hormone|SIMPLE_SEGMENT|13706,13719|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Organic Chemical|SIMPLE_SEGMENT|13706,13719|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13706,13719|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Event|Event|SIMPLE_SEGMENT|13706,13719|false|false|false|||levothyroxine
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13727,13733|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|13727,13733|false|false|false|||Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13747,13753|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|13747,13753|false|false|false|||Tablet
Drug|Organic Chemical|SIMPLE_SEGMENT|13768,13781|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13768,13781|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Event|Event|SIMPLE_SEGMENT|13768,13781|false|false|false|||acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|13768,13781|false|false|false|C0373527|Acetaminophen measurement|acetaminophen
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13789,13795|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13805,13812|false|false|false|C0039225|Tablet Dosage Form|Tablets
Event|Event|SIMPLE_SEGMENT|13805,13812|false|false|false|||Tablets
Finding|Gene or Genome|SIMPLE_SEGMENT|13819,13822|false|false|false|C1422467|CIAO3 gene|prn
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13826,13835|false|false|false|C0032629|Polyvinyls|polyvinyl
Drug|Organic Chemical|SIMPLE_SEGMENT|13826,13835|false|false|false|C0032629|Polyvinyls|polyvinyl
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13826,13843|false|false|false|C0032623|polyvinyl alcohol|polyvinyl alcohol
Drug|Organic Chemical|SIMPLE_SEGMENT|13836,13843|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13836,13843|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Event|Event|SIMPLE_SEGMENT|13836,13843|false|false|false|||alcohol
Finding|Intellectual Product|SIMPLE_SEGMENT|13836,13843|false|false|false|C1547288|Alcohol - Recreational Drug Use Code|alcohol
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13850,13855|false|false|false|C0991568|Drops - Drug Form|Drops
Event|Event|SIMPLE_SEGMENT|13850,13855|false|false|false|||Drops
Finding|Gene or Genome|SIMPLE_SEGMENT|13878,13881|false|false|false|C1422467|CIAO3 gene|prn
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13885,13892|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|13885,13892|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13885,13892|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|13885,13892|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|13885,13892|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|13885,13892|false|false|false|C0202098|Insulin measurement|insulin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13885,13899|true|false|false|C0293359|insulin lispro|insulin lispro
Drug|Hormone|SIMPLE_SEGMENT|13885,13899|true|false|false|C0293359|insulin lispro|insulin lispro
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13885,13899|true|false|false|C0293359|insulin lispro|insulin lispro
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13893,13899|false|false|false|C0293359|insulin lispro|lispro
Drug|Hormone|SIMPLE_SEGMENT|13893,13899|false|false|false|C0293359|insulin lispro|lispro
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13893,13899|false|false|false|C0293359|insulin lispro|lispro
Event|Event|SIMPLE_SEGMENT|13893,13899|false|false|false|||lispro
Event|Event|SIMPLE_SEGMENT|13904,13908|false|false|false|||unit
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13912,13920|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|Solution
Drug|Substance|SIMPLE_SEGMENT|13912,13920|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|Solution
Event|Event|SIMPLE_SEGMENT|13912,13920|false|false|false|||Solution
Finding|Conceptual Entity|SIMPLE_SEGMENT|13912,13920|false|false|false|C2699488|Resolution|Solution
Event|Event|SIMPLE_SEGMENT|13924,13927|false|false|false|||TID
Finding|Functional Concept|SIMPLE_SEGMENT|13928,13935|false|false|false|C0332246|Sliding|Sliding
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|13928,13941|false|false|false|C2937251|sliding scale|Sliding scale
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|13936,13941|false|false|false|C0222045|Integumentary scale|scale
Event|Activity|SIMPLE_SEGMENT|13936,13941|false|false|false|C1947916|Scaling|scale
Event|Event|SIMPLE_SEGMENT|13936,13941|false|false|false|||scale
Finding|Conceptual Entity|SIMPLE_SEGMENT|13936,13941|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Finding|Intellectual Product|SIMPLE_SEGMENT|13936,13941|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|scale
Finding|Functional Concept|SIMPLE_SEGMENT|13950,13962|false|false|false|C1522438|Subcutaneous Route of Administration|Subcutaneous
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13969,13974|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|SIMPLE_SEGMENT|13977,13980|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|13977,13980|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|14105,14109|false|false|false|||call
Finding|Functional Concept|SIMPLE_SEGMENT|14105,14109|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Gene or Genome|SIMPLE_SEGMENT|14105,14109|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Intellectual Product|SIMPLE_SEGMENT|14105,14109|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Mental Process|SIMPLE_SEGMENT|14105,14109|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Drug|Organic Chemical|SIMPLE_SEGMENT|14119,14129|false|false|false|C0025942|miconazole|miconazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14119,14129|false|false|false|C0025942|miconazole|miconazole
Event|Event|SIMPLE_SEGMENT|14119,14129|false|false|false|||miconazole
Drug|Organic Chemical|SIMPLE_SEGMENT|14119,14137|false|false|false|C0086620|miconazole nitrate|miconazole nitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14119,14137|false|false|false|C0086620|miconazole nitrate|miconazole nitrate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|14130,14137|false|false|false|C0028125;C0699857;C3848573|Nitrate;Nitrates;nitrate ion|nitrate
Drug|Inorganic Chemical|SIMPLE_SEGMENT|14130,14137|false|false|false|C0028125;C0699857;C3848573|Nitrate;Nitrates;nitrate ion|nitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14130,14137|false|false|false|C0028125;C0699857;C3848573|Nitrate;Nitrates;nitrate ion|nitrate
Event|Event|SIMPLE_SEGMENT|14130,14137|false|false|false|||nitrate
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|14142,14148|false|false|false|C0032861;C1382110|Powder dose form;powder physical state|Powder
Drug|Substance|SIMPLE_SEGMENT|14142,14148|false|false|false|C0032861;C1382110|Powder dose form;powder physical state|Powder
Event|Event|SIMPLE_SEGMENT|14151,14154|false|false|false|||TID
Finding|Gene or Genome|SIMPLE_SEGMENT|14155,14158|false|false|false|C1422467|CIAO3 gene|prn
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14159,14163|false|false|false|C5779629|Eruption of skin (disorder)|rash
Event|Event|SIMPLE_SEGMENT|14159,14163|false|false|false|||rash
Finding|Pathologic Function|SIMPLE_SEGMENT|14159,14163|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|SIMPLE_SEGMENT|14159,14163|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|14167,14177|false|false|false|C0042313|vancomycin|vancomycin
Drug|Antibiotic|SIMPLE_SEGMENT|14167,14177|false|false|false|C0042313|vancomycin|vancomycin
Event|Event|SIMPLE_SEGMENT|14167,14177|false|false|false|||vancomycin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|14167,14177|false|false|false|C0489941|Vancomycin measurement|vancomycin
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|14185,14192|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|SIMPLE_SEGMENT|14185,14192|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|14185,14192|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Event|Event|SIMPLE_SEGMENT|14198,14201|false|false|false|||Q6H
Drug|Biologically Active Substance|SIMPLE_SEGMENT|14216,14223|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|SIMPLE_SEGMENT|14216,14223|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14216,14223|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Event|Event|SIMPLE_SEGMENT|14216,14223|false|false|false|||heparin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|14216,14233|false|false|false|C0770546|heparin, porcine|heparin (porcine)
Drug|Organic Chemical|SIMPLE_SEGMENT|14216,14233|false|false|false|C0770546|heparin, porcine|heparin (porcine)
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14216,14233|false|false|false|C0770546|heparin, porcine|heparin (porcine)
Event|Event|SIMPLE_SEGMENT|14225,14232|false|false|false|||porcine
Finding|Finding|SIMPLE_SEGMENT|14225,14232|false|false|false|C4554819|Porcine prosthetic valve|porcine
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|14248,14256|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|Solution
Drug|Substance|SIMPLE_SEGMENT|14248,14256|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|Solution
Event|Event|SIMPLE_SEGMENT|14248,14256|false|false|false|||Solution
Finding|Conceptual Entity|SIMPLE_SEGMENT|14248,14256|false|false|false|C2699488|Resolution|Solution
Drug|Organic Chemical|SIMPLE_SEGMENT|14276,14285|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14276,14285|false|false|false|C0001927|albuterol|albuterol
Event|Event|SIMPLE_SEGMENT|14276,14285|false|false|false|||albuterol
Drug|Organic Chemical|SIMPLE_SEGMENT|14276,14293|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14276,14293|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|14286,14293|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|SIMPLE_SEGMENT|14286,14293|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14286,14293|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Event|Event|SIMPLE_SEGMENT|14286,14293|false|false|false|||sulfate
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|14317,14325|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|Solution
Drug|Substance|SIMPLE_SEGMENT|14317,14325|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|Solution
Event|Event|SIMPLE_SEGMENT|14317,14325|false|false|false|||Solution
Finding|Conceptual Entity|SIMPLE_SEGMENT|14317,14325|false|false|false|C2699488|Resolution|Solution
Finding|Gene or Genome|SIMPLE_SEGMENT|14333,14336|false|false|false|C1422467|CIAO3 gene|prn
Event|Event|SIMPLE_SEGMENT|14338,14341|false|false|false|||SOB
Finding|Sign or Symptom|SIMPLE_SEGMENT|14338,14341|false|false|false|C0013404|Dyspnea|SOB
Drug|Organic Chemical|SIMPLE_SEGMENT|14346,14357|false|false|false|C0027235|ipratropium|ipratropium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14346,14357|false|false|false|C0027235|ipratropium|ipratropium
Drug|Organic Chemical|SIMPLE_SEGMENT|14346,14365|false|false|false|C0700580|ipratropium bromide|ipratropium bromide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14346,14365|false|false|false|C0700580|ipratropium bromide|ipratropium bromide
Drug|Inorganic Chemical|SIMPLE_SEGMENT|14358,14365|false|false|false|C0006222|Bromides|bromide
Event|Event|SIMPLE_SEGMENT|14358,14365|false|false|false|||bromide
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|14358,14365|false|false|false|C0202341|Bromides measurement|bromide
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|14373,14381|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|Solution
Drug|Substance|SIMPLE_SEGMENT|14373,14381|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|Solution
Event|Event|SIMPLE_SEGMENT|14373,14381|false|false|false|||Solution
Finding|Conceptual Entity|SIMPLE_SEGMENT|14373,14381|false|false|false|C2699488|Resolution|Solution
Event|Event|SIMPLE_SEGMENT|14384,14388|false|false|false|||q6hr
Finding|Gene or Genome|SIMPLE_SEGMENT|14389,14392|false|false|false|C1422467|CIAO3 gene|prn
Event|Event|SIMPLE_SEGMENT|14393,14396|false|false|false|||SOB
Finding|Sign or Symptom|SIMPLE_SEGMENT|14393,14396|false|false|false|C0013404|Dyspnea|SOB
Event|Event|SIMPLE_SEGMENT|14399,14408|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|14399,14408|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|14399,14408|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|14399,14408|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|14399,14408|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|14399,14420|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14409,14420|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14409,14420|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|14409,14420|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|14409,14420|false|false|false|C4284232|Medications|Medications
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|14425,14435|false|false|false|C0042313|vancomycin|Vancomycin
Drug|Antibiotic|SIMPLE_SEGMENT|14425,14435|false|false|false|C0042313|vancomycin|Vancomycin
Event|Event|SIMPLE_SEGMENT|14425,14435|false|false|false|||Vancomycin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|14425,14435|false|false|false|C0489941|Vancomycin measurement|Vancomycin
Drug|Clinical Drug|SIMPLE_SEGMENT|14425,14440|false|false|false|C0360373||Vancomycin Oral
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|14436,14440|false|false|false|C0226896|Oral cavity|Oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|14436,14440|false|false|false|C1272919|Oral Dosage Form|Oral
Finding|Finding|SIMPLE_SEGMENT|14436,14440|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Finding|Functional Concept|SIMPLE_SEGMENT|14436,14440|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|14436,14447|false|false|false|C1273619|Oral Liquid Product|Oral Liquid
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|14441,14447|false|false|false|C0302908;C1697794|Liquid Dosage Form;Liquid substance|Liquid
Drug|Substance|SIMPLE_SEGMENT|14441,14447|false|false|false|C0302908;C1697794|Liquid Dosage Form;Liquid substance|Liquid
Event|Event|SIMPLE_SEGMENT|14441,14447|false|false|false|||Liquid
Finding|Finding|SIMPLE_SEGMENT|14441,14447|false|false|false|C1304698|Liquid (finding)|Liquid
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|14441,14447|false|false|false|C0301571|Liquid diet|Liquid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14462,14470|false|false|false|C0720099|Duration brand of oxymetazoline|Duration
Event|Event|SIMPLE_SEGMENT|14462,14470|false|false|false|||Duration
Event|Event|SIMPLE_SEGMENT|14486,14489|false|false|false|||day
Finding|Idea or Concept|SIMPLE_SEGMENT|14486,14489|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|14486,14489|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|SIMPLE_SEGMENT|14500,14511|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14500,14511|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|SIMPLE_SEGMENT|14500,14511|false|false|false|||Fluticasone
Drug|Organic Chemical|SIMPLE_SEGMENT|14500,14522|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14500,14522|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|SIMPLE_SEGMENT|14512,14522|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Event|Event|SIMPLE_SEGMENT|14532,14536|false|false|false|||PUFF
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|14540,14543|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|14540,14543|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|14540,14543|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|14540,14543|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|14540,14543|false|false|false|C1332410|BID gene|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|14548,14561|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Hormone|SIMPLE_SEGMENT|14548,14561|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Organic Chemical|SIMPLE_SEGMENT|14548,14561|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14548,14561|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Event|Event|SIMPLE_SEGMENT|14548,14561|false|false|false|||Levothyroxine
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|14548,14568|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Hormone|SIMPLE_SEGMENT|14548,14568|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14548,14568|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|14562,14568|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|14562,14568|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14562,14568|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|14562,14568|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|14562,14568|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|14562,14568|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Organic Chemical|SIMPLE_SEGMENT|14589,14602|false|false|false|C0040864|triamcinolone|Triamcinolone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14589,14602|false|false|false|C0040864|triamcinolone|Triamcinolone
Drug|Organic Chemical|SIMPLE_SEGMENT|14589,14612|false|false|false|C0040866|triamcinolone acetonide|Triamcinolone Acetonide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14589,14612|false|false|false|C0040866|triamcinolone acetonide|Triamcinolone Acetonide
Event|Event|SIMPLE_SEGMENT|14603,14612|false|false|false|||Acetonide
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|14620,14625|false|false|false|C0700385;C0705539;C1378128|Cream;Dairy Cream;Emollient Cream|Cream
Drug|Food|SIMPLE_SEGMENT|14620,14625|false|false|false|C0700385;C0705539;C1378128|Cream;Dairy Cream;Emollient Cream|Cream
Finding|Gene or Genome|SIMPLE_SEGMENT|14628,14632|false|false|false|C1858559|APPL1 gene|Appl
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|14636,14639|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|14636,14639|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|14636,14639|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|14636,14639|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|14636,14639|false|false|false|C1332410|BID gene|BID
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14641,14644|false|false|false|C0030360;C0154682;C0205825|Lateral Sclerosis;Liposarcoma, Pleomorphic;Papillon-Lefevre Disease|pls
Disorder|Neoplastic Process|SIMPLE_SEGMENT|14641,14644|false|false|false|C0030360;C0154682;C0205825|Lateral Sclerosis;Liposarcoma, Pleomorphic;Papillon-Lefevre Disease|pls
Event|Event|SIMPLE_SEGMENT|14641,14644|false|false|false|||pls
Finding|Gene or Genome|SIMPLE_SEGMENT|14641,14644|false|false|false|C1413811;C5849001|CTSC gene;CTSC wt Allele|pls
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|14656,14661|false|false|false|C0934502|anatomical layer|layer
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14665,14669|false|false|false|C5779629|Eruption of skin (disorder)|rash
Event|Event|SIMPLE_SEGMENT|14665,14669|false|false|false|||rash
Finding|Pathologic Function|SIMPLE_SEGMENT|14665,14669|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|SIMPLE_SEGMENT|14665,14669|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Drug|Organic Chemical|SIMPLE_SEGMENT|14674,14684|false|false|false|C0025942|miconazole|Miconazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14674,14684|false|false|false|C0025942|miconazole|Miconazole
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|14685,14691|false|false|false|C0032861;C1382110|Powder dose form;powder physical state|Powder
Drug|Substance|SIMPLE_SEGMENT|14685,14691|false|false|false|C0032861;C1382110|Powder dose form;powder physical state|Powder
Event|Event|SIMPLE_SEGMENT|14685,14691|false|false|false|||Powder
Finding|Gene or Genome|SIMPLE_SEGMENT|14697,14701|false|false|false|C1858559|APPL1 gene|Appl
Event|Event|SIMPLE_SEGMENT|14705,14708|false|false|false|||TID
Anatomy|Body Location or Region|SIMPLE_SEGMENT|14713,14718|false|false|false|C0018246;C0816951;C4266533|Inguinal part of abdomen;Inguinal region;Pelvis>Groin|groin
Finding|Finding|SIMPLE_SEGMENT|14713,14723|false|false|false|C0239785|Rash of groin|groin rash
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14719,14723|false|false|false|C5779629|Eruption of skin (disorder)|rash
Event|Event|SIMPLE_SEGMENT|14719,14723|false|false|false|||rash
Finding|Pathologic Function|SIMPLE_SEGMENT|14719,14723|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|SIMPLE_SEGMENT|14719,14723|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|14728,14735|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Hormone|SIMPLE_SEGMENT|14728,14735|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14728,14735|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Event|Event|SIMPLE_SEGMENT|14728,14735|false|false|false|||Insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|14728,14735|false|false|false|C1337112|INS gene|Insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|14728,14735|false|false|false|C0202098|Insulin measurement|Insulin
Finding|Functional Concept|SIMPLE_SEGMENT|14746,14753|false|false|false|C0332246|Sliding|Sliding
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|14746,14759|false|false|false|C2937251|sliding scale|Sliding Scale
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|14754,14759|false|false|false|C0222045|Integumentary scale|Scale
Event|Activity|SIMPLE_SEGMENT|14754,14759|false|false|false|C1947916|Scaling|Scale
Finding|Conceptual Entity|SIMPLE_SEGMENT|14754,14759|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|Scale
Finding|Intellectual Product|SIMPLE_SEGMENT|14754,14759|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|Scale
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|14779,14786|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Hormone|SIMPLE_SEGMENT|14779,14786|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14779,14786|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Event|Event|SIMPLE_SEGMENT|14779,14786|false|false|false|||Insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|14779,14786|false|false|false|C1337112|INS gene|Insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|14779,14786|false|false|false|C0202098|Insulin measurement|Insulin
Finding|Functional Concept|SIMPLE_SEGMENT|14790,14797|false|false|false|C0332246|Sliding|Sliding
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|14790,14803|false|false|false|C2937251|sliding scale|Sliding Scale
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|14798,14803|false|false|false|C0222045|Integumentary scale|Scale
Event|Activity|SIMPLE_SEGMENT|14798,14803|false|false|false|C1947916|Scaling|Scale
Finding|Conceptual Entity|SIMPLE_SEGMENT|14798,14803|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|Scale
Finding|Intellectual Product|SIMPLE_SEGMENT|14798,14803|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|Scale
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|14810,14816|false|false|false|C0293359|insulin lispro|lispro
Drug|Hormone|SIMPLE_SEGMENT|14810,14816|false|false|false|C0293359|insulin lispro|lispro
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14810,14816|false|false|false|C0293359|insulin lispro|lispro
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|14810,14824|false|false|false|C0293359|insulin lispro|lispro Insulin
Drug|Hormone|SIMPLE_SEGMENT|14810,14824|false|false|false|C0293359|insulin lispro|lispro Insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14810,14824|false|false|false|C0293359|insulin lispro|lispro Insulin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|14817,14824|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Hormone|SIMPLE_SEGMENT|14817,14824|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14817,14824|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Event|Event|SIMPLE_SEGMENT|14817,14824|false|false|false|||Insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|14817,14824|false|false|false|C1337112|INS gene|Insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|14817,14824|false|false|false|C0202098|Insulin measurement|Insulin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|14828,14838|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14828,14838|false|false|false|C0065374|lisinopril|Lisinopril
Event|Activity|SIMPLE_SEGMENT|14854,14858|false|false|false|C1948035|Hold (action)|HOLD
Event|Event|SIMPLE_SEGMENT|14854,14858|false|false|false|||HOLD
Finding|Functional Concept|SIMPLE_SEGMENT|14854,14858|false|false|false|C1553387;C3853841|Hold - dosing instruction fragment;hold - Data Operation|HOLD
Finding|Intellectual Product|SIMPLE_SEGMENT|14854,14858|false|false|false|C1553387;C3853841|Hold - dosing instruction fragment;hold - Data Operation|HOLD
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14863,14866|false|false|false|C0871470|Systolic Pressure|SBP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|14863,14866|false|false|false|C0085805|Androgen Binding Protein|SBP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|14863,14866|false|false|false|C0085805|Androgen Binding Protein|SBP
Event|Event|SIMPLE_SEGMENT|14863,14866|false|false|false|||SBP
Finding|Gene or Genome|SIMPLE_SEGMENT|14863,14866|false|false|false|C1705296;C3274833|CCHCR1 wt Allele;SHBG wt Allele|SBP
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|14863,14866|false|false|false|C1306620|Systolic blood pressure measurement|SBP
Drug|Organic Chemical|SIMPLE_SEGMENT|14875,14885|false|false|false|C0015620|famotidine|Famotidine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14875,14885|false|false|false|C0015620|famotidine|Famotidine
Drug|Biologically Active Substance|SIMPLE_SEGMENT|14904,14911|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Drug|Organic Chemical|SIMPLE_SEGMENT|14904,14911|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14904,14911|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Event|Event|SIMPLE_SEGMENT|14917,14921|false|false|false|||UNIT
Event|Event|SIMPLE_SEGMENT|14925,14928|false|false|false|||TID
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|14934,14943|false|false|false|C0032629|Polyvinyls|polyvinyl
Drug|Organic Chemical|SIMPLE_SEGMENT|14934,14943|false|false|false|C0032629|Polyvinyls|polyvinyl
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|14934,14951|false|false|false|C0032623|polyvinyl alcohol|polyvinyl alcohol
Drug|Organic Chemical|SIMPLE_SEGMENT|14944,14951|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14944,14951|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Event|Event|SIMPLE_SEGMENT|14944,14951|false|false|false|||alcohol
Finding|Intellectual Product|SIMPLE_SEGMENT|14944,14951|false|false|false|C1547288|Alcohol - Recreational Drug Use Code|alcohol
Finding|Gene or Genome|SIMPLE_SEGMENT|14976,14979|false|false|false|C1422467|CIAO3 gene|PRN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14980,14988|false|false|false|C0013238;C0022575|Dry Eye Syndromes;Keratoconjunctivitis Sicca|dry eyes
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14980,14988|false|false|false|C0720056|Dry Eyes brand of ocular lubricant|dry eyes
Finding|Sign or Symptom|SIMPLE_SEGMENT|14980,14988|false|false|false|C0314719|Dryness of eye|dry eyes
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|14984,14988|false|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14984,14988|false|false|false|C5848506||eyes
Event|Event|SIMPLE_SEGMENT|14984,14988|false|false|false|||eyes
Drug|Organic Chemical|SIMPLE_SEGMENT|14994,15002|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14994,15002|false|false|false|C1692318|docusate|Docusate
Drug|Organic Chemical|SIMPLE_SEGMENT|14994,15009|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14994,15009|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|15003,15009|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|15003,15009|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15003,15009|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|15003,15009|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|15003,15009|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|15003,15009|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|15011,15017|false|false|false|C0302908;C1697794|Liquid Dosage Form;Liquid substance|Liquid
Drug|Substance|SIMPLE_SEGMENT|15011,15017|false|false|false|C0302908;C1697794|Liquid Dosage Form;Liquid substance|Liquid
Event|Event|SIMPLE_SEGMENT|15011,15017|false|false|false|||Liquid
Finding|Finding|SIMPLE_SEGMENT|15011,15017|false|false|false|C1304698|Liquid (finding)|Liquid
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|15011,15017|false|false|false|C0301571|Liquid diet|Liquid
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|15029,15032|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|15029,15032|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|15029,15032|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|15029,15032|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|15029,15032|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|15038,15048|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15038,15048|false|false|false|C0016860|furosemide|Furosemide
Event|Event|SIMPLE_SEGMENT|15068,15074|false|false|false|||needed
Finding|Intellectual Product|SIMPLE_SEGMENT|15079,15085|false|false|false|C1705102|Volume (publication)|volume
Finding|Pathologic Function|SIMPLE_SEGMENT|15079,15094|false|false|false|C0546817|Hypervolemia (finding)|volume overload
Event|Event|SIMPLE_SEGMENT|15086,15094|false|false|false|||overload
Event|Activity|SIMPLE_SEGMENT|15103,15108|false|false|false|C1283174||check
Finding|Functional Concept|SIMPLE_SEGMENT|15103,15108|false|false|false|C4321547|Check|check
Drug|Inorganic Chemical|SIMPLE_SEGMENT|15109,15121|false|false|false|C0013832;C3536863|Electrolyte [EPC];Electrolytes|electrolytes
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15109,15121|false|false|false|C0013832;C3536863|Electrolyte [EPC];Electrolytes|electrolytes
Event|Event|SIMPLE_SEGMENT|15109,15121|false|false|false|||electrolytes
Drug|Organic Chemical|SIMPLE_SEGMENT|15127,15136|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15127,15136|false|false|false|C0001927|albuterol|Albuterol
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|15144,15147|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|15144,15147|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|15144,15147|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Finding|Cell Function|SIMPLE_SEGMENT|15144,15147|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|SIMPLE_SEGMENT|15144,15147|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|15155,15158|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|SIMPLE_SEGMENT|15155,15158|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|15155,15158|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|SIMPLE_SEGMENT|15155,15158|false|false|false|||NEB
Finding|Cell Function|SIMPLE_SEGMENT|15155,15158|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|SIMPLE_SEGMENT|15155,15158|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|SIMPLE_SEGMENT|15166,15169|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|15170,15176|false|false|false|||wheeze
Finding|Sign or Symptom|SIMPLE_SEGMENT|15170,15176|false|false|false|C0043144|Wheezing|wheeze
Drug|Organic Chemical|SIMPLE_SEGMENT|15182,15193|false|false|false|C0027235|ipratropium|Ipratropium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15182,15193|false|false|false|C0027235|ipratropium|Ipratropium
Event|Event|SIMPLE_SEGMENT|15182,15193|false|false|false|||Ipratropium
Drug|Organic Chemical|SIMPLE_SEGMENT|15182,15201|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15182,15201|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Inorganic Chemical|SIMPLE_SEGMENT|15194,15201|false|false|false|C0006222|Bromides|Bromide
Event|Event|SIMPLE_SEGMENT|15194,15201|false|false|false|||Bromide
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|15194,15201|false|false|false|C0202341|Bromides measurement|Bromide
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|15202,15205|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|15202,15205|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|15202,15205|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Event|Event|SIMPLE_SEGMENT|15202,15205|false|false|false|||Neb
Finding|Cell Function|SIMPLE_SEGMENT|15202,15205|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|SIMPLE_SEGMENT|15202,15205|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|15208,15211|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|SIMPLE_SEGMENT|15208,15211|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|15208,15211|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|SIMPLE_SEGMENT|15208,15211|false|false|false|||NEB
Finding|Cell Function|SIMPLE_SEGMENT|15208,15211|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|SIMPLE_SEGMENT|15208,15211|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|SIMPLE_SEGMENT|15219,15222|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|15223,15229|false|false|false|||wheeze
Finding|Sign or Symptom|SIMPLE_SEGMENT|15223,15229|false|false|false|C0043144|Wheezing|wheeze
Event|Event|SIMPLE_SEGMENT|15234,15243|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|15234,15243|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|15234,15243|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|15234,15243|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|15234,15243|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15234,15255|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|15234,15255|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15244,15255|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|15244,15255|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|15244,15255|false|false|false|C0184758|Patient disposition|Disposition
Finding|Finding|SIMPLE_SEGMENT|15257,15265|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|15257,15265|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Procedure|Health Care Activity|SIMPLE_SEGMENT|15257,15270|false|false|false|C0023977|long-term care|Extended Care
Event|Activity|SIMPLE_SEGMENT|15266,15270|false|false|false|C1947933|care activity|Care
Event|Event|SIMPLE_SEGMENT|15266,15270|false|false|false|||Care
Finding|Finding|SIMPLE_SEGMENT|15266,15270|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|SIMPLE_SEGMENT|15266,15270|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Event|Event|SIMPLE_SEGMENT|15273,15281|false|false|false|||Facility
Finding|Intellectual Product|SIMPLE_SEGMENT|15273,15281|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|SIMPLE_SEGMENT|15289,15298|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|15289,15298|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|15289,15298|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|15289,15298|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|15289,15298|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|15289,15308|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15299,15308|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|15299,15308|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|15299,15308|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|15299,15308|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|15299,15308|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Intellectual Product|SIMPLE_SEGMENT|15310,15315|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|ACUTE
Event|Event|SIMPLE_SEGMENT|15316,15322|false|false|false|||ISSUES
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15339,15350|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|SIMPLE_SEGMENT|15339,15350|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|SIMPLE_SEGMENT|15339,15350|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|SIMPLE_SEGMENT|15339,15350|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15339,15358|false|false|false|C1145670|Respiratory Failure|respiratory failure
Event|Event|SIMPLE_SEGMENT|15351,15358|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|15351,15358|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|15351,15358|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|15351,15358|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15362,15368|false|false|false|C0036690;C0243026|Sepsis;Septicemia|Sepsis
Event|Event|SIMPLE_SEGMENT|15362,15368|false|false|false|||Sepsis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|15376,15383|false|false|false|C0042027|Urinary tract|urinary
Event|Event|SIMPLE_SEGMENT|15384,15390|false|false|false|||source
Finding|Finding|SIMPLE_SEGMENT|15384,15390|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Functional Concept|SIMPLE_SEGMENT|15384,15390|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Intellectual Product|SIMPLE_SEGMENT|15384,15390|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15417,15424|false|false|false|C0009319|Colitis|colitis
Event|Event|SIMPLE_SEGMENT|15417,15424|false|false|false|||colitis
Event|Event|SIMPLE_SEGMENT|15426,15433|false|false|false|||CHRONIC
Finding|Intellectual Product|SIMPLE_SEGMENT|15426,15433|false|false|false|C1547296|Chronic - Admission Level of Care Code|CHRONIC
Procedure|Health Care Activity|SIMPLE_SEGMENT|15426,15433|false|false|false|C1555457|Provision of recurring care for chronic illness|CHRONIC
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15446,15460|false|false|false|C0020676|Hypothyroidism|Hypothyroidism
Event|Event|SIMPLE_SEGMENT|15446,15460|false|false|false|||Hypothyroidism
Finding|Intellectual Product|SIMPLE_SEGMENT|15464,15471|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|15464,15471|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15464,15478|false|false|false|C0581384|Chronic anemia|Chronic anemia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15472,15478|false|false|false|C0002871|Anemia|anemia
Event|Event|SIMPLE_SEGMENT|15472,15478|false|false|false|||anemia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15482,15502|false|false|false|C0026266|Mitral Valve Insufficiency|Mitral regurgitation
Event|Event|SIMPLE_SEGMENT|15489,15502|false|false|false|||regurgitation
Finding|Finding|SIMPLE_SEGMENT|15489,15502|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|SIMPLE_SEGMENT|15489,15502|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|15489,15502|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15506,15518|false|false|false|C0029456|Osteoporosis|Osteoporosis
Event|Event|SIMPLE_SEGMENT|15506,15518|false|false|false|||Osteoporosis
Finding|Finding|SIMPLE_SEGMENT|15506,15518|false|false|false|C2911643|Encounter due to family history of osteoporosis|Osteoporosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15522,15538|false|false|false|C1527336|Sjogren's Syndrome|Sjogren syndrome
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15530,15538|false|false|false|C0039082|Syndrome|syndrome
Event|Event|SIMPLE_SEGMENT|15530,15538|false|false|false|||syndrome
Event|Event|SIMPLE_SEGMENT|15542,15551|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|15542,15551|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|15542,15551|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|15542,15551|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|15542,15551|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15552,15561|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15552,15561|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|15552,15561|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|15552,15561|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|15563,15569|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15563,15576|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|15563,15576|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15570,15576|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|15570,15576|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|15578,15583|false|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|15578,15583|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|15588,15596|false|false|false|||coherent
Finding|Finding|SIMPLE_SEGMENT|15588,15596|false|false|false|C4068804|Coherent|coherent
Event|Event|SIMPLE_SEGMENT|15598,15603|false|false|false|||Level
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15598,15620|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|15598,15620|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|SIMPLE_SEGMENT|15607,15620|false|false|false|||Consciousness
Finding|Finding|SIMPLE_SEGMENT|15607,15620|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|15607,15620|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15622,15627|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|15622,15627|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|15622,15627|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|15622,15627|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|15622,15627|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|15622,15627|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|15622,15627|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|15632,15643|false|false|false|||interactive
Finding|Functional Concept|SIMPLE_SEGMENT|15632,15643|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|15645,15653|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|15645,15653|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|15645,15653|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15654,15660|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|15654,15660|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|15654,15660|false|false|false|C1546481|What subject filter - Status|Status
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15669,15672|false|false|false|C3159311|BORNHOLM EYE DISEASE|Bed
Event|Event|SIMPLE_SEGMENT|15669,15672|false|false|false|||Bed
Finding|Intellectual Product|SIMPLE_SEGMENT|15669,15672|false|false|false|C2346952|Bachelor of Education|Bed
Event|Event|SIMPLE_SEGMENT|15678,15688|false|false|false|||assistance
Finding|Social Behavior|SIMPLE_SEGMENT|15678,15688|false|false|false|C0018896|Helping Behavior|assistance
Event|Event|SIMPLE_SEGMENT|15702,15712|false|false|false|||wheelchair
Finding|Finding|SIMPLE_SEGMENT|15702,15712|false|false|false|C2135586;C4321408|Wheelchair Usually Used;has wheelchair at home (history)|wheelchair
Event|Event|SIMPLE_SEGMENT|15717,15726|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|15717,15726|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|15717,15726|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|15717,15726|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|15717,15726|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15717,15739|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|15717,15739|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|15717,15739|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15727,15739|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|15727,15739|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|15727,15739|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Finding|Gene or Genome|SIMPLE_SEGMENT|15741,15745|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|SIMPLE_SEGMENT|15766,15774|false|false|false|||pleasure
Finding|Intellectual Product|SIMPLE_SEGMENT|15766,15774|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|SIMPLE_SEGMENT|15766,15774|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|SIMPLE_SEGMENT|15798,15802|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|15798,15802|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|15798,15802|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|15798,15802|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Event|Event|SIMPLE_SEGMENT|15825,15833|false|false|false|||admitted
Finding|Idea or Concept|SIMPLE_SEGMENT|15841,15849|false|false|false|C1547192|Organization unit type - Hospital|hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|15856,15867|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|SIMPLE_SEGMENT|15856,15867|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|SIMPLE_SEGMENT|15856,15867|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|SIMPLE_SEGMENT|15856,15867|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15856,15875|false|false|false|C1145670|Respiratory Failure|respiratory failure
Event|Event|SIMPLE_SEGMENT|15868,15875|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|15868,15875|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|15868,15875|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|15868,15875|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|SIMPLE_SEGMENT|15886,15896|false|false|false|||intubation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|15886,15896|false|false|false|C0021925|Intubation (procedure)|intubation
Event|Event|SIMPLE_SEGMENT|15901,15911|false|false|false|||mechanical
Finding|Functional Concept|SIMPLE_SEGMENT|15901,15911|false|false|false|C0443254|mechanical method|mechanical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|15901,15911|false|false|false|C0699886|Mechanical Treatments|mechanical
Event|Event|SIMPLE_SEGMENT|15913,15924|false|false|false|||ventilation
Finding|Physiologic Function|SIMPLE_SEGMENT|15913,15924|false|false|false|C0035203;C2945579|Respiration;Ventilation, function (observable entity)|ventilation
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|15913,15924|false|false|false|C0042491|Environmental air flow|ventilation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|15913,15924|false|false|false|C0554804|Assisted breathing|ventilation
Finding|Finding|SIMPLE_SEGMENT|15935,15941|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|15935,15941|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|SIMPLE_SEGMENT|15951,15962|false|false|false|||combination
Finding|Finding|SIMPLE_SEGMENT|15951,15962|false|false|false|C3811910|combination - answer to question|combination
Event|Event|SIMPLE_SEGMENT|15966,15972|false|false|false|||severe
Finding|Finding|SIMPLE_SEGMENT|15966,15972|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|15966,15972|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Event|Event|SIMPLE_SEGMENT|15974,15982|false|false|false|||weakness
Finding|Sign or Symptom|SIMPLE_SEGMENT|15974,15982|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Finding|Intellectual Product|SIMPLE_SEGMENT|15993,16000|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|15993,16000|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|15993,16008|false|false|false|C0008679|Chronic disease|chronic illness
Finding|Finding|SIMPLE_SEGMENT|15993,16008|false|false|false|C2186378|Reported history of chronic illness|chronic illness
Event|Event|SIMPLE_SEGMENT|16001,16008|false|false|false|||illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|16001,16008|false|false|false|C0221423|Illness (finding)|illness
Anatomy|Tissue|SIMPLE_SEGMENT|16010,16017|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|16010,16017|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Pathologic Function|SIMPLE_SEGMENT|16010,16027|false|false|false|C0032227|Pleural effusion (disorder)|pleural effusions
Event|Event|SIMPLE_SEGMENT|16018,16027|false|false|false|||effusions
Finding|Pathologic Function|SIMPLE_SEGMENT|16018,16027|false|false|false|C0013687|effusion|effusions
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|16033,16042|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|16033,16042|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|16033,16042|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|16033,16048|false|false|false|C0034063|Pulmonary Edema|pulmonary edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|16043,16048|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|16043,16048|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|16043,16048|false|false|false|C0013604|Edema|edema
Drug|Substance|SIMPLE_SEGMENT|16050,16055|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|16050,16055|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|16050,16055|false|false|false|C1546638|Fluid Specimen Code|fluid
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|16064,16069|false|false|false|C0024109|Lung|lungs
Event|Event|SIMPLE_SEGMENT|16086,16091|false|false|false|||found
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|16103,16110|false|false|false|C0042027|Urinary tract|urinary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|16103,16116|false|false|false|C0042027;C1508753|Urinary system;Urinary tract|urinary tract
Anatomy|Body System|SIMPLE_SEGMENT|16103,16116|false|false|false|C0042027;C1508753|Urinary system;Urinary tract|urinary tract
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|16103,16126|false|false|false|C0042029|Urinary tract infection|urinary tract infection
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|16111,16116|false|false|false|C1185740|Tract|tract
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|16117,16126|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|16117,16126|false|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|16117,16126|false|false|false|C3714514|Infection|infection
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|16135,16141|false|false|false|C0036690;C0243026|Sepsis;Septicemia|sepsis
Event|Event|SIMPLE_SEGMENT|16135,16141|false|false|false|||sepsis
Event|Event|SIMPLE_SEGMENT|16143,16154|false|false|false|||bloodstream
Finding|Physiologic Function|SIMPLE_SEGMENT|16143,16154|false|false|false|C0005775|Blood Circulation|bloodstream
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|16156,16165|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|16156,16165|false|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|16156,16165|false|false|false|C3714514|Infection|infection
Finding|Finding|SIMPLE_SEGMENT|16174,16180|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|16174,16180|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|SIMPLE_SEGMENT|16186,16197|false|false|false|||contributed
Attribute|Clinical Attribute|SIMPLE_SEGMENT|16206,16217|false|false|false|C0231832|Respiratory rate|respiratory
Event|Event|SIMPLE_SEGMENT|16206,16217|false|false|false|||respiratory
Finding|Body Substance|SIMPLE_SEGMENT|16206,16217|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|SIMPLE_SEGMENT|16206,16217|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|SIMPLE_SEGMENT|16206,16217|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Event|Event|SIMPLE_SEGMENT|16219,16226|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|16219,16226|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|16219,16226|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|16219,16226|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|SIMPLE_SEGMENT|16237,16244|false|false|false|||treated
Drug|Antibiotic|SIMPLE_SEGMENT|16250,16261|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|SIMPLE_SEGMENT|16250,16261|false|false|false|||antibiotics
Event|Event|SIMPLE_SEGMENT|16268,16276|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|16268,16276|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|16268,16276|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|SIMPLE_SEGMENT|16282,16291|false|false|false|||breathing
Event|Event|SIMPLE_SEGMENT|16292,16300|false|false|false|||improved
Event|Event|SIMPLE_SEGMENT|16328,16337|false|false|false|||extubated
Event|Event|SIMPLE_SEGMENT|16359,16369|false|false|false|||discharged
Event|Event|SIMPLE_SEGMENT|16373,16378|false|false|false|||rehab
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|16373,16378|false|false|false|C0034991|Rehabilitation therapy|rehab
Event|Event|SIMPLE_SEGMENT|16402,16411|false|false|false|||intensive
Finding|Finding|SIMPLE_SEGMENT|16413,16421|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Finding|Functional Concept|SIMPLE_SEGMENT|16413,16421|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|16413,16421|false|false|false|C0031809|Physical Examination|physical
Finding|Intellectual Product|SIMPLE_SEGMENT|16413,16429|false|false|false|C1547999|Diagnostic Service Section ID - Physical Therapy|physical therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|16413,16429|false|false|false|C0949766|Physical therapy|physical therapy
Event|Event|SIMPLE_SEGMENT|16422,16429|false|false|false|||therapy
Finding|Finding|SIMPLE_SEGMENT|16422,16429|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|SIMPLE_SEGMENT|16422,16429|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|16422,16429|false|false|false|C0087111|Therapeutic procedure|therapy
Event|Event|SIMPLE_SEGMENT|16439,16448|false|false|false|||nutrition
Finding|Finding|SIMPLE_SEGMENT|16439,16448|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|nutrition
Finding|Intellectual Product|SIMPLE_SEGMENT|16439,16448|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|nutrition
Finding|Organism Function|SIMPLE_SEGMENT|16439,16448|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|nutrition
Procedure|Research Activity|SIMPLE_SEGMENT|16439,16448|false|false|false|C0600072;C1521729|Feeding and dietary regimes;Nutritional Study|nutrition
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|16439,16448|false|false|false|C0600072;C1521729|Feeding and dietary regimes;Nutritional Study|nutrition
Event|Event|SIMPLE_SEGMENT|16457,16466|false|false|false|||optimized
Event|Event|SIMPLE_SEGMENT|16470,16474|false|false|false|||help
Finding|Intellectual Product|SIMPLE_SEGMENT|16470,16474|false|false|false|C1552861|Help document|help
Event|Event|SIMPLE_SEGMENT|16480,16488|false|false|false|||continue
Event|Event|SIMPLE_SEGMENT|16499,16507|false|false|false|||strength
Finding|Idea or Concept|SIMPLE_SEGMENT|16499,16507|false|false|false|C0808080|Strength (attribute)|strength
Event|Event|SIMPLE_SEGMENT|16525,16535|false|false|false|||discharged
Event|Event|SIMPLE_SEGMENT|16541,16546|false|false|false|||rehab
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|16541,16546|false|false|false|C0034991|Rehabilitation therapy|rehab
Event|Event|SIMPLE_SEGMENT|16557,16561|false|false|false|||need
Event|Event|SIMPLE_SEGMENT|16565,16571|false|false|false|||follow
Finding|Intellectual Product|SIMPLE_SEGMENT|16586,16598|false|false|false|C1547426|Location Service Code - Primary Care|primary care
Procedure|Health Care Activity|SIMPLE_SEGMENT|16586,16598|false|false|false|C0033137|Primary Health Care|primary care
Event|Activity|SIMPLE_SEGMENT|16594,16598|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|16594,16598|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|16594,16598|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|16594,16598|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|16599,16605|false|false|false|C2348314|Doctor - Title|doctor
Event|Event|SIMPLE_SEGMENT|16617,16621|false|false|false|||made
Event|Event|SIMPLE_SEGMENT|16636,16643|false|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|16636,16643|false|false|false|C0392747|Changing|changes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|16652,16663|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16652,16663|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|16652,16663|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|16652,16663|false|false|false|C4284232|Medications|medications
Drug|Organic Chemical|SIMPLE_SEGMENT|16677,16687|false|false|false|C0015620|famotidine|famotidine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16677,16687|false|false|false|C0015620|famotidine|famotidine
Event|Event|SIMPLE_SEGMENT|16677,16687|false|false|false|||famotidine
Finding|Functional Concept|SIMPLE_SEGMENT|16693,16701|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|16696,16701|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|16696,16701|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|16718,16727|false|false|false|C0017168|Gastroesophageal reflux disease|heartburn
Event|Event|SIMPLE_SEGMENT|16718,16727|false|false|false|||heartburn
Finding|Sign or Symptom|SIMPLE_SEGMENT|16718,16727|false|false|false|C0018834|Heartburn|heartburn
Event|Event|SIMPLE_SEGMENT|16731,16738|false|false|false|||STARTED
Drug|Organic Chemical|SIMPLE_SEGMENT|16739,16752|false|false|false|C0040864|triamcinolone|triamcinolone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16739,16752|false|false|false|C0040864|triamcinolone|triamcinolone
Drug|Organic Chemical|SIMPLE_SEGMENT|16739,16762|false|false|false|C0040866|triamcinolone acetonide|triamcinolone acetonide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16739,16762|false|false|false|C0040866|triamcinolone acetonide|triamcinolone acetonide
Event|Event|SIMPLE_SEGMENT|16753,16762|false|false|false|||acetonide
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|16770,16775|false|false|false|C0700385;C0705539;C1378128|Cream;Dairy Cream;Emollient Cream|cream
Drug|Food|SIMPLE_SEGMENT|16770,16775|false|false|false|C0700385;C0705539;C1378128|Cream;Dairy Cream;Emollient Cream|cream
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|16782,16787|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Event|Event|SIMPLE_SEGMENT|16782,16787|false|false|false|||times
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|16799,16803|false|false|false|C5779629|Eruption of skin (disorder)|rash
Event|Event|SIMPLE_SEGMENT|16799,16803|false|false|false|||rash
Finding|Pathologic Function|SIMPLE_SEGMENT|16799,16803|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|SIMPLE_SEGMENT|16799,16803|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|16817,16827|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16817,16827|false|false|false|C0065374|lisinopril|lisinopril
Event|Event|SIMPLE_SEGMENT|16817,16827|false|false|false|||lisinopril
Finding|Functional Concept|SIMPLE_SEGMENT|16832,16840|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|16835,16840|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|16835,16840|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Finding|SIMPLE_SEGMENT|16851,16855|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|SIMPLE_SEGMENT|16851,16855|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|SIMPLE_SEGMENT|16851,16855|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|16856,16861|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|16856,16861|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|16856,16861|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Event|SIMPLE_SEGMENT|16863,16871|false|false|false|||pressure
Finding|Finding|SIMPLE_SEGMENT|16863,16871|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|16863,16871|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|16863,16871|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|16863,16871|false|false|false|C0033095||pressure
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|16876,16881|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|16876,16881|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|16876,16881|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|16876,16889|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Event|Event|SIMPLE_SEGMENT|16882,16889|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|16882,16889|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|16882,16889|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|16882,16889|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Drug|Organic Chemical|SIMPLE_SEGMENT|16901,16909|false|false|false|C1692318|docusate|docusate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16901,16909|false|false|false|C1692318|docusate|docusate
Event|Event|SIMPLE_SEGMENT|16901,16909|false|false|false|||docusate
Drug|Organic Chemical|SIMPLE_SEGMENT|16911,16917|false|false|false|C0282139|Colace|Colace
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|16911,16917|false|false|false|C0282139|Colace|Colace
Finding|Functional Concept|SIMPLE_SEGMENT|16925,16933|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|16928,16933|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|16928,16933|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Event|SIMPLE_SEGMENT|16951,16963|false|false|false|||constipation
Finding|Sign or Symptom|SIMPLE_SEGMENT|16951,16963|false|false|false|C0009806|Constipation|constipation
Finding|Idea or Concept|SIMPLE_SEGMENT|16967,16976|false|false|false|C0549178|Continuous|CONTINUED
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|16977,16987|false|false|false|C0042313|vancomycin|vancomycin
Drug|Antibiotic|SIMPLE_SEGMENT|16977,16987|false|false|false|C0042313|vancomycin|vancomycin
Event|Event|SIMPLE_SEGMENT|16977,16987|false|false|false|||vancomycin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|16977,16987|false|false|false|C0489941|Vancomycin measurement|vancomycin
Drug|Clinical Drug|SIMPLE_SEGMENT|16977,16992|false|false|false|C0360373||vancomycin oral
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|16988,16992|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|16988,16992|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|16988,16992|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|16988,16992|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|16988,16999|false|false|false|C1273619|Oral Liquid Product|oral liquid
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|16993,16999|false|false|false|C0302908;C1697794|Liquid Dosage Form;Liquid substance|liquid
Drug|Substance|SIMPLE_SEGMENT|16993,16999|false|false|false|C0302908;C1697794|Liquid Dosage Form;Liquid substance|liquid
Event|Event|SIMPLE_SEGMENT|16993,16999|false|false|false|||liquid
Finding|Finding|SIMPLE_SEGMENT|16993,16999|false|false|false|C1304698|Liquid (finding)|liquid
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|16993,16999|false|false|false|C0301571|Liquid diet|liquid
Finding|Functional Concept|SIMPLE_SEGMENT|17004,17012|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|17007,17012|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|17007,17012|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Event|SIMPLE_SEGMENT|17034,17037|false|false|false|||day
Finding|Idea or Concept|SIMPLE_SEGMENT|17034,17037|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|17034,17037|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Food|SIMPLE_SEGMENT|17048,17053|false|false|false|C0452588|Start brand of breakfast cereal|START
Event|Event|SIMPLE_SEGMENT|17048,17053|false|false|false|||START
Finding|Intellectual Product|SIMPLE_SEGMENT|17048,17053|false|false|false|C1552850|start - HtmlLinkType|START
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|17048,17053|false|false|false|C5447432|Collagen Tile Brachytherapy|START
Finding|Gene or Genome|SIMPLE_SEGMENT|17074,17077|false|false|false|C1422467|CIAO3 gene|prn
Finding|Intellectual Product|SIMPLE_SEGMENT|17078,17084|false|false|false|C1705102|Volume (publication)|volume
Finding|Pathologic Function|SIMPLE_SEGMENT|17078,17093|false|false|false|C0546817|Hypervolemia (finding)|volume overload
Event|Event|SIMPLE_SEGMENT|17085,17093|false|false|false|||overload
Procedure|Health Care Activity|SIMPLE_SEGMENT|17096,17104|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|17105,17117|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|17105,17117|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|17105,17117|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

