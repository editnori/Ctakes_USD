 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|39,48|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|39,48|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|39,53|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|73,82|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|73,82|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|73,82|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|73,82|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|73,82|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|73,87|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|105,110|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|105,110|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|105,110|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|129,132|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|140,147|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|140,147|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|149,157|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|Allergies|181,190|false|false|false|C1717415||Allergies
Event|Event|Allergies|181,190|false|false|false|||Allergies
Finding|Pathologic Function|Allergies|181,190|false|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|Allergies|193,215|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|Allergies|201,205|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|Allergies|201,205|false|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|Allergies|201,215|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Event|Event|Allergies|206,215|false|false|false|||Reactions
Event|Event|Allergies|218,227|false|false|false|||Attending
Finding|Functional Concept|Allergies|218,227|false|false|false|C1999232|Attending (action)|Attending
Event|Event|Chief Complaint|253,260|false|false|false|||fatigue
Finding|Sign or Symptom|Chief Complaint|253,260|false|false|false|C0015672|Fatigue|fatigue
Disorder|Disease or Syndrome|Chief Complaint|262,268|false|false|false|C0002871|Anemia|anemia
Event|Event|Chief Complaint|262,268|false|false|false|||anemia
Finding|Classification|Chief Complaint|271,276|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|277,285|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|277,285|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|289,307|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|298,307|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|298,307|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|298,307|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|298,307|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|298,307|false|false|false|C0184661|Interventional procedure|Procedure
Finding|Idea or Concept|History of Present Illness|362,366|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|History of Present Illness|362,366|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|History of Present Illness|367,370|false|false|false|||old
Event|Event|History of Present Illness|389,396|false|false|false|||medical
Finding|Functional Concept|History of Present Illness|389,396|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|History of Present Illness|389,396|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|History of Present Illness|389,396|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|History of Present Illness|389,396|false|false|false|C0199168|Medical service|medical
Event|Event|History of Present Illness|398,405|false|false|false|||history
Finding|Conceptual Entity|History of Present Illness|398,405|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|398,405|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|398,405|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|398,408|false|false|false|C0262926|Medical History|history of
Finding|Gene or Genome|History of Present Illness|409,413|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Intellectual Product|History of Present Illness|409,413|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Disorder|Disease or Syndrome|History of Present Illness|420,432|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|History of Present Illness|420,432|false|false|false|||hypertension
Attribute|Clinical Attribute|History of Present Illness|434,439|false|false|false|C1300072|Tumor stage|stage
Finding|Intellectual Product|History of Present Illness|434,442|false|false|false|C0441772|Stage level 4|stage IV
Disorder|Disease or Syndrome|History of Present Illness|443,446|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Event|Event|History of Present Illness|443,446|false|false|false|||CKD
Disorder|Disease or Syndrome|History of Present Illness|448,451|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|448,451|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|History of Present Illness|448,451|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|History of Present Illness|448,451|false|false|false|||CAD
Finding|Gene or Genome|History of Present Illness|448,451|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|History of Present Illness|448,451|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|History of Present Illness|448,451|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|448,451|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Finding|Pathologic Function|History of Present Illness|457,464|false|false|false|C5441917|Distant Metastasis|distant
Drug|Inorganic Chemical|History of Present Illness|477,482|false|false|false|C0025552|Metals|metal
Event|Event|History of Present Illness|483,488|false|false|false|||stent
Disorder|Disease or Syndrome|History of Present Illness|490,496|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|History of Present Illness|490,496|false|false|false|||stroke
Finding|Finding|History of Present Illness|490,496|false|false|false|C5977286|Stroke (heart beat)|stroke
Disorder|Disease or Syndrome|History of Present Illness|516,520|false|false|false|C0151950|Deep thrombophlebitis|DVTs
Event|Event|History of Present Illness|516,520|false|false|false|||DVTs
Drug|Organic Chemical|History of Present Illness|525,533|false|false|false|C0699129|Coumadin|Coumadin
Drug|Pharmacologic Substance|History of Present Illness|525,533|false|false|false|C0699129|Coumadin|Coumadin
Procedure|Diagnostic Procedure|History of Present Illness|546,554|false|false|false|C0203057|Upper gastrointestinal tract series|upper GI
Finding|Pathologic Function|History of Present Illness|546,563|false|false|false|C0041909|Upper gastrointestinal hemorrhage|upper GI bleeding
Finding|Pathologic Function|History of Present Illness|552,563|false|false|false|C0017181|Gastrointestinal Hemorrhage|GI bleeding
Event|Event|History of Present Illness|555,563|false|false|false|||bleeding
Finding|Pathologic Function|History of Present Illness|555,563|false|false|false|C0019080|Hemorrhage|bleeding
Event|Event|History of Present Illness|573,577|false|false|false|||sent
Attribute|Clinical Attribute|History of Present Illness|593,602|false|false|false|C0804815||physician
Disorder|Disease or Syndrome|History of Present Illness|607,613|false|false|false|C0002871|Anemia|anemia
Event|Event|History of Present Illness|607,613|false|false|false|||anemia
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|615,618|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|History of Present Illness|615,618|false|false|false|C0019046|Hemoglobin|Hgb
Event|Event|History of Present Illness|615,618|false|false|false|||Hgb
Finding|Gene or Genome|History of Present Illness|615,618|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|History of Present Illness|615,618|false|false|false|C0019029|Hemoglobin concentration|Hgb
Finding|Body Substance|History of Present Illness|630,637|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|630,637|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|630,637|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|642,650|false|false|false|||admitted
Anatomy|Body Location or Region|History of Present Illness|692,697|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|History of Present Illness|692,697|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|692,707|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|698,707|false|false|false|C0015385|Limb structure|extremity
Disorder|Disease or Syndrome|History of Present Illness|708,712|false|false|false|C0151950|Deep thrombophlebitis|DVTs
Event|Event|History of Present Illness|708,712|false|false|false|||DVTs
Event|Event|History of Present Illness|722,729|false|false|false|||started
Drug|Biologically Active Substance|History of Present Illness|733,740|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|History of Present Illness|733,740|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|History of Present Illness|733,740|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Event|Event|History of Present Illness|733,740|false|false|false|||heparin
Event|Event|History of Present Illness|748,757|false|false|false|||inpatient
Finding|Idea or Concept|History of Present Illness|748,757|false|true|false|C1548438;C1549404|Patient Class - Inpatient;Referral category - Inpatient|inpatient
Procedure|Health Care Activity|History of Present Illness|748,757|false|true|false|C1555324|inpatient encounter|inpatient
Event|Event|History of Present Illness|763,778|false|false|false|||anticoagulation
Finding|Finding|History of Present Illness|763,778|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|History of Present Illness|763,778|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|763,778|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Event|Event|History of Present Illness|783,794|false|false|false|||complicated
Finding|Finding|History of Present Illness|798,806|false|false|false|C0205082|Severe (severity modifier)|severely
Finding|Finding|History of Present Illness|808,820|false|false|false|C0240671|Partial thromboplastin time increased (finding)|elevated PTT
Disorder|Neoplastic Process|History of Present Illness|817,820|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|History of Present Illness|817,820|false|false|false|||PTT
Procedure|Laboratory Procedure|History of Present Illness|817,820|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Procedure|Diagnostic Procedure|History of Present Illness|832,840|false|false|false|C0203057|Upper gastrointestinal tract series|upper GI
Finding|Pathologic Function|History of Present Illness|832,846|false|false|false|C0041909|Upper gastrointestinal hemorrhage|upper GI bleed
Finding|Pathologic Function|History of Present Illness|838,846|false|false|false|C0017181|Gastrointestinal Hemorrhage|GI bleed
Event|Event|History of Present Illness|841,846|false|false|false|||bleed
Finding|Pathologic Function|History of Present Illness|841,846|false|false|false|C0019080|Hemorrhage|bleed
Event|Event|History of Present Illness|848,857|false|false|false|||Endoscopy
Procedure|Diagnostic Procedure|History of Present Illness|848,857|false|false|false|C0014245;C0079278|Endoscopy (procedure);Endoscopy, Gastrointestinal|Endoscopy
Event|Event|History of Present Illness|862,869|false|false|false|||notable
Finding|Idea or Concept|History of Present Illness|875,886|false|false|false|C0750502|Significant|significant
Disorder|Disease or Syndrome|History of Present Illness|887,895|false|false|false|C0041834|Erythema|erythema
Event|Event|History of Present Illness|887,895|false|false|false|||erythema
Disorder|Disease or Syndrome|History of Present Illness|897,919|false|false|false|C0333307|Superficial ulcer|superficial ulceration
Event|Event|History of Present Illness|909,919|false|false|false|||ulceration
Finding|Pathologic Function|History of Present Illness|909,919|false|false|false|C0041582;C3887532|Ulcer;Ulceration|ulceration
Disorder|Disease or Syndrome|History of Present Illness|925,934|false|false|false|C0017152|Gastritis|gastritis
Event|Event|History of Present Illness|925,934|false|false|false|||gastritis
Event|Event|History of Present Illness|951,959|false|false|false|||bleeding
Finding|Pathologic Function|History of Present Illness|951,959|true|false|false|C0019080|Hemorrhage|bleeding
Event|Event|History of Present Illness|969,975|false|false|false|||placed
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|979,982|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|979,982|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|History of Present Illness|979,982|false|false|false|C1530795|BID protein, human|BID
Event|Event|History of Present Illness|979,982|false|false|false|||BID
Finding|Gene or Genome|History of Present Illness|979,982|false|false|false|C1332410|BID gene|BID
Drug|Pharmacologic Substance|History of Present Illness|983,986|false|false|false|C0358591|Proton Pump Inhibitors|PPI
Event|Event|History of Present Illness|983,986|false|false|false|||PPI
Finding|Physiologic Function|History of Present Illness|983,986|false|false|false|C0871125|Prepulse Inhibition|PPI
Event|Event|History of Present Illness|987,998|false|false|false|||prophylaxis
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|987,998|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Event|Event|History of Present Illness|1020,1027|false|false|false|||bridged
Drug|Organic Chemical|History of Present Illness|1031,1039|false|false|false|C0699129|Coumadin|Coumadin
Drug|Pharmacologic Substance|History of Present Illness|1031,1039|false|false|false|C0699129|Coumadin|Coumadin
Event|Event|History of Present Illness|1031,1039|false|false|false|||Coumadin
Event|Event|History of Present Illness|1046,1053|false|false|false|||planned
Event|Event|History of Present Illness|1056,1061|false|false|false|||month
Finding|Idea or Concept|History of Present Illness|1056,1061|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|History of Present Illness|1056,1061|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Event|Event|History of Present Illness|1063,1069|false|false|false|||course
Attribute|Clinical Attribute|History of Present Illness|1075,1078|false|false|false|C0368980|Coagulation tissue factor induced.INR|INR
Event|Event|History of Present Illness|1075,1078|false|false|false|||INR
Procedure|Laboratory Procedure|History of Present Illness|1075,1078|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1075,1078|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Event|Event|History of Present Illness|1082,1089|false|false|false|||managed
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1097,1102|false|false|false|C0034991|Rehabilitation therapy|rehab
Event|Event|History of Present Illness|1103,1111|false|false|false|||facility
Finding|Intellectual Product|History of Present Illness|1103,1111|false|false|false|C4695111|ADMIN.FACILITY|facility
Event|Event|History of Present Illness|1125,1133|false|false|false|||followed
Event|Event|History of Present Illness|1193,1198|false|false|false|||noted
Event|Event|History of Present Illness|1210,1217|false|false|false|||fatigue
Finding|Sign or Symptom|History of Present Illness|1210,1217|false|false|false|C0015672|Fatigue|fatigue
Event|Event|History of Present Illness|1230,1239|false|false|false|||shortness
Attribute|Clinical Attribute|History of Present Illness|1230,1249|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|History of Present Illness|1230,1249|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|History of Present Illness|1243,1249|false|false|false|C0225386|Breath|breath
Event|Event|History of Present Illness|1251,1261|false|false|false|||exertional
Finding|Sign or Symptom|History of Present Illness|1251,1261|false|false|false|C0239313|exercise induced|exertional
Anatomy|Body Location or Region|History of Present Illness|1274,1279|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|1274,1279|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|1274,1284|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|1274,1284|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|1280,1284|false|true|false|C2598155||pain
Event|Event|History of Present Illness|1280,1284|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|1280,1284|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1280,1284|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|1286,1294|false|false|false|||relieved
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1300,1304|false|false|false|C1742913|REST protein, human|rest
Drug|Biologically Active Substance|History of Present Illness|1300,1304|false|false|false|C1742913|REST protein, human|rest
Event|Event|History of Present Illness|1300,1304|false|false|false|||rest
Finding|Daily or Recreational Activity|History of Present Illness|1300,1304|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Gene or Genome|History of Present Illness|1300,1304|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Molecular Function|History of Present Illness|1300,1304|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Finding|History of Present Illness|1310,1321|false|false|false|C0332516|Symmetrical|symmetrical
Anatomy|Body Location or Region|History of Present Illness|1322,1327|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|History of Present Illness|1322,1327|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1322,1337|false|false|false|C0023216|Lower Extremity|lower extremity
Finding|Pathologic Function|History of Present Illness|1322,1346|false|false|false|C0581394|Swelling of lower limb|lower extremity swelling
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1328,1337|false|false|false|C0015385|Limb structure|extremity
Finding|Sign or Symptom|History of Present Illness|1328,1346|false|false|false|C0158369|Swelling of limb|extremity swelling
Event|Event|History of Present Illness|1338,1346|false|false|false|||swelling
Finding|Finding|History of Present Illness|1338,1346|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|History of Present Illness|1338,1346|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Event|Event|History of Present Illness|1361,1367|false|false|false|||period
Finding|Organism Function|History of Present Illness|1361,1367|false|false|false|C0025344|Menstruation|period
Procedure|Research Activity|History of Present Illness|1361,1367|false|false|false|C2347804|Clinical Trial Period|period
Event|Event|History of Present Illness|1372,1379|false|false|false|||reports
Event|Event|History of Present Illness|1389,1397|false|false|false|||appetite
Finding|Organism Function|History of Present Illness|1389,1397|false|false|false|C0003618|Desire for food|appetite
Event|Event|History of Present Illness|1398,1406|false|false|false|||remained
Event|Event|History of Present Illness|1407,1411|false|false|false|||good
Finding|Idea or Concept|History of Present Illness|1407,1411|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1421,1426|false|false|false|C0021853|Intestines|bowel
Finding|Organism Function|History of Present Illness|1421,1435|false|false|false|C0011135|Defecation|bowel function
Event|Event|History of Present Illness|1427,1435|false|false|false|||function
Finding|Finding|History of Present Illness|1427,1435|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|History of Present Illness|1427,1435|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|History of Present Illness|1427,1435|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|History of Present Illness|1427,1435|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Event|Event|History of Present Illness|1440,1446|false|false|false|||normal
Event|Event|History of Present Illness|1452,1458|false|false|false|||denies
Finding|Finding|History of Present Illness|1459,1465|false|false|false|C4554530|Bloody|bloody
Finding|Sign or Symptom|History of Present Illness|1459,1472|true|false|false|C1321898|Blood in stool|bloody stools
Attribute|Clinical Attribute|History of Present Illness|1466,1472|true|false|false|C0489144||stools
Event|Event|History of Present Illness|1466,1472|false|false|false|||stools
Finding|Body Substance|History of Present Illness|1466,1472|true|false|false|C0015733|Feces|stools
Finding|Sign or Symptom|History of Present Illness|1477,1487|false|false|false|C0474585||dark stool
Event|Event|History of Present Illness|1482,1487|false|false|false|||stool
Finding|Body Substance|History of Present Illness|1482,1487|false|false|false|C0015733|Feces|stool
Event|Event|History of Present Illness|1500,1509|false|false|false|||presented
Disorder|Disease or Syndrome|History of Present Illness|1517,1520|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|1517,1520|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|History of Present Illness|1517,1520|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1517,1520|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|History of Present Illness|1517,1520|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|History of Present Illness|1517,1520|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|History of Present Illness|1517,1520|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|History of Present Illness|1517,1520|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|History of Present Illness|1517,1520|false|false|false|||PCP
Finding|Gene or Genome|History of Present Illness|1517,1520|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|History of Present Illness|1517,1520|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|History of Present Illness|1521,1527|false|false|false|||office
Finding|Idea or Concept|History of Present Illness|1521,1527|false|false|false|C1549636|Address type - Office|office
Event|Event|History of Present Illness|1533,1538|false|false|false|||rehab
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1533,1538|false|false|false|C0034991|Rehabilitation therapy|rehab
Event|Event|History of Present Illness|1540,1549|false|false|false|||reporting
Event|Event|History of Present Illness|1561,1570|false|false|false|||shortness
Attribute|Clinical Attribute|History of Present Illness|1561,1580|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|History of Present Illness|1561,1580|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|History of Present Illness|1574,1580|false|false|false|C0225386|Breath|breath
Event|Event|History of Present Illness|1585,1592|false|false|false|||fatigue
Finding|Sign or Symptom|History of Present Illness|1585,1592|false|false|false|C0015672|Fatigue|fatigue
Event|Event|History of Present Illness|1603,1608|false|false|false|||found
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1619,1622|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|History of Present Illness|1619,1622|false|false|false|C0019046|Hemoglobin|Hgb
Event|Event|History of Present Illness|1619,1622|false|false|false|||Hgb
Finding|Gene or Genome|History of Present Illness|1619,1622|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|History of Present Illness|1619,1622|false|false|false|C0019029|Hemoglobin concentration|Hgb
Event|Event|History of Present Illness|1652,1655|false|false|false|||CXR
Procedure|Diagnostic Procedure|History of Present Illness|1652,1655|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|History of Present Illness|1666,1670|false|false|false|||sent
Event|Event|History of Present Illness|1682,1684|false|false|false|||ED
Finding|Idea or Concept|History of Present Illness|1702,1709|false|false|false|C1555582|Initial (abbreviation)|initial
Event|Event|History of Present Illness|1710,1716|false|false|false|||vitals
Event|Event|History of Present Illness|1730,1731|false|false|false|||P
Attribute|Clinical Attribute|History of Present Illness|1755,1759|false|false|false|C2317096|Saturation of Peripheral Oxygen|SPO2
Event|Event|History of Present Illness|1770,1774|false|false|false|||Exam
Finding|Functional Concept|History of Present Illness|1770,1774|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|History of Present Illness|1770,1774|false|false|false|C0582103|Medical Examination|Exam
Event|Event|History of Present Illness|1779,1786|false|false|false|||notable
Event|Event|History of Present Illness|1797,1805|false|false|false|||negative
Finding|Classification|History of Present Illness|1797,1805|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|History of Present Illness|1797,1805|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|History of Present Illness|1797,1805|false|false|false|C5237010|Expression Negative|negative
Event|Event|History of Present Illness|1806,1811|false|false|false|||stool
Finding|Body Substance|History of Present Illness|1806,1811|false|false|false|C0015733|Feces|stool
Event|Event|History of Present Illness|1814,1821|false|false|false|||Imaging
Finding|Finding|History of Present Illness|1814,1821|false|false|false|C0740845|Imaging problem|Imaging
Procedure|Diagnostic Procedure|History of Present Illness|1814,1821|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|Imaging
Event|Event|History of Present Illness|1826,1833|false|false|false|||notable
Attribute|Clinical Attribute|History of Present Illness|1857,1861|false|false|false|C4318566|Deep Resection Margin|deep
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1857,1866|false|false|false|C0226514|Structure of deep vein|deep vein
Disorder|Disease or Syndrome|History of Present Illness|1857,1877|false|false|false|C0149871;C0340708|Deep Vein Thrombosis;Deep vein thrombosis of lower limb|deep vein thrombosis
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1862,1866|false|false|false|C0042449|Veins|vein
Finding|Pathologic Function|History of Present Illness|1862,1877|false|false|false|C0042487|Venous Thrombosis|vein thrombosis
Event|Event|History of Present Illness|1867,1877|false|false|false|||thrombosis
Finding|Pathologic Function|History of Present Illness|1867,1877|false|false|false|C0040053|Thrombosis|thrombosis
Disorder|Disease or Syndrome|History of Present Illness|1900,1909|false|false|false|C0751438|Posterior pituitary disease|posterior
Event|Event|History of Present Illness|1900,1909|false|false|false|||posterior
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1900,1922|false|false|false|C0226832|Structure of posterior tibial vein|posterior tibial veins
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1910,1916|false|false|false|C0040184|Bone structure of tibia|tibial
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1910,1922|false|false|false|C0447138|Tibial vein structure|tibial veins
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1917,1922|false|false|false|C0042449|Veins|veins
Event|Event|History of Present Illness|1917,1922|false|false|false|||veins
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1917,1922|false|false|false|C0398102|Procedure on vein|veins
Event|Event|History of Present Illness|1950,1958|false|false|false|||thrombus
Finding|Pathologic Function|History of Present Illness|1950,1958|false|false|false|C0087086;C0302148|Blood Clot;Thrombus|thrombus
Event|Event|History of Present Illness|1976,1985|false|false|false|||decreased
Finding|Finding|History of Present Illness|1990,1993|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|History of Present Illness|1990,1993|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Attribute|Clinical Attribute|History of Present Illness|1994,1998|true|false|false|C4318566|Deep Resection Margin|deep
Disorder|Disease or Syndrome|History of Present Illness|1994,2016|true|false|false|C0149871|Deep Vein Thrombosis|deep venous thrombosis
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1999,2005|false|false|false|C0042449|Veins|venous
Finding|Finding|History of Present Illness|1999,2016|true|false|false|C0042487;C0517555|Venous Thrombosis;Venous thrombosis after immobility|venous thrombosis
Finding|Pathologic Function|History of Present Illness|1999,2016|true|false|false|C0042487;C0517555|Venous Thrombosis;Venous thrombosis after immobility|venous thrombosis
Event|Event|History of Present Illness|2006,2016|false|false|false|||thrombosis
Finding|Pathologic Function|History of Present Illness|2006,2016|true|false|false|C0040053|Thrombosis|thrombosis
Anatomy|Body Location or Region|History of Present Illness|2028,2033|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|History of Present Illness|2028,2033|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2028,2043|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2034,2043|false|false|false|C0015385|Limb structure|extremity
Event|Event|History of Present Illness|2050,2055|false|false|false|||Right
Finding|Functional Concept|History of Present Illness|2050,2055|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Drug|Chemical Viewed Structurally|History of Present Illness|2056,2063|false|false|false|C1704241|complex (molecular entity)|complex
Event|Event|History of Present Illness|2056,2063|false|false|false|||complex
Disorder|Anatomical Abnormality|History of Present Illness|2068,2072|false|false|false|C0010709|Cyst|cyst
Event|Event|History of Present Illness|2068,2072|false|false|false|||cyst
Finding|Body Substance|History of Present Illness|2068,2072|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Finding|Intellectual Product|History of Present Illness|2068,2072|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Finding|Body Substance|History of Present Illness|2080,2087|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|2080,2087|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|2080,2087|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|2092,2102|false|false|false|||transfused
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|2119,2124|false|false|false|C2316467|Packed red blood cells|pRBCs
Drug|Pharmacologic Substance|History of Present Illness|2119,2124|false|false|false|C2316467|Packed red blood cells|pRBCs
Event|Event|History of Present Illness|2144,2152|false|false|false|||increase
Finding|Functional Concept|History of Present Illness|2144,2152|false|false|false|C0442805|Increase|increase
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|2156,2159|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|History of Present Illness|2156,2159|false|false|false|C0019046|Hemoglobin|Hgb
Event|Event|History of Present Illness|2156,2159|false|false|false|||Hgb
Finding|Gene or Genome|History of Present Illness|2156,2159|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|History of Present Illness|2156,2159|false|false|false|C0019029|Hemoglobin concentration|Hgb
Event|Event|History of Present Illness|2178,2189|false|false|false|||transfusion
Finding|Functional Concept|History of Present Illness|2178,2189|false|false|false|C0199960||transfusion
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|2178,2189|false|false|false|C0005841;C1879316|Blood Transfusion;Transfusion (procedure)|transfusion
Finding|Functional Concept|History of Present Illness|2194,2200|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Event|Event|History of Present Illness|2201,2204|false|false|false|||CXR
Procedure|Diagnostic Procedure|History of Present Illness|2201,2204|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|History of Present Illness|2209,2216|false|false|false|||notable
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2221,2230|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|History of Present Illness|2221,2230|false|false|false|C2707265||pulmonary
Finding|Finding|History of Present Illness|2221,2230|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|History of Present Illness|2221,2236|false|false|false|C0034063|Pulmonary Edema|pulmonary edema
Attribute|Clinical Attribute|History of Present Illness|2231,2236|false|false|false|C1717255||edema
Event|Event|History of Present Illness|2231,2236|false|false|false|||edema
Finding|Pathologic Function|History of Present Illness|2231,2236|false|false|false|C0013604|Edema|edema
Anatomy|Tissue|History of Present Illness|2253,2260|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|History of Present Illness|2253,2260|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Pathologic Function|History of Present Illness|2253,2270|false|false|false|C0032227|Pleural effusion (disorder)|pleural effusions
Event|Event|History of Present Illness|2261,2270|false|false|false|||effusions
Finding|Pathologic Function|History of Present Illness|2261,2270|false|false|false|C0013687|effusion|effusions
Drug|Organic Chemical|History of Present Illness|2294,2299|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|History of Present Illness|2294,2299|false|false|false|C0699992|Lasix|Lasix
Drug|Organic Chemical|History of Present Illness|2312,2317|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|History of Present Illness|2312,2317|false|false|false|C0699992|Lasix|Lasix
Event|Event|History of Present Illness|2334,2342|false|false|false|||decision
Finding|Mental Process|History of Present Illness|2334,2342|false|false|false|C0679006|Decision|decision
Procedure|Health Care Activity|History of Present Illness|2355,2360|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admit
Finding|Body Substance|History of Present Illness|2365,2372|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|2365,2372|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|2365,2372|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Disorder|Disease or Syndrome|History of Present Illness|2377,2383|false|false|false|C0002871|Anemia|anemia
Event|Event|History of Present Illness|2377,2383|false|false|false|||anemia
Event|Event|History of Present Illness|2389,2394|false|false|false|||flash
Finding|Gene or Genome|History of Present Illness|2389,2394|false|false|false|C1413133;C4284306|CASP8AP2 gene;CASP8AP2 wt Allele|flash
Procedure|Diagnostic Procedure|History of Present Illness|2389,2394|false|false|false|C0262485|Flash|flash
Disorder|Disease or Syndrome|History of Present Illness|2389,2410|false|false|false|C1168329|Flash pulmonary oedema|flash pulmonary edema
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2395,2404|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|History of Present Illness|2395,2404|false|false|false|C2707265||pulmonary
Finding|Finding|History of Present Illness|2395,2404|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|History of Present Illness|2395,2410|false|false|false|C0034063|Pulmonary Edema|pulmonary edema
Attribute|Clinical Attribute|History of Present Illness|2405,2410|false|false|false|C1717255||edema
Event|Event|History of Present Illness|2405,2410|false|false|false|||edema
Finding|Pathologic Function|History of Present Illness|2405,2410|false|false|false|C0013604|Edema|edema
Anatomy|Anatomical Structure|History of Present Illness|2421,2426|false|false|false|C3714591|Floor (anatomic)|floor
Event|Event|History of Present Illness|2435,2442|false|false|false|||notable
Event|Event|History of Present Illness|2488,2492|false|false|false|||FSBG
Event|Event|History of Present Illness|2502,2509|false|false|false|||reports
Finding|Intellectual Product|History of Present Illness|2513,2518|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|History of Present Illness|2519,2529|false|false|false|||complaints
Finding|Finding|History of Present Illness|2519,2529|false|false|false|C5441521|Complaint (finding)|complaints
Event|Event|History of Present Illness|2545,2554|false|false|false|||shortness
Attribute|Clinical Attribute|History of Present Illness|2545,2564|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|History of Present Illness|2545,2564|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|History of Present Illness|2558,2564|false|false|false|C0225386|Breath|breath
Event|Event|History of Present Illness|2569,2577|false|false|false|||resolved
Event|Event|History of Present Illness|2583,2589|false|false|false|||denies
Anatomy|Body Location or Region|History of Present Illness|2590,2595|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|2590,2595|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|2590,2600|true|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|2590,2600|true|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|2596,2600|true|false|false|C2598155||pain
Event|Event|History of Present Illness|2596,2600|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|2596,2600|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|2596,2600|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|2603,2612|false|false|false|||dizziness
Finding|Sign or Symptom|History of Present Illness|2603,2612|false|false|false|C0012833;C0042571|Dizziness;Vertigo|dizziness
Event|Event|History of Present Illness|2614,2629|false|false|false|||lightheadedness
Finding|Sign or Symptom|History of Present Illness|2614,2629|false|false|false|C0220870|Lightheadedness|lightheadedness
Disorder|Disease or Syndrome|Past Medical History|2657,2669|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|Past Medical History|2657,2669|false|false|false|||hypertension
Disorder|Disease or Syndrome|Past Medical History|2674,2682|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|diabetes
Event|Event|Past Medical History|2674,2682|false|false|false|||diabetes
Disorder|Disease or Syndrome|Past Medical History|2690,2693|false|false|false|C0001365;C0038454|Acute ill-defined cerebrovascular disease;Cerebrovascular accident|CVA
Drug|Pharmacologic Substance|Past Medical History|2690,2693|false|false|false|C5779650|Cyclophosphamide/Doxorubicin/Vincristine|CVA
Event|Event|Past Medical History|2690,2693|false|false|false|||CVA
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2695,2705|false|false|false|C0007765|Cerebellum|cerebellar
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2706,2715|false|false|false|C0001629;C0025148;C1550278|Adrenal Medulla;Medulla Oblongata;Medullary - body parts|medullary
Disorder|Disease or Syndrome|Past Medical History|2716,2722|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|Past Medical History|2716,2722|false|false|false|||stroke
Finding|Finding|Past Medical History|2716,2722|false|false|false|C5977286|Stroke (heart beat)|stroke
Disorder|Disease or Syndrome|Past Medical History|2734,2737|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Past Medical History|2734,2737|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Past Medical History|2734,2737|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Past Medical History|2734,2737|false|false|false|||CAD
Finding|Gene or Genome|Past Medical History|2734,2737|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Past Medical History|2734,2737|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Past Medical History|2734,2737|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2734,2737|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|Past Medical History|2755,2758|false|false|false|C0006430|Burning Mouth Syndrome|BMS
Event|Event|Past Medical History|2755,2758|false|false|false|||BMS
Disorder|Disease or Syndrome|Past Medical History|2790,2817|false|false|false|C0085096;C1704436|Peripheral Arterial Diseases;Peripheral Vascular Diseases|peripheral arterial disease
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2801,2809|false|false|false|C0003842|Arteries|arterial
Disorder|Disease or Syndrome|Past Medical History|2801,2817|false|false|false|C0852949|Arteriopathic disease|arterial disease
Disorder|Disease or Syndrome|Past Medical History|2810,2817|false|false|false|C0012634|Disease|disease
Event|Event|Past Medical History|2810,2817|false|false|false|||disease
Disorder|Disease or Syndrome|Past Medical History|2819,2831|false|true|false|C0021775|Intermittent Claudication|claudication
Event|Event|Past Medical History|2819,2831|false|false|false|||claudication
Finding|Finding|Past Medical History|2819,2831|false|true|false|C0311395;C1456822|Claudication (finding);Lameness|claudication
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2846,2854|false|false|false|C0005847|Blood Vessel|vascular
Event|Event|Past Medical History|2856,2863|false|false|false|||managed
Attribute|Clinical Attribute|Past Medical History|2881,2886|false|false|false|C1300072|Tumor stage|stage
Finding|Intellectual Product|Past Medical History|2881,2889|false|false|false|C0441772|Stage level 4|stage IV
Disorder|Disease or Syndrome|Past Medical History|2890,2893|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Event|Event|Past Medical History|2890,2893|false|false|false|||CKD
Drug|Biomedical or Dental Material|Past Medical History|2895,2903|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|Past Medical History|2895,2903|false|false|false|||baseline
Finding|Idea or Concept|Past Medical History|2895,2903|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Disorder|Disease or Syndrome|Past Medical History|2917,2921|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|Past Medical History|2917,2921|false|false|false|||GERD
Disorder|Disease or Syndrome|Past Medical History|2922,2932|false|false|false|C0014852|Esophageal Diseases|esophageal
Disorder|Disease or Syndrome|Past Medical History|2922,2938|false|false|false|C0267081|Terminal esophageal web|esophageal rings
Event|Event|Past Medical History|2933,2938|false|false|false|||rings
Event|Activity|Family Medical History|2992,2996|false|false|false|C1947906|Sorting|sort
Event|Event|Family Medical History|2992,2996|false|false|false|||sort
Finding|Cell Function|Family Medical History|2992,2996|false|false|false|C0237886;C0700314|Sorting (Cognition);Sorting - Cell Movement|sort
Finding|Mental Process|Family Medical History|2992,2996|false|false|false|C0237886;C0700314|Sorting (Cognition);Sorting - Cell Movement|sort
Disorder|Neoplastic Process|Family Medical History|3000,3006|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Family Medical History|3000,3006|false|false|false|||cancer
Finding|Conceptual Entity|Family Medical History|3008,3014|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|Family Medical History|3008,3014|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Event|Event|Family Medical History|3015,3019|false|false|false|||died
Anatomy|Body Location or Region|Family Medical History|3039,3043|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3039,3043|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Family Medical History|3039,3043|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Family Medical History|3039,3043|false|false|false|C0740941|Lung Problem|lung
Disorder|Disease or Syndrome|Family Medical History|3039,3051|false|false|false|C0024115|Lung diseases|lung disease
Disorder|Disease or Syndrome|Family Medical History|3044,3051|false|false|false|C0012634|Disease|disease
Event|Event|Family Medical History|3044,3051|false|false|false|||disease
Finding|Idea or Concept|Family Medical History|3054,3060|false|false|false|C1546508|Relationship - Mother|Mother
Event|Event|Family Medical History|3061,3065|false|false|false|||died
Drug|Amino Acid, Peptide, or Protein|Family Medical History|3087,3094|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Immunologic Factor|Family Medical History|3087,3094|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Pharmacologic Substance|Family Medical History|3087,3094|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Event|Event|Family Medical History|3087,3094|false|false|false|||unknown
Finding|Finding|Family Medical History|3087,3094|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Functional Concept|Family Medical History|3087,3094|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Idea or Concept|Family Medical History|3087,3094|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Intellectual Product|Family Medical History|3087,3094|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Event|Event|Family Medical History|3095,3100|false|false|false|||cause
Finding|Conceptual Entity|Family Medical History|3095,3100|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Finding|Functional Concept|Family Medical History|3095,3100|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Disorder|Disease or Syndrome|Family Medical History|3113,3116|true|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Family Medical History|3113,3116|true|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Family Medical History|3113,3116|true|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Family Medical History|3113,3116|false|false|false|||CAD
Finding|Gene or Genome|Family Medical History|3113,3116|true|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Family Medical History|3113,3116|true|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Family Medical History|3113,3116|true|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Family Medical History|3113,3116|true|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Finding|Pathologic Function|Family Medical History|3120,3140|true|false|false|C0085298|Sudden Cardiac Death|sudden cardiac death
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3127,3134|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|Family Medical History|3127,3134|false|false|false|C1314974|Cardiac attachment|cardiac
Finding|Pathologic Function|Family Medical History|3127,3140|true|false|false|C0376297|Cardiac Death|cardiac death
Event|Event|Family Medical History|3135,3140|false|false|false|||death
Finding|Finding|Family Medical History|3135,3140|false|false|false|C0011065;C1306577;C1546949|Cessation of life;Death (finding);Event Consequence - Death|death
Finding|Idea or Concept|Family Medical History|3135,3140|false|false|false|C0011065;C1306577;C1546949|Cessation of life;Death (finding);Event Consequence - Death|death
Finding|Organism Function|Family Medical History|3135,3140|false|false|false|C0011065;C1306577;C1546949|Cessation of life;Death (finding);Event Consequence - Death|death
Event|Event|Family Medical History|3157,3164|false|false|false|||history
Finding|Conceptual Entity|Family Medical History|3157,3164|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|3157,3164|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Family Medical History|3157,3164|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|3157,3167|true|false|false|C0262926|Medical History|history of
Disorder|Neoplastic Process|Family Medical History|3169,3175|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Family Medical History|3169,3175|false|false|false|||cancer
Procedure|Health Care Activity|General Exam|3194,3203|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|General Exam|3204,3212|false|false|false|||PHYSICAL
Finding|Finding|General Exam|3204,3212|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|General Exam|3204,3212|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|General Exam|3204,3212|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|General Exam|3204,3217|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|General Exam|3204,3217|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Event|Event|General Exam|3213,3217|false|false|false|||EXAM
Finding|Functional Concept|General Exam|3213,3217|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|3213,3217|false|false|false|C0582103|Medical Examination|EXAM
Event|Event|General Exam|3269,3273|false|false|false|||FSBG
Event|Event|General Exam|3280,3287|false|false|false|||General
Finding|Classification|General Exam|3280,3287|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|General Exam|3280,3287|false|false|false|C3812897|General medical service|General
Finding|Finding|General Exam|3289,3299|false|false|false|C0497406|Overweight|Overweight
Attribute|Clinical Attribute|General Exam|3307,3312|false|false|false|C5890168||alert
Drug|Organic Chemical|General Exam|3307,3312|false|false|false|C0718338|Alert brand of caffeine|alert
Drug|Pharmacologic Substance|General Exam|3307,3312|false|false|false|C0718338|Alert brand of caffeine|alert
Event|Event|General Exam|3307,3312|false|false|false|||alert
Finding|Finding|General Exam|3307,3312|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Functional Concept|General Exam|3307,3312|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Intellectual Product|General Exam|3307,3312|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Event|Event|General Exam|3314,3322|false|false|false|||oriented
Finding|Finding|General Exam|3314,3322|false|false|false|C1961028|Oriented to place|oriented
Finding|Intellectual Product|General Exam|3327,3332|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|General Exam|3333,3341|false|false|false|||distress
Finding|Finding|General Exam|3333,3341|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|General Exam|3333,3341|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|General Exam|3344,3349|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|General Exam|3351,3357|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|General Exam|3351,3357|false|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|General Exam|3351,3357|false|false|false|||Sclera
Procedure|Health Care Activity|General Exam|3351,3357|false|false|false|C2228481|examination of sclera|Sclera
Event|Event|General Exam|3358,3367|false|false|false|||anicteric
Finding|Finding|General Exam|3358,3367|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|General Exam|3369,3372|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|General Exam|3369,3372|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Location or Region|General Exam|3374,3384|false|false|false|C0521367|Oropharyngeal|oropharynx
Event|Event|General Exam|3385,3390|false|false|false|||clear
Finding|Idea or Concept|General Exam|3385,3390|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Location or Region|General Exam|3393,3397|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|General Exam|3393,3397|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|General Exam|3393,3397|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|General Exam|3399,3405|false|false|false|||supple
Finding|Functional Concept|General Exam|3399,3405|false|false|false|C0332254|Supple|supple
Event|Event|General Exam|3407,3410|false|false|false|||JVP
Finding|Finding|General Exam|3407,3410|false|false|false|C0428897|Jugular venous pressure|JVP
Event|Event|General Exam|3415,3423|false|false|false|||elevated
Anatomy|Body Part, Organ, or Organ Component|General Exam|3426,3431|false|false|false|C0024109|Lung|Lungs
Event|Event|General Exam|3433,3441|false|false|false|||Crackles
Finding|Finding|General Exam|3433,3441|false|false|false|C0034642;C0240859|Basilar Rales;Rales|Crackles
Event|Activity|General Exam|3485,3489|false|false|false|C0871208|Rating (action)|rate
Event|Event|General Exam|3485,3489|false|false|false|||rate
Finding|Idea or Concept|General Exam|3485,3489|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|General Exam|3494,3500|false|false|false|||rhythm
Finding|Finding|General Exam|3494,3500|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|General Exam|3494,3500|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Event|Event|General Exam|3521,3528|false|false|false|||murmurs
Finding|Finding|General Exam|3521,3528|true|false|false|C0018808|Heart murmur|murmurs
Event|Event|General Exam|3533,3540|false|false|false|||gallops
Anatomy|Body Location or Region|General Exam|3543,3550|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|General Exam|3543,3550|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Event|Event|General Exam|3543,3550|false|false|false|||Abdomen
Finding|Finding|General Exam|3543,3550|false|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|General Exam|3552,3556|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|General Exam|3552,3556|false|false|false|||soft
Anatomy|Body Part, Organ, or Organ Component|General Exam|3585,3590|false|false|false|C0021853|Intestines|bowel
Finding|Finding|General Exam|3585,3597|false|false|false|C0232693|Bowel sounds|bowel sounds
Event|Event|General Exam|3591,3597|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|General Exam|3591,3597|false|false|false|C0037709||sounds
Finding|Finding|General Exam|3598,3605|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|General Exam|3598,3605|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Sign or Symptom|General Exam|3611,3629|true|false|false|C0234246|Rebound tenderness|rebound tenderness
Event|Event|General Exam|3619,3629|false|false|false|||tenderness
Finding|Mental Process|General Exam|3619,3629|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|General Exam|3619,3629|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Event|General Exam|3633,3641|false|false|false|||guarding
Finding|Finding|General Exam|3633,3641|true|false|false|C0427198|Protective muscle spasm|guarding
Event|Event|General Exam|3646,3658|false|false|false|||organomegaly
Finding|Finding|General Exam|3646,3658|true|false|false|C4054315|Organomegaly|organomegaly
Disorder|Congenital Abnormality|General Exam|3661,3664|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|General Exam|3661,3664|false|false|false|||Ext
Finding|Gene or Genome|General Exam|3661,3664|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|General Exam|3666,3670|false|false|false|||Warm
Finding|Finding|General Exam|3666,3670|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|3666,3670|false|false|false|C0687712|warming process|Warm
Finding|Finding|General Exam|3672,3676|false|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|3677,3685|false|false|false|||perfused
Drug|Food|General Exam|3690,3696|false|false|false|C5890763||pulses
Event|Event|General Exam|3690,3696|false|false|false|||pulses
Finding|Physiologic Function|General Exam|3690,3696|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|3690,3696|false|false|false|C0034107|Pulse taking|pulses
Disorder|Anatomical Abnormality|General Exam|3701,3709|true|false|false|C0149651|Clubbing|clubbing
Event|Event|General Exam|3701,3709|false|false|false|||clubbing
Event|Event|General Exam|3713,3721|false|false|false|||cyanosis
Finding|Sign or Symptom|General Exam|3713,3721|true|false|false|C0010520|Cyanosis|cyanosis
Finding|Functional Concept|General Exam|3727,3734|false|false|false|C0205323|Pitting|pitting
Finding|Finding|General Exam|3727,3740|false|false|false|C0333243|Pitting edema|pitting edema
Attribute|Clinical Attribute|General Exam|3735,3740|false|false|false|C1717255||edema
Event|Event|General Exam|3735,3740|false|false|false|||edema
Finding|Pathologic Function|General Exam|3735,3740|false|false|false|C0013604|Edema|edema
Finding|Functional Concept|General Exam|3744,3753|false|false|false|C3244310|dependent|dependent
Event|Event|General Exam|3754,3759|false|false|false|||areas
Anatomy|Body Location or Region|General Exam|3767,3775|false|false|false|C0006497|Buttocks|buttocks
Anatomy|Body System|General Exam|3778,3782|false|false|false|C1123023;C4520765|Skin;Skin, Human|Skin
Disorder|Disease or Syndrome|General Exam|3778,3782|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Disorder|Neoplastic Process|General Exam|3778,3782|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Finding|Body Substance|General Exam|3778,3782|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Finding|Intellectual Product|General Exam|3778,3782|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Event|Event|General Exam|3787,3793|false|false|false|||rashes
Finding|Sign or Symptom|General Exam|3787,3793|true|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Event|Event|General Exam|3794,3799|false|false|false|||noted
Event|Event|General Exam|3811,3819|false|false|false|||strength
Finding|Idea or Concept|General Exam|3811,3819|false|false|false|C0808080|Strength (attribute)|strength
Anatomy|Body Part, Organ, or Organ Component|General Exam|3823,3831|false|false|false|C0224234|Structure of deltoid muscle|deltoids
Anatomy|Body Part, Organ, or Organ Component|General Exam|3833,3839|false|false|false|C0559499|Biceps brachii muscle structure|biceps
Anatomy|Body Part, Organ, or Organ Component|General Exam|3841,3848|false|false|false|C0559502;C3146295|Triceps;Triceps brachii muscle structure|triceps
Anatomy|Body Location or Region|General Exam|3850,3855|false|false|false|C0043262;C1322271;C4298907|Upper extremity>Wrist;Wrist;Wrist joint|wrist
Anatomy|Body Space or Junction|General Exam|3850,3855|false|false|false|C0043262;C1322271;C4298907|Upper extremity>Wrist;Wrist;Wrist joint|wrist
Anatomy|Body Location or Region|General Exam|3857,3866|false|false|false|C1184148|Extensor|extensors
Anatomy|Body Part, Organ, or Organ Component|General Exam|3868,3874|false|false|false|C0016129;C0851278;C4299059|Fingers;Fingers not including thumb;Upper extremity>Finger|finger
Anatomy|Body Part, Organ, or Organ Component|General Exam|3868,3884|false|false|false|C5235530|Finger Extensors|finger extensors
Anatomy|Body Location or Region|General Exam|3875,3884|false|false|false|C1184148|Extensor|extensors
Anatomy|Body Part, Organ, or Organ Component|General Exam|3886,3889|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|General Exam|3886,3889|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|General Exam|3886,3889|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|General Exam|3886,3889|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|General Exam|3886,3889|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|General Exam|3886,3889|false|false|false|C1292890|Procedure on hip|hip
Event|Event|General Exam|3890,3897|false|false|false|||flexors
Anatomy|Body Part, Organ, or Organ Component|General Exam|3899,3909|false|false|false|C0584895|Posterior muscle of thigh structure|hamstrings
Anatomy|Body Part, Organ, or Organ Component|General Exam|3912,3922|false|false|false|C0224440|Structure of quadriceps femoris muscle|quadriceps
Event|Event|General Exam|3924,3932|false|false|false|||gastrocs
Anatomy|Body Part, Organ, or Organ Component|General Exam|3934,3942|false|false|false|C1710422|Tibialis Muscle|tibialis
Anatomy|Body Part, Organ, or Organ Component|General Exam|3934,3951|false|false|false|C0242690|Tibialis anterior muscle structure|tibialis anterior
Disorder|Disease or Syndrome|General Exam|3943,3951|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Event|Event|General Exam|3966,3975|false|false|false|||Sensation
Finding|Finding|General Exam|3966,3975|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Finding|Organ or Tissue Function|General Exam|3966,3975|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Procedure|Health Care Activity|General Exam|3966,3975|false|false|false|C2229507|sensory exam|Sensation
Event|Event|General Exam|3977,3983|false|false|false|||intact
Finding|Finding|General Exam|3977,3983|false|false|false|C1554187|Gender Status - Intact|intact
Disorder|Mental or Behavioral Dysfunction|General Exam|3998,4003|false|false|false|C0004936;C1306597|Mental disorders;Psychiatric problem|PSYCH
Event|Event|General Exam|3998,4003|false|false|false|||PSYCH
Attribute|Clinical Attribute|General Exam|4005,4010|false|false|false|C5890168||Alert
Drug|Organic Chemical|General Exam|4005,4010|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|General Exam|4005,4010|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|General Exam|4005,4010|false|false|false|||Alert
Finding|Finding|General Exam|4005,4010|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|General Exam|4005,4010|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|General Exam|4005,4010|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|General Exam|4021,4029|false|false|false|||oriented
Finding|Finding|General Exam|4021,4029|false|false|false|C1961028|Oriented to place|oriented
Attribute|Clinical Attribute|General Exam|4038,4042|false|false|false|C2713234||mood
Event|Event|General Exam|4038,4042|false|false|false|||mood
Finding|Conceptual Entity|General Exam|4038,4042|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|mood
Finding|Finding|General Exam|4038,4042|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|mood
Finding|Mental Process|General Exam|4038,4042|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|mood
Event|Event|General Exam|4047,4053|false|false|false|||affect
Finding|Mental Process|General Exam|4047,4053|false|false|false|C0001721|Affect (mental function)|affect
Procedure|Health Care Activity|General Exam|4047,4053|false|false|false|C2237113|assessment of affect|affect
Event|Event|General Exam|4073,4080|false|false|false|||respond
Event|Event|General Exam|4085,4095|false|false|false|||responding
Event|Event|General Exam|4112,4119|false|false|false|||answers
Event|Event|General Exam|4134,4145|false|false|false|||appropriate
Finding|Body Substance|General Exam|4147,4156|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|4147,4156|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|4147,4156|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|4147,4156|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|General Exam|4157,4165|false|false|false|||PHYSICAL
Finding|Finding|General Exam|4157,4165|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|General Exam|4157,4165|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|General Exam|4157,4165|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|General Exam|4157,4170|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|General Exam|4157,4170|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Event|Event|General Exam|4166,4170|false|false|false|||EXAM
Finding|Functional Concept|General Exam|4166,4170|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|4166,4170|false|false|false|C0582103|Medical Examination|EXAM
Attribute|Clinical Attribute|General Exam|4224,4228|false|false|false|C2317096|Saturation of Peripheral Oxygen|SPO2
Event|Event|General Exam|4236,4243|false|false|false|||General
Finding|Classification|General Exam|4236,4243|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|General Exam|4236,4243|false|false|false|C3812897|General medical service|General
Finding|Finding|General Exam|4245,4255|false|false|false|C0497406|Overweight|Overweight
Attribute|Clinical Attribute|General Exam|4263,4268|false|false|false|C5890168||alert
Drug|Organic Chemical|General Exam|4263,4268|false|false|false|C0718338|Alert brand of caffeine|alert
Drug|Pharmacologic Substance|General Exam|4263,4268|false|false|false|C0718338|Alert brand of caffeine|alert
Event|Event|General Exam|4263,4268|false|false|false|||alert
Finding|Finding|General Exam|4263,4268|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Functional Concept|General Exam|4263,4268|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Intellectual Product|General Exam|4263,4268|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Event|Event|General Exam|4270,4278|false|false|false|||oriented
Finding|Finding|General Exam|4270,4278|false|false|false|C1961028|Oriented to place|oriented
Finding|Intellectual Product|General Exam|4283,4288|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|General Exam|4289,4297|false|false|false|||distress
Finding|Finding|General Exam|4289,4297|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|General Exam|4289,4297|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|General Exam|4300,4305|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|General Exam|4307,4313|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|General Exam|4307,4313|false|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|General Exam|4307,4313|false|false|false|||Sclera
Procedure|Health Care Activity|General Exam|4307,4313|false|false|false|C2228481|examination of sclera|Sclera
Event|Event|General Exam|4314,4323|false|false|false|||anicteric
Finding|Finding|General Exam|4314,4323|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|General Exam|4325,4328|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|General Exam|4325,4328|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Location or Region|General Exam|4330,4340|false|false|false|C0521367|Oropharyngeal|oropharynx
Event|Event|General Exam|4341,4346|false|false|false|||clear
Finding|Idea or Concept|General Exam|4341,4346|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Location or Region|General Exam|4349,4353|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|General Exam|4349,4353|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|General Exam|4349,4353|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|General Exam|4355,4361|false|false|false|||supple
Finding|Functional Concept|General Exam|4355,4361|false|false|false|C0332254|Supple|supple
Event|Event|General Exam|4363,4366|false|false|false|||JVP
Finding|Finding|General Exam|4363,4366|false|false|false|C0428897|Jugular venous pressure|JVP
Event|Event|General Exam|4371,4379|false|false|false|||elevated
Anatomy|Body Part, Organ, or Organ Component|General Exam|4382,4387|false|false|false|C0024109|Lung|Lungs
Event|Event|General Exam|4389,4394|false|false|false|||Clear
Finding|Idea or Concept|General Exam|4389,4394|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|General Exam|4398,4410|false|false|false|||auscultation
Procedure|Diagnostic Procedure|General Exam|4398,4410|false|false|false|C0004339|Auscultation|auscultation
Event|Activity|General Exam|4435,4439|false|false|false|C0871208|Rating (action)|rate
Event|Event|General Exam|4435,4439|false|false|false|||rate
Finding|Idea or Concept|General Exam|4435,4439|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|General Exam|4444,4450|false|false|false|||rhythm
Finding|Finding|General Exam|4444,4450|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|General Exam|4444,4450|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Event|Event|General Exam|4471,4478|false|false|false|||murmurs
Finding|Finding|General Exam|4471,4478|true|false|false|C0018808|Heart murmur|murmurs
Event|Event|General Exam|4483,4490|false|false|false|||gallops
Anatomy|Body Location or Region|General Exam|4493,4500|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|General Exam|4493,4500|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Event|Event|General Exam|4493,4500|false|false|false|||Abdomen
Finding|Finding|General Exam|4493,4500|false|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|General Exam|4502,4506|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|General Exam|4502,4506|false|false|false|||soft
Anatomy|Body Part, Organ, or Organ Component|General Exam|4535,4540|false|false|false|C0021853|Intestines|bowel
Finding|Finding|General Exam|4535,4547|false|false|false|C0232693|Bowel sounds|bowel sounds
Event|Event|General Exam|4541,4547|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|General Exam|4541,4547|false|false|false|C0037709||sounds
Finding|Finding|General Exam|4548,4555|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|General Exam|4548,4555|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Sign or Symptom|General Exam|4561,4579|true|false|false|C0234246|Rebound tenderness|rebound tenderness
Event|Event|General Exam|4569,4579|false|false|false|||tenderness
Finding|Mental Process|General Exam|4569,4579|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|General Exam|4569,4579|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Event|General Exam|4583,4591|false|false|false|||guarding
Finding|Finding|General Exam|4583,4591|true|false|false|C0427198|Protective muscle spasm|guarding
Event|Event|General Exam|4596,4608|false|false|false|||organomegaly
Finding|Finding|General Exam|4596,4608|true|false|false|C4054315|Organomegaly|organomegaly
Disorder|Congenital Abnormality|General Exam|4611,4614|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|General Exam|4611,4614|false|false|false|||Ext
Finding|Gene or Genome|General Exam|4611,4614|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|General Exam|4616,4620|false|false|false|||Warm
Finding|Finding|General Exam|4616,4620|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|4616,4620|false|false|false|C0687712|warming process|Warm
Finding|Finding|General Exam|4622,4626|false|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|4627,4635|false|false|false|||perfused
Drug|Food|General Exam|4640,4646|false|false|false|C5890763||pulses
Event|Event|General Exam|4640,4646|false|false|false|||pulses
Finding|Physiologic Function|General Exam|4640,4646|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|4640,4646|false|false|false|C0034107|Pulse taking|pulses
Disorder|Anatomical Abnormality|General Exam|4651,4659|true|false|false|C0149651|Clubbing|clubbing
Event|Event|General Exam|4651,4659|false|false|false|||clubbing
Event|Event|General Exam|4663,4671|false|false|false|||cyanosis
Finding|Sign or Symptom|General Exam|4663,4671|true|false|false|C0010520|Cyanosis|cyanosis
Finding|Functional Concept|General Exam|4677,4684|false|false|false|C0205323|Pitting|pitting
Finding|Finding|General Exam|4677,4690|false|false|false|C0333243|Pitting edema|pitting edema
Attribute|Clinical Attribute|General Exam|4685,4690|false|false|false|C1717255||edema
Event|Event|General Exam|4685,4690|false|false|false|||edema
Finding|Pathologic Function|General Exam|4685,4690|false|false|false|C0013604|Edema|edema
Anatomy|Body Location or Region|General Exam|4694,4699|false|false|false|C0230444|Shin|shins
Anatomy|Body System|General Exam|4712,4716|false|false|false|C1123023;C4520765|Skin;Skin, Human|Skin
Disorder|Disease or Syndrome|General Exam|4712,4716|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Disorder|Neoplastic Process|General Exam|4712,4716|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Finding|Body Substance|General Exam|4712,4716|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Finding|Intellectual Product|General Exam|4712,4716|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Event|Event|General Exam|4721,4727|false|false|false|||rashes
Finding|Sign or Symptom|General Exam|4721,4727|true|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Event|Event|General Exam|4728,4733|false|false|false|||noted
Attribute|Clinical Attribute|General Exam|4756,4766|false|false|false|C2598148||LABORATORY
Finding|Functional Concept|General Exam|4756,4766|false|false|false|C1548427;C1571737;C3244292|Diagnostic Service Section ID - Laboratory;Laboratory domain;Referral type - Laboratory|LABORATORY
Finding|Intellectual Product|General Exam|4756,4766|false|false|false|C1548427;C1571737;C3244292|Diagnostic Service Section ID - Laboratory;Laboratory domain;Referral type - Laboratory|LABORATORY
Lab|Laboratory or Test Result|General Exam|4756,4766|false|false|false|C4283904|Laboratory observation|LABORATORY
Procedure|Laboratory Procedure|General Exam|4756,4774|false|false|false|C0681827|laboratory studies|LABORATORY STUDIES
Event|Event|General Exam|4767,4774|false|false|false|||STUDIES
Procedure|Research Activity|General Exam|4767,4774|false|false|false|C0947630|Scientific Study|STUDIES
Procedure|Health Care Activity|General Exam|4778,4787|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Anatomy|Cell|General Exam|4848,4851|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|4856,4859|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|4856,4859|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|4856,4859|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|4866,4869|false|false|false|C0019046|Hemoglobin|HGB
Drug|Biologically Active Substance|General Exam|4866,4869|false|false|false|C0019046|Hemoglobin|HGB
Event|Event|General Exam|4866,4869|false|false|false|||HGB
Finding|Gene or Genome|General Exam|4866,4869|false|false|false|C1424337|CYGB gene|HGB
Lab|Laboratory or Test Result|General Exam|4866,4869|false|false|false|C0019029|Hemoglobin concentration|HGB
Procedure|Laboratory Procedure|General Exam|4875,4878|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|General Exam|4875,4878|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Disorder|Virus|General Exam|4886,4889|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|4886,4889|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|4886,4889|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|4886,4889|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|4886,4889|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|4896,4899|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|4896,4899|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|4896,4899|false|false|false|||MCH
Finding|Gene or Genome|General Exam|4896,4899|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|4896,4899|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|4896,4899|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|4905,4909|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|4905,4909|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Drug|Amino Acid, Peptide, or Protein|General Exam|4970,4977|false|false|false|C0001924;C5966160|Albumin;Albumins|ALBUMIN
Drug|Biologically Active Substance|General Exam|4970,4977|false|false|false|C0001924;C5966160|Albumin;Albumins|ALBUMIN
Drug|Pharmacologic Substance|General Exam|4970,4977|false|false|false|C0001924;C5966160|Albumin;Albumins|ALBUMIN
Event|Event|General Exam|4970,4977|false|false|false|||ALBUMIN
Finding|Gene or Genome|General Exam|4970,4977|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|ALBUMIN
Finding|Physiologic Function|General Exam|4970,4977|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|ALBUMIN
Procedure|Laboratory Procedure|General Exam|4970,4977|false|false|false|C0201838|Albumin measurement|ALBUMIN
Drug|Biologically Active Substance|General Exam|4982,4989|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Element, Ion, or Isotope|General Exam|4982,4989|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Inorganic Chemical|General Exam|4982,4989|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Pharmacologic Substance|General Exam|4982,4989|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Vitamin|General Exam|4982,4989|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Event|Event|General Exam|4982,4989|false|false|false|||CALCIUM
Finding|Physiologic Function|General Exam|4982,4989|false|false|false|C4553026|Calcium metabolic function|CALCIUM
Procedure|Laboratory Procedure|General Exam|4982,4989|false|false|false|C0201925|Calcium measurement|CALCIUM
Drug|Element, Ion, or Isotope|General Exam|4994,5003|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Drug|Inorganic Chemical|General Exam|4994,5003|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Drug|Pharmacologic Substance|General Exam|4994,5003|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Procedure|Laboratory Procedure|General Exam|4994,5003|false|false|false|C0523826|Phosphate measurement|PHOSPHATE
Drug|Biologically Active Substance|General Exam|5010,5014|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|IRON
Drug|Element, Ion, or Isotope|General Exam|5010,5014|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|IRON
Drug|Pharmacologic Substance|General Exam|5010,5014|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|IRON
Event|Event|General Exam|5010,5014|false|false|false|||IRON
Procedure|Laboratory Procedure|General Exam|5010,5014|false|false|false|C0337439|Iron measurement|IRON
Drug|Amino Acid, Peptide, or Protein|General Exam|5044,5052|false|false|false|C0015879|Ferritin|FERRITIN
Drug|Biologically Active Substance|General Exam|5044,5052|false|false|false|C0015879|Ferritin|FERRITIN
Drug|Pharmacologic Substance|General Exam|5044,5052|false|false|false|C0015879|Ferritin|FERRITIN
Event|Event|General Exam|5044,5052|false|false|false|||FERRITIN
Procedure|Laboratory Procedure|General Exam|5044,5052|false|false|false|C0373607|Ferritin measurement|FERRITIN
Drug|Amino Acid, Peptide, or Protein|General Exam|5058,5061|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Biologically Active Substance|General Exam|5058,5061|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Hormone|General Exam|5058,5061|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Pharmacologic Substance|General Exam|5058,5061|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Event|Event|General Exam|5058,5061|false|false|false|||TRF
Finding|Gene or Genome|General Exam|5058,5061|false|false|false|C1334121;C1336604;C1705002|IL5 gene;TERF1 gene;TERF1 wt Allele|TRF
Drug|Biologically Active Substance|General Exam|5080,5084|false|false|false|C0041942|urea|UREA
Drug|Organic Chemical|General Exam|5080,5084|false|false|false|C0041942|urea|UREA
Drug|Pharmacologic Substance|General Exam|5080,5084|false|false|false|C0041942|urea|UREA
Event|Event|General Exam|5080,5084|false|false|false|||UREA
Procedure|Laboratory Procedure|General Exam|5080,5084|false|false|false|C0523961|Urea measurement|UREA
Drug|Biologically Active Substance|General Exam|5102,5108|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Element, Ion, or Isotope|General Exam|5102,5108|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Pharmacologic Substance|General Exam|5102,5108|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Event|Event|General Exam|5102,5108|false|false|false|||SODIUM
Finding|Physiologic Function|General Exam|5102,5108|false|false|false|C4553025|Sodium metabolic function|SODIUM
Procedure|Laboratory Procedure|General Exam|5102,5108|false|false|false|C0337443|Sodium measurement|SODIUM
Drug|Biologically Active Substance|General Exam|5114,5123|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Element, Ion, or Isotope|General Exam|5114,5123|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Food|General Exam|5114,5123|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Inorganic Chemical|General Exam|5114,5123|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Pharmacologic Substance|General Exam|5114,5123|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Event|Event|General Exam|5114,5123|false|false|false|||POTASSIUM
Finding|Physiologic Function|General Exam|5114,5123|false|false|false|C4553027|Potassium metabolic function|POTASSIUM
Procedure|Laboratory Procedure|General Exam|5114,5123|false|false|false|C0202194|Potassium measurement|POTASSIUM
Drug|Element, Ion, or Isotope|General Exam|5128,5136|false|false|false|C0008203;C0596019|Chlorides;chloride ion|CHLORIDE
Event|Event|General Exam|5128,5136|false|false|false|||CHLORIDE
Finding|Physiologic Function|General Exam|5128,5136|false|false|false|C4553021|Chloride metabolic function|CHLORIDE
Procedure|Laboratory Procedure|General Exam|5128,5136|false|false|false|C0201952|Chloride measurement|CHLORIDE
Drug|Biologically Active Substance|General Exam|5148,5151|false|false|false|C0007012|carbon dioxide|CO2
Drug|Inorganic Chemical|General Exam|5148,5151|false|false|false|C0007012|carbon dioxide|CO2
Event|Event|General Exam|5148,5151|false|false|false|||CO2
Finding|Finding|General Exam|5148,5151|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Finding|Gene or Genome|General Exam|5148,5151|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Drug|Element, Ion, or Isotope|General Exam|5155,5160|false|false|false|C0003075|Anions|ANION
Attribute|Clinical Attribute|General Exam|5155,5164|false|false|false|C0003074|Anion Gap|ANION GAP
Lab|Laboratory or Test Result|General Exam|5155,5164|false|false|false|C1509129|Anion gap result|ANION GAP
Procedure|Laboratory Procedure|General Exam|5155,5164|false|false|false|C0201889;C2189246|Anion gap measurement;blood anion gap (lab test)|ANION GAP
Drug|Amino Acid, Peptide, or Protein|General Exam|5161,5164|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Drug|Biologically Active Substance|General Exam|5161,5164|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Event|Event|General Exam|5161,5164|false|false|false|||GAP
Finding|Gene or Genome|General Exam|5161,5164|false|false|false|C1419277;C2984552|RASA1 gene;RASA1 wt Allele|GAP
Event|Event|General Exam|5198,5202|false|false|false|||BILI
Event|Event|General Exam|5236,5243|false|false|false|||IMAGING
Finding|Finding|General Exam|5236,5243|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|General Exam|5236,5243|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Attribute|Clinical Attribute|General Exam|5322,5326|false|false|false|C4318566|Deep Resection Margin|deep
Anatomy|Body Part, Organ, or Organ Component|General Exam|5322,5331|false|false|false|C0226514|Structure of deep vein|deep vein
Disorder|Disease or Syndrome|General Exam|5322,5342|false|false|false|C0149871;C0340708|Deep Vein Thrombosis;Deep vein thrombosis of lower limb|deep vein thrombosis
Anatomy|Body Part, Organ, or Organ Component|General Exam|5327,5331|false|false|false|C0042449|Veins|vein
Finding|Pathologic Function|General Exam|5327,5342|false|false|false|C0042487|Venous Thrombosis|vein thrombosis
Event|Event|General Exam|5332,5342|false|false|false|||thrombosis
Finding|Pathologic Function|General Exam|5332,5342|false|false|false|C0040053|Thrombosis|thrombosis
Disorder|Disease or Syndrome|General Exam|5365,5374|false|false|false|C0751438|Posterior pituitary disease|posterior
Event|Event|General Exam|5365,5374|false|false|false|||posterior
Anatomy|Body Part, Organ, or Organ Component|General Exam|5365,5387|false|false|false|C0226832|Structure of posterior tibial vein|posterior tibial veins
Anatomy|Body Part, Organ, or Organ Component|General Exam|5375,5381|false|false|false|C0040184|Bone structure of tibia|tibial
Anatomy|Body Part, Organ, or Organ Component|General Exam|5375,5387|false|false|false|C0447138|Tibial vein structure|tibial veins
Anatomy|Body Part, Organ, or Organ Component|General Exam|5382,5387|false|false|false|C0042449|Veins|veins
Event|Event|General Exam|5382,5387|false|false|false|||veins
Procedure|Therapeutic or Preventive Procedure|General Exam|5382,5387|false|false|false|C0398102|Procedure on vein|veins
Event|Event|General Exam|5416,5424|false|false|false|||thrombus
Finding|Pathologic Function|General Exam|5416,5424|false|false|false|C0087086;C0302148|Blood Clot;Thrombus|thrombus
Event|Event|General Exam|5442,5451|false|false|false|||decreased
Finding|Finding|General Exam|5457,5460|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|General Exam|5457,5460|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Attribute|Clinical Attribute|General Exam|5461,5465|true|false|false|C4318566|Deep Resection Margin|deep
Disorder|Disease or Syndrome|General Exam|5461,5483|true|false|false|C0149871|Deep Vein Thrombosis|deep venous thrombosis
Anatomy|Body Part, Organ, or Organ Component|General Exam|5466,5472|false|false|false|C0042449|Veins|venous
Finding|Finding|General Exam|5466,5483|true|false|false|C0042487;C0517555|Venous Thrombosis;Venous thrombosis after immobility|venous thrombosis
Finding|Pathologic Function|General Exam|5466,5483|true|false|false|C0042487;C0517555|Venous Thrombosis;Venous thrombosis after immobility|venous thrombosis
Event|Event|General Exam|5473,5483|false|false|false|||thrombosis
Finding|Pathologic Function|General Exam|5473,5483|true|false|false|C0040053|Thrombosis|thrombosis
Anatomy|Body Location or Region|General Exam|5495,5500|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|5495,5500|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|General Exam|5495,5510|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|General Exam|5501,5510|false|false|false|C0015385|Limb structure|extremity
Event|Event|General Exam|5516,5521|false|false|false|||Right
Finding|Functional Concept|General Exam|5516,5521|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Drug|Chemical Viewed Structurally|General Exam|5522,5529|false|false|false|C1704241|complex (molecular entity)|complex
Event|Event|General Exam|5522,5529|false|false|false|||complex
Disorder|Anatomical Abnormality|General Exam|5534,5538|false|false|false|C0010709|Cyst|cyst
Event|Event|General Exam|5534,5538|false|false|false|||cyst
Finding|Body Substance|General Exam|5534,5538|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Finding|Intellectual Product|General Exam|5534,5538|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Event|Event|General Exam|5542,5545|false|false|false|||CXR
Procedure|Diagnostic Procedure|General Exam|5542,5545|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Finding|General Exam|5557,5560|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Finding|Idea or Concept|General Exam|5557,5560|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Finding|Intellectual Product|General Exam|5561,5565|false|false|false|C1547225|Mild Severity of Illness Code|mild
Anatomy|Body Part, Organ, or Organ Component|General Exam|5566,5575|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|General Exam|5566,5575|false|false|false|C2707265||pulmonary
Finding|Finding|General Exam|5566,5575|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|General Exam|5566,5581|false|false|false|C0034063|Pulmonary Edema|pulmonary edema
Attribute|Clinical Attribute|General Exam|5576,5581|false|false|false|C1717255||edema
Event|Event|General Exam|5576,5581|false|false|false|||edema
Finding|Pathologic Function|General Exam|5576,5581|false|false|false|C0013604|Edema|edema
Event|Event|General Exam|5604,5613|false|false|false|||bilateral
Anatomy|Tissue|General Exam|5615,5622|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|General Exam|5615,5622|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Pathologic Function|General Exam|5615,5632|false|false|false|C0032227|Pleural effusion (disorder)|pleural effusions
Event|Event|General Exam|5623,5632|false|false|false|||effusions
Finding|Pathologic Function|General Exam|5623,5632|false|false|false|C0013687|effusion|effusions
Finding|Finding|General Exam|5638,5644|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Finding|Intellectual Product|General Exam|5638,5644|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Event|Event|General Exam|5645,5657|false|false|false|||cardiomegaly
Finding|Finding|General Exam|5645,5657|false|false|false|C0018800|Cardiomegaly|cardiomegaly
Finding|Finding|General Exam|5661,5667|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|General Exam|5661,5667|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|General Exam|5668,5679|false|false|false|||accentuated
Finding|Finding|General Exam|5687,5690|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|General Exam|5687,5690|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Anatomy|Body Location or Region|General Exam|5691,5695|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|General Exam|5691,5695|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|General Exam|5691,5695|false|false|false|C0024115|Lung diseases|lung
Event|Event|General Exam|5691,5695|false|false|false|||lung
Finding|Finding|General Exam|5691,5695|false|false|false|C0740941|Lung Problem|lung
Event|Event|General Exam|5697,5704|false|false|false|||volumes
Finding|Body Substance|General Exam|5709,5716|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|General Exam|5709,5716|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|General Exam|5709,5716|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Procedure|Health Care Activity|General Exam|5709,5728|false|false|false|C1561964|Positioning patient (procedure)|patient positioning
Event|Event|General Exam|5717,5728|false|false|false|||positioning
Procedure|Health Care Activity|General Exam|5717,5728|false|false|false|C0150305;C1561964|Positioning - therapy;Positioning patient (procedure)|positioning
Procedure|Therapeutic or Preventive Procedure|General Exam|5717,5728|false|false|false|C0150305;C1561964|Positioning - therapy;Positioning patient (procedure)|positioning
Event|Event|General Exam|5732,5735|false|false|false|||CXR
Procedure|Diagnostic Procedure|General Exam|5732,5735|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|General Exam|5746,5754|false|false|false|||compared
Anatomy|Body Location or Region|General Exam|5767,5771|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|General Exam|5767,5771|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|General Exam|5767,5771|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|General Exam|5767,5771|false|false|false|C0740941|Lung Problem|lung
Finding|Organ or Tissue Function|General Exam|5767,5779|false|false|false|C0231953|Lung Volumes|lung volumes
Event|Event|General Exam|5772,5779|false|false|false|||volumes
Event|Event|General Exam|5795,5804|false|false|false|||decreased
Event|Event|General Exam|5807,5812|false|false|false|||Signs
Finding|Finding|General Exam|5807,5812|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|Signs
Finding|Functional Concept|General Exam|5807,5812|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|Signs
Finding|Intellectual Product|General Exam|5816,5820|false|false|false|C1547225|Mild Severity of Illness Code|mild
Event|Event|General Exam|5821,5834|false|false|false|||overinflation
Finding|Finding|General Exam|5839,5847|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|General Exam|5839,5847|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Anatomy|Tissue|General Exam|5848,5855|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|General Exam|5848,5855|false|false|false|C0032226|Pleural Diseases|pleural
Event|Event|General Exam|5857,5866|false|false|false|||effusions
Finding|Pathologic Function|General Exam|5857,5866|false|false|false|C0013687|effusion|effusions
Event|Event|General Exam|5867,5874|false|false|false|||persist
Finding|Finding|General Exam|5877,5885|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|General Exam|5877,5885|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Event|Event|General Exam|5886,5898|false|false|false|||cardiomegaly
Finding|Finding|General Exam|5886,5898|false|false|false|C0018800|Cardiomegaly|cardiomegaly
Event|Event|General Exam|5901,5911|false|false|false|||Elongation
Finding|Functional Concept|General Exam|5920,5930|false|false|false|C1547177|Sequencing - Descending|descending
Anatomy|Body Part, Organ, or Organ Component|General Exam|5920,5936|false|false|false|C0011666;C1305624|Descending aorta|descending aorta
Anatomy|Body Part, Organ, or Organ Component|General Exam|5931,5936|false|false|false|C0003483;C4037978|Aorta;Chest+Abdomen>Aorta|aorta
Procedure|Health Care Activity|General Exam|5931,5936|false|false|false|C0869784|Procedure on aorta|aorta
Disorder|Disease or Syndrome|General Exam|5942,5951|true|false|false|C0032285|Pneumonia|pneumonia
Event|Event|General Exam|5942,5951|false|false|false|||pneumonia
Event|Event|General Exam|5966,5973|false|false|false|||STUDIES
Procedure|Research Activity|General Exam|5966,5973|false|false|false|C0947630|Scientific Study|STUDIES
Event|Event|General Exam|5977,5986|false|false|false|||DISCHARGE
Finding|Body Substance|General Exam|5977,5986|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|5977,5986|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|5977,5986|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|5977,5986|false|false|false|C0030685|Patient Discharge|DISCHARGE
Disorder|Disease or Syndrome|General Exam|6046,6051|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|6046,6051|false|false|false|||BLOOD
Finding|Body Substance|General Exam|6046,6051|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|6052,6055|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|6061,6064|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|6061,6064|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|6061,6064|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|6071,6074|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|6071,6074|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|6071,6074|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|6071,6074|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|6080,6083|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|6080,6083|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|6091,6094|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|6091,6094|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|6091,6094|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|6091,6094|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|6091,6094|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|6098,6101|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|6098,6101|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|6098,6101|false|false|false|||MCH
Finding|Gene or Genome|General Exam|6098,6101|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|6098,6101|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|6098,6101|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|6107,6111|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|6107,6111|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|6140,6143|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|6160,6165|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|6160,6165|false|false|false|||BLOOD
Finding|Body Substance|General Exam|6160,6165|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|6170,6173|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|General Exam|6170,6173|false|false|false|||PTT
Procedure|Laboratory Procedure|General Exam|6170,6173|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|General Exam|6195,6200|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|6195,6200|false|false|false|||BLOOD
Finding|Body Substance|General Exam|6195,6200|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|6195,6208|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|6195,6208|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|6195,6208|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|6201,6208|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|6201,6208|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|6201,6208|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|6201,6208|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|6201,6208|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|6201,6208|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|6256,6260|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|6256,6260|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|6256,6260|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|6285,6290|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|6285,6290|false|false|false|||BLOOD
Finding|Body Substance|General Exam|6285,6290|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|6294,6297|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Drug|Enzyme|General Exam|6294,6297|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Event|Event|General Exam|6294,6297|false|false|false|||LDH
Finding|Finding|General Exam|6294,6297|false|false|false|C0851148|Lifetime Drinking History|LDH
Procedure|Laboratory Procedure|General Exam|6294,6297|false|false|false|C0202113|Lactate dehydrogenase measurement|LDH
Disorder|Disease or Syndrome|General Exam|6327,6332|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|6327,6332|false|false|false|||BLOOD
Finding|Body Substance|General Exam|6327,6332|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|6327,6340|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|General Exam|6333,6340|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|6333,6340|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|6333,6340|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|6333,6340|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|6333,6340|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|General Exam|6333,6340|false|false|false|||Calcium
Finding|Physiologic Function|General Exam|6333,6340|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|6333,6340|false|false|false|C0201925|Calcium measurement|Calcium
Finding|Idea or Concept|Hospital Course|6404,6408|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|Hospital Course|6404,6408|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|Hospital Course|6409,6412|false|false|false|||old
Event|Event|Hospital Course|6431,6438|false|false|false|||medical
Finding|Functional Concept|Hospital Course|6431,6438|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|Hospital Course|6431,6438|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|Hospital Course|6431,6438|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|Hospital Course|6431,6438|false|false|false|C0199168|Medical service|medical
Event|Event|Hospital Course|6440,6447|false|false|false|||history
Finding|Conceptual Entity|Hospital Course|6440,6447|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|6440,6447|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|6440,6447|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|6440,6450|false|false|false|C0262926|Medical History|history of
Finding|Gene or Genome|Hospital Course|6451,6455|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Intellectual Product|Hospital Course|6451,6455|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Disorder|Disease or Syndrome|Hospital Course|6462,6474|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|Hospital Course|6462,6474|false|false|false|||hypertension
Attribute|Clinical Attribute|Hospital Course|6476,6481|false|false|false|C1300072|Tumor stage|stage
Finding|Intellectual Product|Hospital Course|6476,6484|false|false|false|C0441772|Stage level 4|stage IV
Disorder|Disease or Syndrome|Hospital Course|6485,6488|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Event|Event|Hospital Course|6485,6488|false|false|false|||CKD
Disorder|Disease or Syndrome|Hospital Course|6490,6493|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6490,6493|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|6490,6493|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Hospital Course|6490,6493|false|false|false|||CAD
Finding|Gene or Genome|Hospital Course|6490,6493|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|6490,6493|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|6490,6493|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6490,6493|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Finding|Pathologic Function|Hospital Course|6499,6506|false|false|false|C5441917|Distant Metastasis|distant
Drug|Inorganic Chemical|Hospital Course|6519,6524|false|false|false|C0025552|Metals|metal
Event|Event|Hospital Course|6525,6530|false|false|false|||stent
Disorder|Disease or Syndrome|Hospital Course|6532,6538|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|Hospital Course|6532,6538|false|false|false|||stroke
Finding|Finding|Hospital Course|6532,6538|false|false|false|C5977286|Stroke (heart beat)|stroke
Disorder|Disease or Syndrome|Hospital Course|6558,6562|false|false|false|C0151950|Deep thrombophlebitis|DVTs
Event|Event|Hospital Course|6558,6562|false|false|false|||DVTs
Drug|Organic Chemical|Hospital Course|6567,6575|false|false|false|C0699129|Coumadin|Coumadin
Drug|Pharmacologic Substance|Hospital Course|6567,6575|false|false|false|C0699129|Coumadin|Coumadin
Procedure|Diagnostic Procedure|Hospital Course|6588,6596|false|false|false|C0203057|Upper gastrointestinal tract series|upper GI
Finding|Pathologic Function|Hospital Course|6588,6602|false|false|false|C0041909|Upper gastrointestinal hemorrhage|upper GI bleed
Finding|Pathologic Function|Hospital Course|6594,6602|false|false|false|C0017181|Gastrointestinal Hemorrhage|GI bleed
Event|Event|Hospital Course|6597,6602|false|false|false|||bleed
Finding|Pathologic Function|Hospital Course|6597,6602|false|false|false|C0019080|Hemorrhage|bleed
Event|Event|Hospital Course|6612,6616|false|false|false|||sent
Attribute|Clinical Attribute|Hospital Course|6632,6641|false|false|false|C0804815||physician
Disorder|Disease or Syndrome|Hospital Course|6646,6652|false|false|false|C0002871|Anemia|anemia
Event|Event|Hospital Course|6646,6652|false|false|false|||anemia
Disorder|Disease or Syndrome|Hospital Course|6658,6664|false|false|false|C0002871|Anemia|Anemia
Event|Event|Hospital Course|6658,6664|false|false|false|||Anemia
Finding|Body Substance|Hospital Course|6667,6674|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|6667,6674|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|6667,6674|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|6675,6684|false|false|false|||presented
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6690,6693|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Hospital Course|6690,6693|false|false|false|C0019046|Hemoglobin|Hgb
Event|Event|Hospital Course|6690,6693|false|false|false|||Hgb
Finding|Gene or Genome|Hospital Course|6690,6693|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Hospital Course|6690,6693|false|false|false|C0019029|Hemoglobin concentration|Hgb
Drug|Biomedical or Dental Material|Hospital Course|6723,6731|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|Hospital Course|6723,6731|false|false|false|||baseline
Finding|Idea or Concept|Hospital Course|6723,6731|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|Hospital Course|6755,6770|false|false|false|||hospitalization
Procedure|Health Care Activity|Hospital Course|6755,6770|false|false|false|C0019993|Hospitalization|hospitalization
Event|Event|Hospital Course|6777,6789|false|false|false|||presentation
Finding|Idea or Concept|Hospital Course|6777,6789|false|false|false|C0449450|Presentation|presentation
Finding|Finding|Hospital Course|6801,6804|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Hospital Course|6801,6804|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Finding|Hospital Course|6805,6815|false|false|false|C0302845|Mean corpuscular volume above reference range|macrocytic
Disorder|Disease or Syndrome|Hospital Course|6805,6822|false|false|false|C0002886|Anemia, Macrocytic|macrocytic anemia
Finding|Gene or Genome|Hospital Course|6805,6822|false|false|false|C1420653|TCN2 gene|macrocytic anemia
Disorder|Disease or Syndrome|Hospital Course|6816,6822|false|false|false|C0002871|Anemia|anemia
Event|Event|Hospital Course|6816,6822|false|false|false|||anemia
Finding|Cell Function|Hospital Course|6824,6833|false|false|false|C0019054;C1553188;C2937287;C2945560|Hemolysis (biological function);Hemolysis (disorder);Hemolysis (finding)|Hemolysis
Finding|Finding|Hospital Course|6824,6833|false|false|false|C0019054;C1553188;C2937287;C2945560|Hemolysis (biological function);Hemolysis (disorder);Hemolysis (finding)|Hemolysis
Finding|Pathologic Function|Hospital Course|6824,6833|false|false|false|C0019054;C1553188;C2937287;C2945560|Hemolysis (biological function);Hemolysis (disorder);Hemolysis (finding)|Hemolysis
Event|Event|Hospital Course|6834,6838|false|false|false|||labs
Lab|Laboratory or Test Result|Hospital Course|6834,6838|false|false|false|C0587081|Laboratory test finding|labs
Event|Event|Hospital Course|6844,6852|false|false|false|||negative
Finding|Classification|Hospital Course|6844,6852|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|6844,6852|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|6844,6852|false|false|false|C5237010|Expression Negative|negative
Event|Event|Hospital Course|6859,6867|false|false|false|||received
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6881,6887|false|false|false|C0184967|Insertion of pack (procedure)|packed
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6881,6897|false|false|false|C2316467|Packed red blood cells|packed red cells
Drug|Pharmacologic Substance|Hospital Course|6881,6897|false|false|false|C2316467|Packed red blood cells|packed red cells
Finding|Finding|Hospital Course|6888,6891|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Finding|Gene or Genome|Hospital Course|6888,6891|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Anatomy|Cell|Hospital Course|6888,6897|false|false|false|C0014792|Erythrocytes|red cells
Drug|Pharmacologic Substance|Hospital Course|6888,6897|false|false|false|C0014792|Erythrocytes|red cells
Anatomy|Cell|Hospital Course|6892,6897|false|false|false|C0007634|Cells|cells
Event|Event|Hospital Course|6892,6897|false|false|false|||cells
Drug|Organic Chemical|Hospital Course|6918,6922|false|false|false|C0246719|risedronate|rise
Drug|Pharmacologic Substance|Hospital Course|6918,6922|false|false|false|C0246719|risedronate|rise
Event|Event|Hospital Course|6918,6922|false|false|false|||rise
Finding|Intellectual Product|Hospital Course|6918,6922|false|false|false|C4321377|Relational and Item-Specific Encoding Task|rise
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6931,6934|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Hospital Course|6931,6934|false|false|false|C0019046|Hemoglobin|Hgb
Event|Event|Hospital Course|6931,6934|false|false|false|||Hgb
Finding|Gene or Genome|Hospital Course|6931,6934|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Hospital Course|6931,6934|false|false|false|C0019029|Hemoglobin concentration|Hgb
Event|Event|Hospital Course|6943,6948|false|false|false|||Stool
Finding|Body Substance|Hospital Course|6943,6948|false|false|false|C0015733|Feces|Stool
Event|Event|Hospital Course|6959,6967|false|false|false|||negative
Finding|Classification|Hospital Course|6959,6967|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|6959,6967|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|6959,6967|false|false|false|C5237010|Expression Negative|negative
Event|Event|Hospital Course|6977,6984|false|false|false|||reports
Finding|Intellectual Product|Hospital Course|6977,6984|true|false|false|C0684224|Report (document)|reports
Procedure|Health Care Activity|Hospital Course|6977,6984|true|false|false|C0700287|Reporting|reports
Finding|Sign or Symptom|Hospital Course|6989,6999|false|false|false|C0474585||dark stool
Event|Event|Hospital Course|6994,6999|false|false|false|||stool
Finding|Body Substance|Hospital Course|6994,6999|false|false|false|C0015733|Feces|stool
Disorder|Disease or Syndrome|Hospital Course|7003,7008|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Hospital Course|7003,7008|false|false|false|||blood
Finding|Body Substance|Hospital Course|7003,7008|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Disorder|Disease or Syndrome|Hospital Course|7003,7017|false|false|false|C0018932|Hematochezia|blood in stool
Finding|Sign or Symptom|Hospital Course|7003,7017|false|false|false|C1321898|Blood in stool|blood in stool
Event|Event|Hospital Course|7012,7017|false|false|false|||stool
Finding|Body Substance|Hospital Course|7012,7017|false|false|false|C0015733|Feces|stool
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7023,7033|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Biologically Active Substance|Hospital Course|7023,7033|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Organic Chemical|Hospital Course|7023,7033|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Pharmacologic Substance|Hospital Course|7023,7033|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Event|Event|Hospital Course|7023,7033|false|false|false|||hemoglobin
Finding|Finding|Hospital Course|7023,7033|false|false|false|C1561562|Hemoglobin finding|hemoglobin
Procedure|Laboratory Procedure|Hospital Course|7023,7033|false|false|false|C0518015|Hemoglobin measurement|hemoglobin
Event|Event|Hospital Course|7034,7042|false|false|false|||remained
Event|Event|Hospital Course|7043,7049|false|false|false|||stable
Finding|Intellectual Product|Hospital Course|7043,7049|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|Hospital Course|7085,7093|false|false|false|||bleeding
Finding|Pathologic Function|Hospital Course|7085,7093|true|false|false|C0019080|Hemorrhage|bleeding
Event|Event|Hospital Course|7103,7108|false|false|false|||stool
Finding|Body Substance|Hospital Course|7103,7108|false|false|false|C0015733|Feces|stool
Event|Event|Hospital Course|7113,7118|false|false|false|||guiac
Event|Event|Hospital Course|7120,7128|false|false|false|||negative
Finding|Classification|Hospital Course|7120,7128|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|7120,7128|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|7120,7128|false|false|false|C5237010|Expression Negative|negative
Event|Event|Hospital Course|7136,7147|false|false|false|||transfusion
Finding|Functional Concept|Hospital Course|7136,7147|false|false|false|C0199960||transfusion
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7136,7147|false|false|false|C0005841;C1879316|Blood Transfusion;Transfusion (procedure)|transfusion
Finding|Body Substance|Hospital Course|7152,7159|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|7152,7159|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|7152,7159|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|7160,7168|false|false|false|||reported
Event|Event|Hospital Course|7169,7180|false|false|false|||significant
Finding|Idea or Concept|Hospital Course|7169,7180|false|false|false|C0750502|Significant|significant
Event|Event|Hospital Course|7182,7193|false|false|false|||improvement
Finding|Conceptual Entity|Hospital Course|7182,7193|false|false|false|C2986411|Improvement|improvement
Event|Event|Hospital Course|7201,7210|false|false|false|||shortness
Attribute|Clinical Attribute|Hospital Course|7201,7220|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|Hospital Course|7201,7220|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|Hospital Course|7214,7220|false|false|false|C0225386|Breath|breath
Event|Event|Hospital Course|7225,7232|false|false|false|||fatigue
Finding|Sign or Symptom|Hospital Course|7225,7232|false|false|false|C0015672|Fatigue|fatigue
Event|Event|Hospital Course|7245,7252|false|false|false|||history
Finding|Conceptual Entity|Hospital Course|7245,7252|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|7245,7252|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|7245,7252|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|7245,7255|false|false|false|C0262926|Medical History|history of
Finding|Finding|Hospital Course|7245,7265|false|false|false|C4041078|History of gastritis|history of gastritis
Disorder|Disease or Syndrome|Hospital Course|7256,7265|false|false|false|C0017152|Gastritis|gastritis
Event|Event|Hospital Course|7256,7265|false|false|false|||gastritis
Disorder|Disease or Syndrome|Hospital Course|7270,7284|false|false|false|C1510475|Diverticulosis|diverticulosis
Event|Event|Hospital Course|7270,7284|false|false|false|||diverticulosis
Finding|Pathologic Function|Hospital Course|7288,7296|false|false|false|C0017181|Gastrointestinal Hemorrhage|GI bleed
Event|Event|Hospital Course|7291,7296|false|false|false|||bleed
Finding|Pathologic Function|Hospital Course|7291,7296|false|false|false|C0019080|Hemorrhage|bleed
Event|Event|Hospital Course|7301,7309|false|false|false|||believed
Event|Event|Hospital Course|7311,7322|false|false|false|||responsible
Finding|Finding|Hospital Course|7311,7322|false|false|false|C1273518|Responsible to (attribute)|responsible
Disorder|Disease or Syndrome|Hospital Course|7331,7337|false|false|false|C0002871|Anemia|anemia
Event|Event|Hospital Course|7331,7337|false|false|false|||anemia
Finding|Body Substance|Hospital Course|7339,7346|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|7339,7346|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|7339,7346|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|7362,7364|false|false|false|||an
Event|Event|Hospital Course|7366,7369|false|false|false|||EGD
Procedure|Diagnostic Procedure|Hospital Course|7366,7369|false|false|false|C0079304|Esophagogastroduodenoscopy|EGD
Event|Event|Hospital Course|7370,7381|false|false|false|||colonoscopy
Procedure|Diagnostic Procedure|Hospital Course|7370,7381|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Procedure|Health Care Activity|Hospital Course|7370,7381|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Event|Event|Hospital Course|7388,7398|false|false|false|||outpatient
Finding|Classification|Hospital Course|7388,7398|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|7388,7398|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Intellectual Product|Hospital Course|7404,7409|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Finding|Finding|Hospital Course|7404,7422|false|false|false|C0743630|exacerbation acute|Acute exacerbation
Event|Event|Hospital Course|7410,7422|false|false|false|||exacerbation
Finding|Finding|Hospital Course|7410,7422|false|false|false|C4086268|Exacerbation|exacerbation
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7426,7431|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Hospital Course|7426,7431|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Hospital Course|7426,7431|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|Hospital Course|7426,7439|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Event|Event|Hospital Course|7432,7439|false|false|false|||failure
Finding|Functional Concept|Hospital Course|7432,7439|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|Hospital Course|7432,7439|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|Hospital Course|7432,7439|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Attribute|Clinical Attribute|Hospital Course|7455,7463|false|false|false|C0812388|Ejection time|ejection
Event|Event|Hospital Course|7455,7463|false|false|false|||ejection
Finding|Daily or Recreational Activity|Hospital Course|7455,7463|false|false|false|C0336969|Ejection as a Sports activity|ejection
Phenomenon|Phenomenon or Process|Hospital Course|7455,7463|false|false|false|C0302131|Ejection as a Circumstance of Injury|ejection
Event|Event|Hospital Course|7465,7473|false|false|false|||fraction
Finding|Intellectual Product|Hospital Course|7465,7473|false|false|false|C1554103|MDFAttributeType - Fraction|fraction
Finding|Body Substance|Hospital Course|7480,7487|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|7480,7487|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|7480,7487|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|7497,7502|false|false|false|||found
Event|Event|Hospital Course|7518,7524|false|false|false|||volume
Finding|Intellectual Product|Hospital Course|7518,7524|false|false|false|C1705102|Volume (publication)|volume
Event|Event|Hospital Course|7546,7553|false|false|false|||treated
Event|Event|Hospital Course|7559,7565|false|false|false|||2x40mg
Drug|Organic Chemical|Hospital Course|7569,7574|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|Hospital Course|7569,7574|false|false|false|C0699992|Lasix|Lasix
Event|Event|Hospital Course|7569,7574|false|false|false|||Lasix
Finding|Idea or Concept|Hospital Course|7581,7585|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Finding|Body Substance|Hospital Course|7586,7591|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|Hospital Course|7586,7591|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|Hospital Course|7586,7591|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Attribute|Clinical Attribute|Hospital Course|7586,7598|false|false|false|C0232856;C0489132||urine output
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7586,7598|false|false|false|C2094175|monitoring of urine output for fluid balance|urine output
Event|Event|Hospital Course|7592,7598|false|false|false|||output
Finding|Conceptual Entity|Hospital Course|7592,7598|false|false|false|C1709366|system output|output
Procedure|Health Care Activity|Hospital Course|7592,7598|false|false|false|C3251815|Measurement of fluid output|output
Finding|Functional Concept|Hospital Course|7604,7615|false|false|false|C0231220|Symptomatic|symptomatic
Event|Event|Hospital Course|7616,7627|false|false|false|||improvement
Finding|Conceptual Entity|Hospital Course|7616,7627|false|false|false|C2986411|Improvement|improvement
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7633,7642|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Hospital Course|7633,7642|false|false|false|C2707265||pulmonary
Finding|Finding|Hospital Course|7633,7642|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|Hospital Course|7633,7648|false|false|false|C0034063|Pulmonary Edema|pulmonary edema
Attribute|Clinical Attribute|Hospital Course|7643,7648|false|false|false|C1717255||edema
Event|Event|Hospital Course|7643,7648|false|false|false|||edema
Finding|Pathologic Function|Hospital Course|7643,7648|false|false|false|C0013604|Edema|edema
Attribute|Clinical Attribute|Hospital Course|7665,7670|false|false|false|C1717255||edema
Event|Event|Hospital Course|7665,7670|false|false|false|||edema
Finding|Pathologic Function|Hospital Course|7665,7670|false|false|false|C0013604|Edema|edema
Event|Event|Hospital Course|7671,7679|false|false|false|||resolved
Event|Event|Hospital Course|7685,7693|false|false|false|||diuresis
Finding|Organ or Tissue Function|Hospital Course|7685,7693|false|false|false|C0012797|Diuresis|diuresis
Event|Event|Hospital Course|7696,7703|false|false|false|||CHRONIC
Finding|Intellectual Product|Hospital Course|7696,7703|false|false|false|C1547296|Chronic - Admission Level of Care Code|CHRONIC
Procedure|Health Care Activity|Hospital Course|7696,7703|false|false|false|C1555457|Provision of recurring care for chronic illness|CHRONIC
Event|Event|Hospital Course|7721,7731|false|false|false|||ulceration
Finding|Pathologic Function|Hospital Course|7721,7731|false|false|false|C0041582;C3887532|Ulcer;Ulceration|ulceration
Event|Event|Hospital Course|7734,7743|false|false|false|||Continued
Finding|Idea or Concept|Hospital Course|7747,7751|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|7747,7751|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|7747,7751|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|7752,7764|false|false|false|C0081876|pantoprazole|pantoprazole
Drug|Pharmacologic Substance|Hospital Course|7752,7764|false|false|false|C0081876|pantoprazole|pantoprazole
Event|Event|Hospital Course|7752,7764|false|false|false|||pantoprazole
Disorder|Mental or Behavioral Dysfunction|Hospital Course|7765,7768|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7765,7768|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|7765,7768|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|7765,7768|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|7765,7768|false|false|false|C1332410|BID gene|BID
Disorder|Disease or Syndrome|Hospital Course|7772,7784|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|Hospital Course|7772,7784|false|false|false|||Hypertension
Event|Event|Hospital Course|7786,7795|false|false|false|||Continued
Finding|Idea or Concept|Hospital Course|7799,7803|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|7799,7803|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|7799,7803|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|7804,7814|false|false|false|C0028066|nifedipine|nifedipine
Drug|Pharmacologic Substance|Hospital Course|7804,7814|false|false|false|C0028066|nifedipine|nifedipine
Event|Event|Hospital Course|7804,7814|false|false|false|||nifedipine
Event|Event|Hospital Course|7816,7826|false|false|false|||carvadilol
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7828,7838|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|Hospital Course|7828,7838|false|false|false|C0065374|lisinopril|lisinopril
Event|Event|Hospital Course|7828,7838|false|false|false|||lisinopril
Attribute|Clinical Attribute|Hospital Course|7843,7848|false|false|false|C1300072|Tumor stage|Stage
Finding|Intellectual Product|Hospital Course|7843,7851|false|false|false|C0441772|Stage level 4|Stage IV
Finding|Intellectual Product|Hospital Course|7852,7859|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|Hospital Course|7852,7859|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Disorder|Disease or Syndrome|Hospital Course|7852,7874|false|false|false|C1561643|Chronic Kidney Diseases|Chronic Kidney Disease
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7860,7866|false|false|false|C0022646;C0227665|Both kidneys;Kidney|Kidney
Disorder|Neoplastic Process|Hospital Course|7860,7866|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|Kidney
Finding|Sign or Symptom|Hospital Course|7860,7866|false|false|false|C0812426|Kidney problem|Kidney
Procedure|Diagnostic Procedure|Hospital Course|7860,7866|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|Kidney
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7860,7866|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|Kidney
Disorder|Disease or Syndrome|Hospital Course|7860,7874|false|false|false|C0022658|Kidney Diseases|Kidney Disease
Disorder|Disease or Syndrome|Hospital Course|7867,7874|false|false|false|C0012634|Disease|Disease
Event|Event|Hospital Course|7867,7874|false|false|false|||Disease
Drug|Biologically Active Substance|Hospital Course|7877,7887|false|false|false|C0010294|creatinine|Creatinine
Drug|Organic Chemical|Hospital Course|7877,7887|false|false|false|C0010294|creatinine|Creatinine
Event|Event|Hospital Course|7877,7887|false|false|false|||Creatinine
Finding|Physiologic Function|Hospital Course|7877,7887|false|false|false|C4551889|Creatinine metabolic function|Creatinine
Procedure|Laboratory Procedure|Hospital Course|7877,7887|false|false|false|C0201975|Creatinine measurement|Creatinine
Event|Event|Hospital Course|7888,7896|false|false|false|||remained
Drug|Biomedical or Dental Material|Hospital Course|7900,7908|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|Hospital Course|7900,7908|false|false|false|||baseline
Finding|Idea or Concept|Hospital Course|7900,7908|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|Hospital Course|7934,7943|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|7934,7943|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Idea or Concept|Hospital Course|7946,7958|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Finding|Body Substance|Hospital Course|7991,7998|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|7991,7998|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|7991,7998|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Disorder|Disease or Syndrome|Hospital Course|8001,8007|false|false|false|C0002871|Anemia|Anemia
Event|Event|Hospital Course|8001,8007|false|false|false|||Anemia
Event|Event|Hospital Course|8011,8018|false|false|false|||thought
Finding|Pathologic Function|Hospital Course|8037,8045|false|false|false|C0017181|Gastrointestinal Hemorrhage|GI bleed
Finding|Pathologic Function|Hospital Course|8040,8045|false|false|false|C0019080|Hemorrhage|bleed
Event|Event|Hospital Course|8053,8060|false|false|false|||history
Finding|Conceptual Entity|Hospital Course|8053,8060|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|8053,8060|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|8053,8060|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|8053,8063|false|false|false|C0262926|Medical History|history of
Finding|Finding|Hospital Course|8053,8073|false|false|false|C4041078|History of gastritis|history of gastritis
Disorder|Disease or Syndrome|Hospital Course|8064,8073|false|false|false|C0017152|Gastritis|gastritis
Event|Event|Hospital Course|8064,8073|false|false|false|||gastritis
Disorder|Disease or Syndrome|Hospital Course|8078,8092|false|false|false|C1510475|Diverticulosis|diverticulosis
Event|Event|Hospital Course|8078,8092|false|false|false|||diverticulosis
Event|Event|Hospital Course|8101,8109|false|false|false|||schedule
Finding|Intellectual Product|Hospital Course|8101,8109|false|false|false|C0086960|Schedule (document)|schedule
Procedure|Health Care Activity|Hospital Course|8101,8109|false|false|false|C1446911|Scheduling (procedure)|schedule
Event|Event|Hospital Course|8111,8114|false|false|false|||EGD
Procedure|Diagnostic Procedure|Hospital Course|8111,8114|false|false|false|C0079304|Esophagogastroduodenoscopy|EGD
Event|Event|Hospital Course|8115,8126|false|false|false|||colonoscopy
Procedure|Diagnostic Procedure|Hospital Course|8115,8126|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Procedure|Health Care Activity|Hospital Course|8115,8126|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Finding|Idea or Concept|Hospital Course|8138,8142|false|false|false|C1552851|next - HtmlLinkType|next
Finding|Idea or Concept|Hospital Course|8143,8148|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|Hospital Course|8143,8148|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Body Substance|Hospital Course|8151,8158|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|8151,8158|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|8151,8158|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|8159,8168|false|false|false|||continued
Drug|Organic Chemical|Hospital Course|8172,8180|false|false|false|C0699129|Coumadin|Coumadin
Drug|Pharmacologic Substance|Hospital Course|8172,8180|false|false|false|C0699129|Coumadin|Coumadin
Event|Event|Hospital Course|8172,8180|false|false|false|||Coumadin
Disorder|Disease or Syndrome|Hospital Course|8195,8199|false|false|false|C0151950|Deep thrombophlebitis|DVTs
Event|Event|Hospital Course|8195,8199|false|false|false|||DVTs
Event|Event|Hospital Course|8209,8217|false|false|false|||continue
Event|Event|Hospital Course|8221,8226|false|false|false|||weigh
Event|Event|Hospital Course|8231,8236|false|false|false|||risks
Finding|Idea or Concept|Hospital Course|8231,8236|false|false|false|C0035647|Risk|risks
Event|Event|Hospital Course|8241,8249|false|false|false|||benefits
Event|Event|Hospital Course|8253,8268|false|false|false|||anticoagulation
Finding|Finding|Hospital Course|8253,8268|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|Hospital Course|8253,8268|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8253,8268|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Event|Event|Hospital Course|8276,8283|false|false|false|||history
Finding|Conceptual Entity|Hospital Course|8276,8283|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|8276,8283|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|8276,8283|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|8276,8286|false|false|false|C0262926|Medical History|history of
Event|Event|Hospital Course|8287,8292|false|false|false|||bleed
Finding|Pathologic Function|Hospital Course|8287,8292|false|false|false|C0019080|Hemorrhage|bleed
Event|Event|Hospital Course|8296,8305|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|8296,8305|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|8296,8305|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|8296,8305|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|8296,8305|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|8306,8312|false|false|false|C0944911||weight
Event|Event|Hospital Course|8306,8312|false|false|false|||weight
Finding|Finding|Hospital Course|8306,8312|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|Hospital Course|8306,8312|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|Hospital Course|8306,8312|false|false|false|C1305866|Weighing patient|weight
Event|Activity|Hospital Course|8323,8330|false|false|false|C3812666|Personal Contact|CONTACT
Event|Event|Hospital Course|8323,8330|false|false|false|||CONTACT
Finding|Functional Concept|Hospital Course|8323,8330|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Idea or Concept|Hospital Course|8323,8330|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Intellectual Product|Hospital Course|8323,8330|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Phenomenon|Phenomenon or Process|Hospital Course|8323,8330|false|false|false|C0392367|Physical contact|CONTACT
Event|Event|Hospital Course|8342,8346|false|false|false|||CODE
Event|Occupational Activity|Hospital Course|8342,8346|false|false|false|C0009219|Coding|CODE
Finding|Intellectual Product|Hospital Course|8342,8346|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|CODE
Event|Event|Hospital Course|8354,8363|false|false|false|||confirmed
Attribute|Clinical Attribute|Hospital Course|8366,8377|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|8366,8377|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|8366,8377|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|8366,8377|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|8366,8390|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|8381,8390|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|8381,8390|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|Hospital Course|8409,8419|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Hospital Course|8409,8419|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|Hospital Course|8409,8424|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|Hospital Course|8420,8424|false|false|false|||list
Finding|Intellectual Product|Hospital Course|8420,8424|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|Hospital Course|8432,8442|false|false|false|||inaccurate
Event|Event|Hospital Course|8447,8455|false|false|false|||requires
Event|Event|Hospital Course|8464,8477|false|false|false|||investigation
Finding|Intellectual Product|Hospital Course|8464,8477|false|false|false|C1552578|Act Class - investigation|investigation
Procedure|Health Care Activity|Hospital Course|8464,8477|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|investigation
Drug|Organic Chemical|Hospital Course|8482,8493|false|false|false|C0002144|allopurinol|Allopurinol
Drug|Pharmacologic Substance|Hospital Course|8482,8493|false|false|false|C0002144|allopurinol|Allopurinol
Event|Event|Hospital Course|8516,8519|false|false|false|||DAY
Finding|Idea or Concept|Hospital Course|8516,8519|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|DAY
Finding|Intellectual Product|Hospital Course|8516,8519|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|DAY
Drug|Organic Chemical|Hospital Course|8524,8531|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Hospital Course|8524,8531|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|Hospital Course|8551,8563|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|8551,8563|false|false|false|C0286651|atorvastatin|Atorvastatin
Event|Event|Hospital Course|8573,8576|false|false|false|||QPM
Drug|Organic Chemical|Hospital Course|8581,8591|false|false|false|C0054836|carvedilol|Carvedilol
Drug|Pharmacologic Substance|Hospital Course|8581,8591|false|false|false|C0054836|carvedilol|Carvedilol
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8603,8606|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8603,8606|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8603,8606|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|8603,8606|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|8603,8606|false|false|false|C1332410|BID gene|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8611,8621|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|Hospital Course|8611,8621|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Organic Chemical|Hospital Course|8641,8654|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|Hospital Course|8641,8654|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|Hospital Course|8641,8654|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Event|Event|Hospital Course|8641,8654|false|false|false|||Multivitamins
Drug|Biomedical or Dental Material|Hospital Course|8657,8660|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|Hospital Course|8657,8660|false|false|false|||TAB
Drug|Organic Chemical|Hospital Course|8674,8684|false|false|false|C0028066|nifedipine|NIFEdipine
Drug|Pharmacologic Substance|Hospital Course|8674,8684|false|false|false|C0028066|nifedipine|NIFEdipine
Event|Event|Hospital Course|8674,8684|false|false|false|||NIFEdipine
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8697,8700|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8697,8700|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8697,8700|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|8697,8700|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|8697,8700|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|8705,8712|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|8705,8712|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|8705,8712|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|Hospital Course|8705,8714|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|Hospital Course|8705,8714|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|Hospital Course|8705,8714|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|Hospital Course|8705,8714|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|Hospital Course|8705,8714|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|Hospital Course|8713,8714|false|false|false|||D
Event|Event|Hospital Course|8719,8723|false|false|false|||UNIT
Drug|Organic Chemical|Hospital Course|8737,8745|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|8737,8745|false|false|false|C1692318|docusate|Docusate
Event|Event|Hospital Course|8737,8745|false|false|false|||Docusate
Drug|Organic Chemical|Hospital Course|8737,8752|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|Hospital Course|8737,8752|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|Hospital Course|8746,8752|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|8746,8752|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|8746,8752|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|8746,8752|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|8746,8752|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|8746,8752|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8763,8766|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8763,8766|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8763,8766|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|8763,8766|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|8763,8766|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|8772,8782|false|false|false|C0060926|gabapentin|Gabapentin
Drug|Pharmacologic Substance|Hospital Course|8772,8782|false|false|false|C0060926|gabapentin|Gabapentin
Finding|Finding|Hospital Course|8797,8813|false|false|false|C0027796;C3714625|Neuralgia;Neuropathic pain|neuropathic pain
Finding|Sign or Symptom|Hospital Course|8797,8813|false|false|false|C0027796;C3714625|Neuralgia;Neuropathic pain|neuropathic pain
Attribute|Clinical Attribute|Hospital Course|8809,8813|false|false|false|C2598155||pain
Event|Event|Hospital Course|8809,8813|false|false|false|||pain
Finding|Functional Concept|Hospital Course|8809,8813|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|8809,8813|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|8819,8831|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Pharmacologic Substance|Hospital Course|8819,8831|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Organic Chemical|Hospital Course|8851,8856|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|Hospital Course|8851,8856|false|false|false|C3489575|sennosides, USP|Senna
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8867,8870|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8867,8870|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8867,8870|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|8867,8870|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|8867,8870|false|false|false|C1332410|BID gene|BID
Event|Event|Hospital Course|8871,8883|false|false|false|||constipation
Finding|Sign or Symptom|Hospital Course|8871,8883|false|false|false|C0009806|Constipation|constipation
Drug|Hazardous or Poisonous Substance|Hospital Course|8889,8897|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|Hospital Course|8889,8897|false|false|false|C0043031|warfarin|Warfarin
Drug|Pharmacologic Substance|Hospital Course|8889,8897|false|false|false|C0043031|warfarin|Warfarin
Finding|Intellectual Product|Hospital Course|8909,8913|false|false|false|C1561540|Transaction counts and value totals - week|WEEK
Drug|Organic Chemical|Hospital Course|8925,8938|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Pharmacologic Substance|Hospital Course|8925,8938|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Event|Event|Hospital Course|8925,8938|false|false|false|||Nitroglycerin
Finding|Gene or Genome|Hospital Course|8958,8961|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Location or Region|Hospital Course|8962,8967|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|8962,8967|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|8962,8972|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Hospital Course|8962,8972|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Hospital Course|8968,8972|false|true|false|C2598155||pain
Event|Event|Hospital Course|8968,8972|false|false|false|||pain
Finding|Functional Concept|Hospital Course|8968,8972|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|8968,8972|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|8978,8988|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|Hospital Course|8978,8988|false|false|false|C0016860|furosemide|Furosemide
Drug|Biomedical or Dental Material|Hospital Course|9009,9021|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Drug|Organic Chemical|Hospital Course|9009,9021|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Event|Event|Hospital Course|9009,9021|false|false|false|||Polyethylene
Drug|Organic Chemical|Hospital Course|9009,9028|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Pharmacologic Substance|Hospital Course|9009,9028|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Hazardous or Poisonous Substance|Hospital Course|9022,9028|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Drug|Organic Chemical|Hospital Course|9022,9028|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Drug|Organic Chemical|Hospital Course|9048,9061|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|9048,9061|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Hospital Course|9048,9061|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|9048,9061|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|Hospital Course|9080,9083|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|9084,9088|false|false|false|C2598155||pain
Event|Event|Hospital Course|9084,9088|false|false|false|||pain
Finding|Functional Concept|Hospital Course|9084,9088|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|9084,9088|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|9092,9097|false|false|false|||fever
Finding|Finding|Hospital Course|9092,9097|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|Hospital Course|9092,9097|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Drug|Hazardous or Poisonous Substance|Hospital Course|9103,9111|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|Hospital Course|9103,9111|false|false|false|C0043031|warfarin|Warfarin
Drug|Pharmacologic Substance|Hospital Course|9103,9111|false|false|false|C0043031|warfarin|Warfarin
Finding|Intellectual Product|Hospital Course|9123,9127|false|false|false|C1561540|Transaction counts and value totals - week|WEEK
Event|Event|Hospital Course|9154,9160|false|false|false|||Dinner
Finding|Daily or Recreational Activity|Hospital Course|9154,9160|false|false|false|C4048877|Dinner|Dinner
Event|Event|Hospital Course|9164,9173|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|9164,9173|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|9164,9173|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|9164,9173|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|9164,9173|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|9164,9185|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|9174,9185|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|9174,9185|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|9174,9185|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|9174,9185|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|9190,9203|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|9190,9203|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Hospital Course|9190,9203|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|9190,9203|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|Hospital Course|9222,9225|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|9226,9230|false|false|false|C2598155||pain
Event|Event|Hospital Course|9226,9230|false|false|false|||pain
Finding|Functional Concept|Hospital Course|9226,9230|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|9226,9230|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|9234,9239|false|false|false|||fever
Finding|Finding|Hospital Course|9234,9239|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|Hospital Course|9234,9239|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Drug|Organic Chemical|Hospital Course|9245,9258|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Drug|Pharmacologic Substance|Hospital Course|9245,9258|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Event|Event|Hospital Course|9245,9258|false|false|false|||acetaminophen
Procedure|Laboratory Procedure|Hospital Course|9245,9258|false|false|false|C0373527|Acetaminophen measurement|acetaminophen
Drug|Biomedical or Dental Material|Hospital Course|9270,9276|false|false|false|C0039225|Tablet Dosage Form|tablet
Event|Event|Hospital Course|9270,9276|false|false|false|||tablet
Finding|Functional Concept|Hospital Course|9280,9288|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|9283,9288|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|9283,9288|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Gene or Genome|Hospital Course|9293,9296|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|9297,9301|false|false|false|||Disp
Drug|Biomedical or Dental Material|Hospital Course|9309,9315|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|9316,9323|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|9316,9323|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|9330,9337|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Hospital Course|9330,9337|false|false|false|C0004057|aspirin|Aspirin
Event|Event|Hospital Course|9354,9356|false|false|false|||RX
Drug|Organic Chemical|Hospital Course|9358,9365|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|Hospital Course|9358,9365|false|false|false|C0004057|aspirin|aspirin
Event|Event|Hospital Course|9358,9365|false|false|false|||aspirin
Drug|Biomedical or Dental Material|Hospital Course|9374,9380|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|9384,9392|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|9387,9392|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|9387,9392|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Biomedical or Dental Material|Hospital Course|9409,9415|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|9409,9415|false|false|false|||Tablet
Event|Event|Hospital Course|9417,9424|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|9417,9424|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|9431,9443|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|9431,9443|false|false|false|C0286651|atorvastatin|Atorvastatin
Event|Event|Hospital Course|9453,9456|false|false|false|||QPM
Drug|Organic Chemical|Hospital Course|9462,9474|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|Hospital Course|9462,9474|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|Hospital Course|9462,9474|false|false|false|||atorvastatin
Drug|Biomedical or Dental Material|Hospital Course|9483,9489|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|9493,9501|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|9496,9501|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|9496,9501|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Event|Hospital Course|9502,9505|false|false|false|||QPM
Drug|Biomedical or Dental Material|Hospital Course|9516,9522|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|9516,9522|false|false|false|||Tablet
Event|Event|Hospital Course|9524,9531|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|9524,9531|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|9538,9548|false|false|false|C0054836|carvedilol|Carvedilol
Drug|Pharmacologic Substance|Hospital Course|9538,9548|false|false|false|C0054836|carvedilol|Carvedilol
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9560,9563|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9560,9563|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9560,9563|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|9560,9563|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|9560,9563|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|9569,9579|false|false|false|C0054836|carvedilol|carvedilol
Drug|Pharmacologic Substance|Hospital Course|9569,9579|false|false|false|C0054836|carvedilol|carvedilol
Event|Event|Hospital Course|9569,9579|false|false|false|||carvedilol
Drug|Biomedical or Dental Material|Hospital Course|9590,9596|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|9600,9608|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|9603,9608|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|9603,9608|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|Hospital Course|9617,9620|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|9617,9620|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Activity|Hospital Course|9621,9625|false|false|false|C1880359|Dispense (activity)|Disp
Finding|Gene or Genome|Hospital Course|9621,9625|false|false|false|C2828567|PRSS30P gene|Disp
Drug|Biomedical or Dental Material|Hospital Course|9632,9638|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|9639,9646|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|9639,9646|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|9653,9661|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|9653,9661|false|false|false|C1692318|docusate|Docusate
Event|Event|Hospital Course|9653,9661|false|false|false|||Docusate
Drug|Organic Chemical|Hospital Course|9653,9668|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|Hospital Course|9653,9668|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|Hospital Course|9662,9668|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|9662,9668|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|9662,9668|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|9662,9668|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|9662,9668|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|9662,9668|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9679,9682|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9679,9682|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9679,9682|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|9679,9682|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|9679,9682|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|9688,9696|false|false|false|C1692318|docusate|docusate
Drug|Pharmacologic Substance|Hospital Course|9688,9696|false|false|false|C1692318|docusate|docusate
Drug|Organic Chemical|Hospital Course|9688,9703|false|false|false|C0243237|docusate sodium|docusate sodium
Drug|Pharmacologic Substance|Hospital Course|9688,9703|false|false|false|C0243237|docusate sodium|docusate sodium
Drug|Biologically Active Substance|Hospital Course|9697,9703|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|Hospital Course|9697,9703|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|Hospital Course|9697,9703|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Event|Event|Hospital Course|9697,9703|false|false|false|||sodium
Finding|Physiologic Function|Hospital Course|9697,9703|false|false|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|Hospital Course|9697,9703|false|false|false|C0337443|Sodium measurement|sodium
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9713,9720|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|Hospital Course|9713,9720|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|Hospital Course|9713,9720|false|false|false|C0006935|capsule (pharmacologic)|capsule
Finding|Functional Concept|Hospital Course|9724,9732|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|9727,9732|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|9727,9732|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|Hospital Course|9741,9744|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|9741,9744|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9756,9763|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|9756,9763|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|9756,9763|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Event|Event|Hospital Course|9764,9771|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|9764,9771|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|9778,9788|false|false|false|C0060926|gabapentin|Gabapentin
Drug|Pharmacologic Substance|Hospital Course|9778,9788|false|false|false|C0060926|gabapentin|Gabapentin
Finding|Finding|Hospital Course|9803,9819|false|false|false|C0027796;C3714625|Neuralgia;Neuropathic pain|neuropathic pain
Finding|Sign or Symptom|Hospital Course|9803,9819|false|false|false|C0027796;C3714625|Neuralgia;Neuropathic pain|neuropathic pain
Attribute|Clinical Attribute|Hospital Course|9815,9819|false|false|false|C2598155||pain
Event|Event|Hospital Course|9815,9819|false|false|false|||pain
Finding|Functional Concept|Hospital Course|9815,9819|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|9815,9819|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|9825,9835|false|false|false|C0060926|gabapentin|gabapentin
Drug|Pharmacologic Substance|Hospital Course|9825,9835|false|false|false|C0060926|gabapentin|gabapentin
Event|Event|Hospital Course|9825,9835|false|false|false|||gabapentin
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9845,9852|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|Hospital Course|9845,9852|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|Hospital Course|9845,9852|false|false|false|C0006935|capsule (pharmacologic)|capsule
Finding|Functional Concept|Hospital Course|9856,9864|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|9859,9864|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|9859,9864|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9887,9894|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|9887,9894|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|9887,9894|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Event|Event|Hospital Course|9895,9902|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|9895,9902|false|false|false|C0807726|refill|Refills
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9909,9919|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|Hospital Course|9909,9919|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9940,9950|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|Hospital Course|9940,9950|false|false|false|C0065374|lisinopril|lisinopril
Event|Event|Hospital Course|9940,9950|false|false|false|||lisinopril
Drug|Biomedical or Dental Material|Hospital Course|9959,9965|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|9969,9977|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|9972,9977|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|9972,9977|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Biomedical or Dental Material|Hospital Course|9994,10000|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|9994,10000|false|false|false|||Tablet
Event|Event|Hospital Course|10002,10009|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|10002,10009|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|10016,10029|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|Hospital Course|10016,10029|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|Hospital Course|10016,10029|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Event|Event|Hospital Course|10016,10029|false|false|false|||Multivitamins
Drug|Biomedical or Dental Material|Hospital Course|10032,10035|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|Hospital Course|10032,10035|false|false|false|||TAB
Event|Event|Hospital Course|10046,10048|false|false|false|||RX
Drug|Organic Chemical|Hospital Course|10050,10062|false|false|false|C0301532|Multivitamin preparation|multivitamin
Drug|Pharmacologic Substance|Hospital Course|10050,10062|false|false|false|C0301532|Multivitamin preparation|multivitamin
Drug|Vitamin|Hospital Course|10050,10062|false|false|false|C0301532|Multivitamin preparation|multivitamin
Event|Event|Hospital Course|10050,10062|false|false|false|||multivitamin
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10066,10073|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|Hospital Course|10066,10073|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|Hospital Course|10066,10073|false|false|false|C0006935|capsule (pharmacologic)|capsule
Finding|Functional Concept|Hospital Course|10077,10085|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|10080,10085|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|10080,10085|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10102,10109|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|10102,10109|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|10102,10109|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Event|Event|Hospital Course|10111,10118|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|10111,10118|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|10125,10135|false|false|false|C0028066|nifedipine|NIFEdipine
Drug|Pharmacologic Substance|Hospital Course|10125,10135|false|false|false|C0028066|nifedipine|NIFEdipine
Event|Event|Hospital Course|10125,10135|false|false|false|||NIFEdipine
Disorder|Mental or Behavioral Dysfunction|Hospital Course|10148,10151|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10148,10151|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|10148,10151|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|10148,10151|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|10148,10151|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|10157,10167|false|false|false|C0028066|nifedipine|nifedipine
Drug|Pharmacologic Substance|Hospital Course|10157,10167|false|false|false|C0028066|nifedipine|nifedipine
Event|Event|Hospital Course|10157,10167|false|false|false|||nifedipine
Drug|Biomedical or Dental Material|Hospital Course|10176,10182|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|10186,10194|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|10189,10194|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|10189,10194|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|Hospital Course|10203,10206|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|10203,10206|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biomedical or Dental Material|Hospital Course|10218,10224|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|10225,10232|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|10225,10232|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|10240,10253|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Pharmacologic Substance|Hospital Course|10240,10253|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Event|Event|Hospital Course|10240,10253|false|false|false|||Nitroglycerin
Finding|Gene or Genome|Hospital Course|10273,10276|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Location or Region|Hospital Course|10277,10282|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|10277,10282|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|10277,10287|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Hospital Course|10277,10287|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Hospital Course|10283,10287|false|true|false|C2598155||pain
Event|Event|Hospital Course|10283,10287|false|false|false|||pain
Finding|Functional Concept|Hospital Course|10283,10287|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|10283,10287|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|10289,10291|false|false|false|||RX
Drug|Organic Chemical|Hospital Course|10293,10306|false|false|false|C0017887|nitroglycerin|nitroglycerin
Drug|Pharmacologic Substance|Hospital Course|10293,10306|false|false|false|C0017887|nitroglycerin|nitroglycerin
Event|Event|Hospital Course|10293,10306|false|false|false|||nitroglycerin
Drug|Organic Chemical|Hospital Course|10308,10317|false|false|false|C0699241|Nitrostat|Nitrostat
Drug|Pharmacologic Substance|Hospital Course|10308,10317|false|false|false|C0699241|Nitrostat|Nitrostat
Drug|Biomedical or Dental Material|Hospital Course|10328,10334|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Gene or Genome|Hospital Course|10358,10361|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Biomedical or Dental Material|Hospital Course|10372,10378|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|10379,10386|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|10379,10386|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|10394,10406|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Pharmacologic Substance|Hospital Course|10394,10406|false|false|false|C0081876|pantoprazole|Pantoprazole
Event|Event|Hospital Course|10422,10424|false|false|false|||RX
Drug|Organic Chemical|Hospital Course|10426,10438|false|false|false|C0081876|pantoprazole|pantoprazole
Drug|Pharmacologic Substance|Hospital Course|10426,10438|false|false|false|C0081876|pantoprazole|pantoprazole
Event|Event|Hospital Course|10426,10438|false|false|false|||pantoprazole
Drug|Biomedical or Dental Material|Hospital Course|10447,10453|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|10457,10465|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|10460,10465|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|10460,10465|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Biomedical or Dental Material|Hospital Course|10501,10507|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|10508,10515|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|10508,10515|false|false|false|C0807726|refill|Refills
Drug|Biomedical or Dental Material|Hospital Course|10523,10535|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Drug|Organic Chemical|Hospital Course|10523,10535|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Event|Event|Hospital Course|10523,10535|false|false|false|||Polyethylene
Drug|Organic Chemical|Hospital Course|10523,10542|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Pharmacologic Substance|Hospital Course|10523,10542|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Hazardous or Poisonous Substance|Hospital Course|10536,10542|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Drug|Organic Chemical|Hospital Course|10536,10542|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Event|Event|Hospital Course|10536,10542|false|false|false|||Glycol
Drug|Biomedical or Dental Material|Hospital Course|10562,10574|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|polyethylene
Drug|Organic Chemical|Hospital Course|10562,10574|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|polyethylene
Drug|Organic Chemical|Hospital Course|10562,10581|false|false|false|C0032483|polyethylene glycols|polyethylene glycol
Drug|Pharmacologic Substance|Hospital Course|10562,10581|false|false|false|C0032483|polyethylene glycols|polyethylene glycol
Drug|Organic Chemical|Hospital Course|10562,10586|false|false|false|C0724672|polyethylene glycol 3350|polyethylene glycol 3350
Drug|Pharmacologic Substance|Hospital Course|10562,10586|false|false|false|C0724672|polyethylene glycol 3350|polyethylene glycol 3350
Drug|Hazardous or Poisonous Substance|Hospital Course|10575,10581|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|glycol
Drug|Organic Chemical|Hospital Course|10575,10581|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|glycol
Event|Event|Hospital Course|10575,10581|false|false|false|||glycol
Drug|Biomedical or Dental Material|Hospital Course|10602,10608|false|false|false|C0032861;C1382110|Powder dose form;powder physical state|powder
Drug|Substance|Hospital Course|10602,10608|false|false|false|C0032861;C1382110|Powder dose form;powder physical state|powder
Event|Event|Hospital Course|10602,10608|false|false|false|||powder
Finding|Functional Concept|Hospital Course|10612,10620|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|10615,10620|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|10615,10620|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Event|Hospital Course|10628,10635|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|10628,10635|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|10643,10648|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|Hospital Course|10643,10648|false|false|false|C3489575|sennosides, USP|Senna
Disorder|Mental or Behavioral Dysfunction|Hospital Course|10659,10662|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10659,10662|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|10659,10662|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|10659,10662|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|10659,10662|false|false|false|C1332410|BID gene|BID
Event|Event|Hospital Course|10663,10675|false|false|false|||constipation
Finding|Sign or Symptom|Hospital Course|10663,10675|false|false|false|C0009806|Constipation|constipation
Drug|Organic Chemical|Hospital Course|10681,10691|false|false|false|C3489575|sennosides, USP|sennosides
Drug|Pharmacologic Substance|Hospital Course|10681,10691|false|false|false|C3489575|sennosides, USP|sennosides
Drug|Organic Chemical|Hospital Course|10693,10698|false|false|false|C3489575|sennosides, USP|senna
Drug|Pharmacologic Substance|Hospital Course|10693,10698|false|false|false|C3489575|sennosides, USP|senna
Event|Event|Hospital Course|10693,10698|false|false|false|||senna
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10709,10716|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|Hospital Course|10709,10716|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|Hospital Course|10709,10716|false|false|false|C0006935|capsule (pharmacologic)|capsule
Finding|Functional Concept|Hospital Course|10717,10725|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|10720,10725|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|10720,10725|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|Hospital Course|10734,10737|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|10734,10737|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10749,10756|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|10749,10756|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|10749,10756|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Event|Event|Hospital Course|10757,10764|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|10757,10764|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|10772,10779|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|10772,10779|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|10772,10779|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|Hospital Course|10772,10781|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|Hospital Course|10772,10781|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|Hospital Course|10772,10781|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|Hospital Course|10772,10781|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|Hospital Course|10772,10781|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|Hospital Course|10780,10781|false|false|false|||D
Event|Event|Hospital Course|10786,10790|false|false|false|||UNIT
Event|Event|Hospital Course|10801,10803|false|false|false|||RX
Drug|Organic Chemical|Hospital Course|10805,10819|false|false|false|C0014695;C3714696|Ergocalciferol Drug Product;ergocalciferol|ergocalciferol
Drug|Pharmacologic Substance|Hospital Course|10805,10819|false|false|false|C0014695;C3714696|Ergocalciferol Drug Product;ergocalciferol|ergocalciferol
Drug|Vitamin|Hospital Course|10805,10819|false|false|false|C0014695;C3714696|Ergocalciferol Drug Product;ergocalciferol|ergocalciferol
Event|Event|Hospital Course|10805,10819|false|false|false|||ergocalciferol
Drug|Organic Chemical|Hospital Course|10805,10832|false|false|false|C0014695|ergocalciferol|ergocalciferol (vitamin D2)
Drug|Pharmacologic Substance|Hospital Course|10805,10832|false|false|false|C0014695|ergocalciferol|ergocalciferol (vitamin D2)
Drug|Vitamin|Hospital Course|10805,10832|false|false|false|C0014695|ergocalciferol|ergocalciferol (vitamin D2)
Drug|Organic Chemical|Hospital Course|10821,10828|false|false|false|C0042890|Vitamins|vitamin
Drug|Pharmacologic Substance|Hospital Course|10821,10828|false|false|false|C0042890|Vitamins|vitamin
Drug|Vitamin|Hospital Course|10821,10828|false|false|false|C0042890|Vitamins|vitamin
Event|Event|Hospital Course|10821,10828|false|false|false|||vitamin
Drug|Organic Chemical|Hospital Course|10821,10831|false|false|false|C0014695|ergocalciferol|vitamin D2
Drug|Pharmacologic Substance|Hospital Course|10821,10831|false|false|false|C0014695|ergocalciferol|vitamin D2
Drug|Vitamin|Hospital Course|10821,10831|false|false|false|C0014695|ergocalciferol|vitamin D2
Drug|Biomedical or Dental Material|Hospital Course|10846,10852|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|10856,10864|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|10859,10864|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|10859,10864|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Biomedical or Dental Material|Hospital Course|10882,10888|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|10889,10896|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|10889,10896|false|false|false|C0807726|refill|Refills
Drug|Hazardous or Poisonous Substance|Hospital Course|10904,10912|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|Hospital Course|10904,10912|false|false|false|C0043031|warfarin|Warfarin
Drug|Pharmacologic Substance|Hospital Course|10904,10912|false|false|false|C0043031|warfarin|Warfarin
Finding|Intellectual Product|Hospital Course|10924,10928|false|false|false|C1561540|Transaction counts and value totals - week|WEEK
Drug|Hazardous or Poisonous Substance|Hospital Course|10940,10948|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|Hospital Course|10940,10948|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|Hospital Course|10940,10948|false|false|false|C0043031|warfarin|warfarin
Event|Event|Hospital Course|10940,10948|false|false|false|||warfarin
Drug|Biomedical or Dental Material|Hospital Course|10956,10962|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|10966,10974|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|10969,10974|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|10969,10974|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Event|Hospital Course|10978,10982|false|false|false|||WEEK
Finding|Intellectual Product|Hospital Course|10978,10982|false|false|false|C1561540|Transaction counts and value totals - week|WEEK
Drug|Biomedical or Dental Material|Hospital Course|10993,10999|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|10993,10999|false|false|false|||Tablet
Event|Event|Hospital Course|11001,11008|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|11001,11008|false|false|false|C0807726|refill|Refills
Drug|Hazardous or Poisonous Substance|Hospital Course|11016,11024|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|Hospital Course|11016,11024|false|false|false|C0043031|warfarin|Warfarin
Drug|Pharmacologic Substance|Hospital Course|11016,11024|false|false|false|C0043031|warfarin|Warfarin
Finding|Intellectual Product|Hospital Course|11036,11040|false|false|false|C1561540|Transaction counts and value totals - week|WEEK
Event|Event|Hospital Course|11048,11050|false|false|false|||RX
Drug|Hazardous or Poisonous Substance|Hospital Course|11052,11060|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|Hospital Course|11052,11060|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|Hospital Course|11052,11060|false|false|false|C0043031|warfarin|warfarin
Event|Event|Hospital Course|11052,11060|false|false|false|||warfarin
Drug|Biomedical or Dental Material|Hospital Course|11068,11074|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|11078,11086|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|11081,11086|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|11081,11086|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Event|Hospital Course|11090,11094|false|false|false|||WEEK
Finding|Intellectual Product|Hospital Course|11090,11094|false|false|false|C1561540|Transaction counts and value totals - week|WEEK
Drug|Biomedical or Dental Material|Hospital Course|11105,11111|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|11105,11111|false|false|false|||Tablet
Event|Event|Hospital Course|11113,11120|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|11113,11120|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|11128,11138|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|Hospital Course|11128,11138|false|false|false|C0016860|furosemide|Furosemide
Drug|Organic Chemical|Hospital Course|11159,11169|false|false|false|C0016860|furosemide|furosemide
Drug|Pharmacologic Substance|Hospital Course|11159,11169|false|false|false|C0016860|furosemide|furosemide
Event|Event|Hospital Course|11159,11169|false|false|false|||furosemide
Drug|Biomedical or Dental Material|Hospital Course|11178,11184|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|11188,11196|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|11191,11196|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|11191,11196|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Biomedical or Dental Material|Hospital Course|11213,11219|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|11213,11219|false|false|false|||Tablet
Event|Event|Hospital Course|11221,11228|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|11221,11228|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|11236,11247|false|false|false|C0002144|allopurinol|Allopurinol
Drug|Pharmacologic Substance|Hospital Course|11236,11247|false|false|false|C0002144|allopurinol|Allopurinol
Event|Event|Hospital Course|11270,11273|false|false|false|||DAY
Finding|Idea or Concept|Hospital Course|11270,11273|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|DAY
Finding|Intellectual Product|Hospital Course|11270,11273|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|DAY
Drug|Organic Chemical|Hospital Course|11279,11290|false|false|false|C0002144|allopurinol|allopurinol
Drug|Pharmacologic Substance|Hospital Course|11279,11290|false|false|false|C0002144|allopurinol|allopurinol
Drug|Biomedical or Dental Material|Hospital Course|11300,11306|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|11310,11318|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|11313,11318|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|11313,11318|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Event|Hospital Course|11331,11334|false|false|false|||DAY
Finding|Idea or Concept|Hospital Course|11331,11334|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|DAY
Finding|Intellectual Product|Hospital Course|11331,11334|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|DAY
Event|Activity|Hospital Course|11335,11339|false|false|false|C1880359|Dispense (activity)|Disp
Finding|Gene or Genome|Hospital Course|11335,11339|false|false|false|C2828567|PRSS30P gene|Disp
Drug|Biomedical or Dental Material|Hospital Course|11346,11352|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|11353,11360|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|11353,11360|false|false|false|C0807726|refill|Refills
Event|Event|Hospital Course|11383,11389|false|false|false|||Dinner
Finding|Daily or Recreational Activity|Hospital Course|11383,11389|false|false|false|C4048877|Dinner|Dinner
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11394,11401|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|Hospital Course|11394,11401|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|Hospital Course|11394,11401|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|Hospital Course|11394,11401|false|false|false|||insulin
Finding|Gene or Genome|Hospital Course|11394,11401|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|Hospital Course|11394,11401|false|false|false|C0202098|Insulin measurement|insulin
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11394,11405|false|false|false|C0021658|insulin isophane|insulin NPH
Drug|Hormone|Hospital Course|11394,11405|false|false|false|C0021658|insulin isophane|insulin NPH
Drug|Pharmacologic Substance|Hospital Course|11394,11405|false|false|false|C0021658|insulin isophane|insulin NPH
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11402,11405|false|false|false|C0027442|Nasopharynx|NPH
Disorder|Disease or Syndrome|Hospital Course|11402,11405|false|false|false|C0020258|Hydrocephalus, Normal Pressure|NPH
Event|Event|Hospital Course|11402,11405|false|false|false|||NPH
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11425,11432|false|false|false|C0020171;C0020172;C3538423|Humulin;Humulin S;Humulin insulin|Humulin
Drug|Hormone|Hospital Course|11425,11432|false|false|false|C0020171;C0020172;C3538423|Humulin;Humulin S;Humulin insulin|Humulin
Drug|Pharmacologic Substance|Hospital Course|11425,11432|false|false|false|C0020171;C0020172;C3538423|Humulin;Humulin S;Humulin insulin|Humulin
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11425,11438|false|false|false|C0306367|HumuLIN 70/30|Humulin 70/30
Drug|Hormone|Hospital Course|11425,11438|false|false|false|C0306367|HumuLIN 70/30|Humulin 70/30
Drug|Pharmacologic Substance|Hospital Course|11425,11438|false|false|false|C0306367|HumuLIN 70/30|Humulin 70/30
Drug|Clinical Drug|Hospital Course|11425,11446|false|false|false|C2683543|3 ML insulin isophane, human 70 UNT/ML / insulin, regular, human 30 UNT/ML Pen Injector [Humulin]|Humulin 70/30 KwikPen
Event|Event|Hospital Course|11478,11480|false|false|false|||SC
Event|Event|Hospital Course|11481,11485|false|false|false|||Take
Event|Activity|Hospital Course|11508,11512|false|false|false|C1880359|Dispense (activity)|Disp
Finding|Gene or Genome|Hospital Course|11508,11512|false|false|false|C2828567|PRSS30P gene|Disp
Finding|Intellectual Product|Hospital Course|11518,11525|false|false|false|C1704709|Computer program package|Package
Event|Event|Hospital Course|11526,11533|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|11526,11533|false|false|false|C0807726|refill|Refills
Event|Event|Hospital Course|11540,11549|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|11540,11549|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|11540,11549|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|11540,11549|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|11540,11549|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|11540,11561|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|11540,11561|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|11550,11561|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|11550,11561|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|11550,11561|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|Hospital Course|11563,11567|false|false|false|||Home
Finding|Idea or Concept|Hospital Course|11563,11567|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|11563,11567|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|11563,11567|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|Hospital Course|11573,11580|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|Hospital Course|11573,11580|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|Hospital Course|11583,11591|false|false|false|||Facility
Finding|Intellectual Product|Hospital Course|11583,11591|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|Hospital Course|11599,11608|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|11599,11608|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|11599,11608|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|11599,11608|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|11599,11608|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|11599,11618|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|11609,11618|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|11609,11618|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|11609,11618|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|11609,11618|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|11609,11618|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Disease or Syndrome|Principle Diagnosis|11639,11645|false|false|false|C0002871|Anemia|Anemia
Event|Event|Principle Diagnosis|11639,11645|false|false|false|||Anemia
Disorder|Disease or Syndrome|Principle Diagnosis|11646,11670|false|false|false|C0018802|Congestive heart failure|Congestive heart failure
Finding|Finding|Principle Diagnosis|11646,11683|false|false|false|C3532952|Exacerbation of congestive heart failure|Congestive heart failure exacerbation
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|11657,11662|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Principle Diagnosis|11657,11662|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Principle Diagnosis|11657,11662|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|Principle Diagnosis|11657,11670|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Event|Event|Principle Diagnosis|11663,11670|false|false|false|||failure
Finding|Functional Concept|Principle Diagnosis|11663,11670|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|Principle Diagnosis|11663,11670|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|Principle Diagnosis|11663,11670|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|Principle Diagnosis|11671,11683|false|false|false|||exacerbation
Finding|Finding|Principle Diagnosis|11671,11683|false|false|false|C4086268|Exacerbation|exacerbation
Disorder|Neoplastic Process|Principle Diagnosis|11685,11694|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Event|Event|Principle Diagnosis|11685,11694|false|false|false|||Secondary
Finding|Functional Concept|Principle Diagnosis|11685,11694|false|false|false|C1522484|metastatic qualifier|Secondary
Attribute|Clinical Attribute|Principle Diagnosis|11685,11704|false|false|false|C4255018||Secondary diagnosis
Finding|Finding|Principle Diagnosis|11685,11704|false|false|false|C0332138|Secondary diagnosis|Secondary diagnosis
Attribute|Clinical Attribute|Principle Diagnosis|11695,11704|false|false|false|C0945731||diagnosis
Event|Event|Principle Diagnosis|11695,11704|false|false|false|||diagnosis
Finding|Classification|Principle Diagnosis|11695,11704|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|Principle Diagnosis|11695,11704|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|Principle Diagnosis|11695,11704|false|false|false|C0011900|Diagnosis|diagnosis
Disorder|Disease or Syndrome|Principle Diagnosis|11706,11718|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|Principle Diagnosis|11706,11718|false|false|false|||Hypertension
Event|Event|Principle Diagnosis|11720,11724|false|false|false|||DMII
Drug|Amino Acid, Peptide, or Protein|Principle Diagnosis|11728,11735|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|Principle Diagnosis|11728,11735|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|Principle Diagnosis|11728,11735|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|Principle Diagnosis|11728,11735|false|false|false|||insulin
Finding|Gene or Genome|Principle Diagnosis|11728,11735|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|Principle Diagnosis|11728,11735|false|false|false|C0202098|Insulin measurement|insulin
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|11737,11745|false|false|false|C0018787|Heart|Coronary
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|11737,11752|false|false|false|C0205042|Coronary artery|Coronary artery
Disorder|Disease or Syndrome|Principle Diagnosis|11737,11760|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|Coronary artery disease
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|11746,11752|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|Principle Diagnosis|11746,11752|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Disorder|Disease or Syndrome|Principle Diagnosis|11746,11760|false|false|false|C0852949|Arteriopathic disease|artery disease
Disorder|Disease or Syndrome|Principle Diagnosis|11753,11760|false|false|false|C0012634|Disease|disease
Event|Event|Principle Diagnosis|11753,11760|false|false|false|||disease
Attribute|Clinical Attribute|Principle Diagnosis|11762,11767|false|false|false|C1300072|Tumor stage|Stage
Event|Event|Principle Diagnosis|11771,11778|false|false|false|||chronic
Finding|Intellectual Product|Principle Diagnosis|11771,11778|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Principle Diagnosis|11771,11778|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|Principle Diagnosis|11771,11793|false|false|false|C1561643|Chronic Kidney Diseases|chronic kidney disease
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|11779,11785|false|false|false|C0022646;C0227665|Both kidneys;Kidney|kidney
Disorder|Neoplastic Process|Principle Diagnosis|11779,11785|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|kidney
Finding|Sign or Symptom|Principle Diagnosis|11779,11785|false|false|false|C0812426|Kidney problem|kidney
Procedure|Diagnostic Procedure|Principle Diagnosis|11779,11785|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Procedure|Therapeutic or Preventive Procedure|Principle Diagnosis|11779,11785|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Disorder|Disease or Syndrome|Principle Diagnosis|11779,11793|false|false|false|C0022658|Kidney Diseases|kidney disease
Disorder|Disease or Syndrome|Principle Diagnosis|11786,11793|false|false|false|C0012634|Disease|disease
Event|Event|Principle Diagnosis|11786,11793|false|false|false|||disease
Attribute|Clinical Attribute|Principle Diagnosis|11794,11798|false|false|false|C4318566|Deep Resection Margin|Deep
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|11794,11803|false|false|false|C0226514|Structure of deep vein|Deep vein
Disorder|Disease or Syndrome|Principle Diagnosis|11794,11814|false|false|false|C0149871;C0340708|Deep Vein Thrombosis;Deep vein thrombosis of lower limb|Deep vein thrombosis
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|11799,11803|false|false|false|C0042449|Veins|vein
Finding|Pathologic Function|Principle Diagnosis|11799,11814|false|false|false|C0042487|Venous Thrombosis|vein thrombosis
Event|Event|Principle Diagnosis|11804,11814|false|false|false|||thrombosis
Finding|Pathologic Function|Principle Diagnosis|11804,11814|false|false|false|C0040053|Thrombosis|thrombosis
Finding|Mental Process|Discharge Condition|11839,11845|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|11839,11852|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|11839,11852|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|11846,11852|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|11846,11852|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|11854,11859|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|11854,11859|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|11864,11872|false|false|false|||coherent
Finding|Finding|Discharge Condition|11864,11872|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|11874,11879|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|11874,11896|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|11874,11896|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|11883,11896|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|11883,11896|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|11883,11896|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|11898,11903|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|11898,11903|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|11898,11903|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|11898,11903|false|false|false|||Alert
Finding|Finding|Discharge Condition|11898,11903|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|11898,11903|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|11898,11903|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|11908,11919|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|11908,11919|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|11921,11929|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|11921,11929|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|11921,11929|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|11930,11936|false|false|false|C5889824||Status
Event|Event|Discharge Condition|11930,11936|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|11930,11936|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|Discharge Condition|11938,11948|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|11938,11948|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|11938,11948|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|11938,11948|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|11951,11959|false|false|false|||requires
Event|Event|Discharge Condition|11960,11970|false|false|false|||assistance
Finding|Social Behavior|Discharge Condition|11960,11970|false|false|false|C0018896|Helping Behavior|assistance
Drug|Amino Acid, Peptide, or Protein|Discharge Condition|11974,11977|false|false|false|C1454018|AICDA protein, human|aid
Drug|Enzyme|Discharge Condition|11974,11977|false|false|false|C1454018|AICDA protein, human|aid
Event|Event|Discharge Condition|11974,11977|false|false|false|||aid
Finding|Gene or Genome|Discharge Condition|11974,11977|false|false|false|C1421876;C3540469|AICDA gene;AICDA wt Allele|aid
Procedure|Therapeutic or Preventive Procedure|Discharge Condition|11974,11977|false|false|false|C0021588;C0280108|AID - Artificial insemination by donor;dacarbazine/doxorubicin/ifosfamide protocol|aid
Event|Event|Discharge Condition|11979,11985|false|false|false|||walker
Finding|Gene or Genome|Discharge Instructions|12024,12028|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|Discharge Instructions|12044,12052|false|false|false|||pleasure
Finding|Intellectual Product|Discharge Instructions|12044,12052|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|Discharge Instructions|12044,12052|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Event|Discharge Instructions|12053,12059|false|false|false|||caring
Event|Event|Discharge Instructions|12078,12086|false|false|false|||admitted
Event|Event|Discharge Instructions|12095,12103|false|false|false|||hospital
Finding|Idea or Concept|Discharge Instructions|12095,12103|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|Discharge Instructions|12109,12116|false|false|false|||fatigue
Finding|Sign or Symptom|Discharge Instructions|12109,12116|false|false|false|C0015672|Fatigue|fatigue
Anatomy|Body Location or Region|Discharge Instructions|12118,12123|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Discharge Instructions|12118,12123|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Discharge Instructions|12118,12128|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Discharge Instructions|12118,12128|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Discharge Instructions|12124,12128|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|12124,12128|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|12124,12128|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|12124,12128|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Discharge Instructions|12134,12143|false|false|false|||shortness
Attribute|Clinical Attribute|Discharge Instructions|12134,12153|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|Discharge Instructions|12134,12153|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|Discharge Instructions|12147,12153|false|false|false|C0225386|Breath|breath
Event|Event|Discharge Instructions|12165,12170|false|false|false|||found
Finding|Gene or Genome|Discharge Instructions|12179,12186|false|false|false|C1825291|FEZF2 gene|too few
Finding|Finding|Discharge Instructions|12187,12190|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Finding|Gene or Genome|Discharge Instructions|12187,12190|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Anatomy|Cell|Discharge Instructions|12187,12202|false|false|false|C0014792|Erythrocytes|red blood cells
Drug|Pharmacologic Substance|Discharge Instructions|12187,12202|false|false|false|C0014792;C1277078|Erythrocytes;Red blood cells, blood product|red blood cells
Disorder|Disease or Syndrome|Discharge Instructions|12191,12196|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Discharge Instructions|12191,12196|false|false|false|||blood
Finding|Body Substance|Discharge Instructions|12191,12196|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Anatomy|Cell|Discharge Instructions|12191,12202|false|false|false|C0005773|Blood Cells|blood cells
Anatomy|Cell|Discharge Instructions|12197,12202|false|false|false|C0007634|Cells|cells
Disorder|Disease or Syndrome|Discharge Instructions|12204,12210|false|false|false|C0002871|Anemia|anemia
Event|Event|Discharge Instructions|12204,12210|false|false|false|||anemia
Disorder|Disease or Syndrome|Discharge Instructions|12226,12231|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Discharge Instructions|12226,12231|false|false|false|||blood
Finding|Body Substance|Discharge Instructions|12226,12231|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Event|Discharge Instructions|12242,12250|false|false|false|||symptoms
Finding|Functional Concept|Discharge Instructions|12242,12250|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Discharge Instructions|12242,12250|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|Discharge Instructions|12251,12259|false|false|false|||improved
Event|Event|Discharge Instructions|12284,12289|false|false|false|||found
Finding|Finding|Discharge Instructions|12299,12307|false|false|false|C3843660|Too much|too much
Finding|Finding|Discharge Instructions|12303,12307|false|false|false|C4281574|Much|much
Drug|Substance|Discharge Instructions|12308,12313|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|Discharge Instructions|12308,12313|false|false|false|||fluid
Finding|Intellectual Product|Discharge Instructions|12308,12313|false|false|false|C1546638|Fluid Specimen Code|fluid
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|12322,12326|false|false|false|C1140621|Leg|legs
Attribute|Clinical Attribute|Discharge Instructions|12322,12326|false|false|false|C5781420||legs
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|12331,12336|false|false|false|C0024109|Lung|lungs
Event|Event|Discharge Instructions|12341,12348|false|false|false|||treated
Drug|Pharmacologic Substance|Discharge Instructions|12361,12369|false|false|false|C0012798;C5399719|Diuretic [APC];Diuretics|diuretic
Event|Event|Discharge Instructions|12361,12369|false|false|false|||diuretic
Event|Event|Discharge Instructions|12377,12383|false|false|false|||helped
Event|Event|Discharge Instructions|12384,12393|false|false|false|||eliminate
Drug|Substance|Discharge Instructions|12398,12403|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|Discharge Instructions|12398,12403|false|false|false|||fluid
Finding|Intellectual Product|Discharge Instructions|12398,12403|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|Discharge Instructions|12437,12441|false|false|false|||call
Attribute|Clinical Attribute|Discharge Instructions|12448,12454|false|false|false|C0944911||weight
Event|Event|Discharge Instructions|12448,12454|false|false|false|||weight
Finding|Finding|Discharge Instructions|12448,12454|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|Discharge Instructions|12448,12454|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|Discharge Instructions|12448,12454|false|false|false|C1305866|Weighing patient|weight
Event|Event|Discharge Instructions|12455,12459|false|false|false|||goes
Procedure|Laboratory Procedure|Discharge Instructions|12476,12479|false|false|false|C3161851|liquid-based cytology (procedure)|lbs
Procedure|Health Care Activity|Discharge Instructions|12509,12517|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|12518,12530|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|12518,12530|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|12518,12530|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

