 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|29,33
No|34,36
:|36,37
_|40,41
_|41,42
_|42,43
<EOL>|43,44
<EOL>|45,46
Admission|46,55
Date|56,60
:|60,61
_|63,64
_|64,65
_|65,66
Discharge|80,89
Date|90,94
:|94,95
_|98,99
_|99,100
_|100,101
<EOL>|101,102
<EOL>|103,104
Date|104,108
of|109,111
Birth|112,117
:|117,118
_|120,121
_|121,122
_|122,123
Sex|136,139
:|139,140
F|143,144
<EOL>|144,145
<EOL>|146,147
Service|147,154
:|154,155
NEUROSURGERY|156,168
<EOL>|168,169
<EOL>|170,171
Penicillins|183,194
/|195,196
Paxil|197,202
/|203,204
Wellbutrin|205,215
<EOL>|215,216
<EOL>|217,218
Attending|218,227
:|227,228
_|229,230
_|230,231
_|231,232
.|232,233
<EOL>|233,234
<EOL>|235,236
exposed|253,260
craniotomy|261,271
hardware|272,280
<EOL>|280,281
<EOL>|282,283
Major|283,288
Surgical|289,297
or|298,300
Invasive|301,309
Procedure|310,319
:|319,320
<EOL>|320,321
wound|321,326
revision|327,335
and|336,339
hardware|340,348
removal|349,356
<EOL>|356,357
<EOL>|357,358
<EOL>|359,360
This|388,392
is|393,395
a|396,397
_|398,399
_|399,400
_|400,401
year|402,406
old|407,410
female|411,417
with|418,422
prior|423,428
surgery|429,436
which|437,442
<EOL>|442,443
includes|443,451
right|452,457
parietal|458,466
anaplastic|467,477
astrocytoma|478,489
with|490,494
Craniotomy|495,505
<EOL>|505,506
for|506,509
resection|510,519
on|520,522
_|523,524
_|524,525
_|525,526
by|527,529
Dr.|530,533
_|534,535
_|535,536
_|536,537
in|538,540
_|541,542
_|542,543
_|543,544
<EOL>|545,546
followed|546,554
<EOL>|554,555
by|555,557
involved|558,566
-|566,567
field|567,572
irradiation|573,584
to|585,587
6,120|588,593
cGy|594,597
_|598,599
_|599,600
_|600,601
in|602,604
_|605,606
_|606,607
_|607,608
,|608,609
<EOL>|609,610
3|610,611
cycles|612,618
of|619,621
Temodar|622,629
ended|630,635
_|636,637
_|637,638
_|638,639
and|640,643
a|644,645
second|646,652
craniotomy|653,663
for|664,667
tumor|668,673
<EOL>|673,674
recurrence|674,684
on|685,687
_|688,689
_|689,690
_|690,691
by|692,694
Dr.|695,698
_|699,700
_|700,701
_|701,702
at|703,705
_|706,707
_|707,708
_|708,709
with|710,714
PCV|715,718
(|718,719
comb|719,723
chemo|724,729
)|729,730
<EOL>|730,731
_|731,732
_|732,733
_|733,734
-|735,736
_|737,738
_|738,739
_|739,740
.|740,741
<EOL>|743,744
<EOL>|744,745
The|745,748
patient|749,756
presents|757,765
today|766,771
with|772,776
_|777,778
_|778,779
_|779,780
month|781,786
history|787,794
of|795,797
pruritus|798,806
on|807,809
<EOL>|809,810
the|810,813
top|814,817
of|818,820
her|821,824
head|825,829
.|829,830
She|832,835
reports|836,843
that|844,848
she|849,852
had|853,856
her|857,860
husband|861,868
look|869,873
<EOL>|873,874
at|874,876
the|877,880
top|881,884
of|885,887
her|888,891
head|892,896
_|897,898
_|898,899
_|899,900
days|901,905
ago|906,909
and|910,913
saw|914,917
that|918,922
metal|923,928
hardware|929,937
<EOL>|937,938
from|938,942
her|943,946
prior|947,952
surgery|953,960
was|961,964
present|965,972
.|972,973
The|975,978
patient|979,986
and|987,990
her|991,994
husband|995,1002
<EOL>|1002,1003
presented|1003,1012
to|1013,1015
their|1016,1021
local|1022,1027
Emergency|1028,1037
and|1038,1041
was|1042,1045
told|1046,1050
to|1051,1053
follow|1054,1060
up|1061,1063
<EOL>|1063,1064
here|1064,1068
.|1068,1069
The|1071,1074
patient|1075,1082
denies|1083,1089
fever|1090,1095
,|1095,1096
chills|1097,1103
,|1103,1104
nausea|1105,1111
vomiting|1112,1120
,|1120,1121
nuchal|1122,1128
<EOL>|1128,1129
rigidity|1129,1137
,|1137,1138
numbness|1139,1147
or|1148,1150
tingling|1151,1159
sensation|1160,1169
,|1169,1170
vision|1171,1177
or|1178,1180
hearing|1181,1188
<EOL>|1188,1189
changes|1189,1196
,|1196,1197
bowel|1198,1203
or|1204,1206
bladder|1207,1214
incontinence|1215,1227
.|1227,1228
She|1230,1233
denies|1234,1240
new|1241,1244
onset|1245,1250
<EOL>|1250,1251
weakness|1251,1259
.|1259,1260
She|1262,1265
reports|1266,1273
baseline|1274,1282
tremors|1283,1290
in|1291,1293
arms|1294,1298
due|1299,1302
to|1303,1305
her|1306,1309
<EOL>|1309,1310
hyperthyroid|1310,1322
disease|1323,1330
and|1331,1334
baseline|1335,1343
left|1344,1348
sided|1349,1354
weakness|1355,1363
since|1364,1369
her|1370,1373
<EOL>|1373,1374
initial|1374,1381
surgery|1382,1389
.|1389,1390
She|1392,1395
does|1396,1400
not|1401,1404
ambulate|1405,1413
with|1414,1418
a|1419,1420
walker|1421,1427
<EOL>|1428,1429
<EOL>|1429,1430
<EOL>|1431,1432
right|1454,1459
parietal|1460,1468
anaplastic|1469,1479
astrocytoma|1480,1491
,|1491,1492
Craniotomy|1492,1502
_|1503,1504
_|1504,1505
_|1505,1506
by|1507,1509
<EOL>|1509,1510
Dr.|1510,1513
_|1514,1515
_|1515,1516
_|1516,1517
in|1518,1520
_|1521,1522
_|1522,1523
_|1523,1524
irradiation|1525,1536
to|1537,1539
6,120|1540,1545
<EOL>|1545,1546
cGy|1546,1549
_|1550,1551
_|1551,1552
_|1552,1553
in|1554,1556
_|1557,1558
_|1558,1559
_|1559,1560
,|1560,1561
3|1561,1562
cycles|1563,1569
of|1570,1572
Temodar|1573,1580
ended|1581,1586
_|1587,1588
_|1588,1589
_|1589,1590
<EOL>|1590,1591
craniotomy|1591,1601
on|1602,1604
_|1605,1606
_|1606,1607
_|1607,1608
by|1609,1611
Dr.|1612,1615
_|1616,1617
_|1617,1618
_|1618,1619
at|1620,1622
_|1623,1624
_|1624,1625
_|1625,1626
_|1627,1628
_|1628,1629
_|1629,1630
-|1631,1632
<EOL>|1632,1633
_|1633,1634
_|1634,1635
_|1635,1636
for|1637,1640
2|1641,1642
weeks|1643,1648
only|1649,1653
_|1654,1655
_|1655,1656
_|1656,1657
disease|1658,1665
since|1666,1671
_|1672,1673
_|1673,1674
_|1674,1675
,|1675,1676
<EOL>|1676,1677
tubal|1677,1682
ligation|1683,1691
,|1691,1692
tonsillectomy|1692,1705
,|1705,1706
bronchitis|1707,1717
,|1717,1718
depression|1719,1729
.|1729,1730
<EOL>|1730,1731
seizures|1731,1739
<EOL>|1739,1740
<EOL>|1740,1741
<EOL>|1742,1743
:|1757,1758
<EOL>|1758,1759
_|1759,1760
_|1760,1761
_|1761,1762
<EOL>|1762,1763
:|1777,1778
<EOL>|1778,1779
NC|1779,1781
<EOL>|1781,1782
<EOL>|1783,1784
O|1799,1800
:|1800,1801
T|1802,1803
:|1803,1804
96.7|1804,1808
BP|1810,1812
:|1812,1813
139|1814,1817
/|1817,1818
73|1818,1820
HR|1822,1824
:|1824,1825
114|1825,1828
R|1832,1833
:|1833,1834
20|1834,1836
O2Sats|1840,1846
:|1846,1847
100|1848,1851
%|1851,1852
ra|1853,1855
<EOL>|1855,1856
Gen|1856,1859
:|1859,1860
WD|1861,1863
/|1863,1864
WN|1864,1866
,|1866,1867
comfortable|1868,1879
,|1879,1880
NAD|1881,1884
.|1884,1885
<EOL>|1885,1886
HEENT|1886,1891
:|1891,1892
Pupils|1893,1899
:|1899,1900
3|1900,1901
-|1901,1902
2mm|1902,1905
bilat|1906,1911
EOMs|1920,1924
:|1924,1925
intact|1926,1932
<EOL>|1932,1933
Neck|1933,1937
:|1937,1938
Supple|1939,1945
.|1945,1946
<EOL>|1946,1947
Extrem|1947,1953
:|1953,1954
Warm|1955,1959
and|1960,1963
well|1964,1968
-|1968,1969
perfused|1969,1977
,|1977,1978
arms|1979,1983
hands|1984,1989
tremulous|1990,1999
-|1999,2000
(|2001,2002
patient|2002,2009
<EOL>|2009,2010
states|2010,2016
this|2017,2021
is|2022,2024
her|2025,2028
baseline|2029,2037
due|2038,2041
to|2042,2044
hyperthyroid|2045,2057
disease|2058,2065
)|2065,2066
<EOL>|2066,2067
Neuro|2067,2072
:|2072,2073
<EOL>|2073,2074
Mental|2074,2080
status|2081,2087
:|2087,2088
Awake|2089,2094
and|2095,2098
alert|2099,2104
,|2104,2105
cooperative|2106,2117
with|2118,2122
exam|2123,2127
,|2127,2128
normal|2129,2135
<EOL>|2135,2136
affect|2136,2142
.|2142,2143
<EOL>|2143,2144
Orientation|2144,2155
:|2155,2156
Oriented|2157,2165
to|2166,2168
person|2169,2175
,|2175,2176
place|2177,2182
,|2182,2183
and|2184,2187
date|2188,2192
.|2192,2193
<EOL>|2193,2194
Recall|2194,2200
:|2200,2201
_|2202,2203
_|2203,2204
_|2204,2205
objects|2206,2213
at|2214,2216
5|2217,2218
minutes|2219,2226
.|2226,2227
<EOL>|2227,2228
Language|2228,2236
:|2236,2237
Speech|2238,2244
fluent|2245,2251
with|2252,2256
good|2257,2261
comprehension|2262,2275
and|2276,2279
repetition|2280,2290
.|2290,2291
<EOL>|2291,2292
Naming|2292,2298
intact|2299,2305
.|2305,2306
No|2307,2309
dysarthria|2310,2320
or|2321,2323
paraphasic|2324,2334
errors|2335,2341
.|2341,2342
<EOL>|2342,2343
<EOL>|2343,2344
Cranial|2344,2351
Nerves|2352,2358
:|2358,2359
<EOL>|2359,2360
I|2360,2361
:|2361,2362
Not|2363,2366
tested|2367,2373
<EOL>|2373,2374
II|2374,2376
:|2376,2377
Pupils|2378,2384
equally|2385,2392
round|2393,2398
and|2399,2402
reactive|2403,2411
to|2412,2414
light|2415,2420
,|2420,2421
3|2423,2424
to|2425,2427
2|2428,2429
<EOL>|2429,2430
mm|2430,2432
bilaterally|2433,2444
.|2444,2445
Visual|2446,2452
fields|2453,2459
are|2460,2463
full|2464,2468
to|2469,2471
confrontation|2472,2485
.|2485,2486
<EOL>|2486,2487
III|2487,2490
,|2490,2491
IV|2492,2494
,|2494,2495
VI|2496,2498
:|2498,2499
Extraocular|2500,2511
movements|2512,2521
intact|2522,2528
bilaterally|2529,2540
without|2541,2548
<EOL>|2548,2549
nystagmus|2549,2558
.|2558,2559
<EOL>|2559,2560
V|2560,2561
,|2561,2562
VII|2563,2566
:|2566,2567
Facial|2568,2574
strength|2575,2583
and|2584,2587
sensation|2588,2597
intact|2598,2604
and|2605,2608
symmetric|2609,2618
.|2618,2619
<EOL>|2619,2620
VIII|2620,2624
:|2624,2625
Hearing|2626,2633
intact|2634,2640
to|2641,2643
voice|2644,2649
.|2649,2650
<EOL>|2650,2651
IX|2651,2653
,|2653,2654
X|2655,2656
:|2656,2657
Palatal|2658,2665
elevation|2666,2675
symmetrical|2676,2687
.|2687,2688
<EOL>|2688,2689
XI|2689,2691
:|2691,2692
Sternocleidomastoid|2693,2712
and|2713,2716
trapezius|2717,2726
normal|2727,2733
bilaterally|2734,2745
.|2745,2746
<EOL>|2746,2747
XII|2747,2750
:|2750,2751
Tongue|2752,2758
midline|2759,2766
without|2767,2774
fasciculations|2775,2789
.|2789,2790
<EOL>|2790,2791
<EOL>|2791,2792
Motor|2792,2797
:|2797,2798
Normal|2799,2805
bulk|2806,2810
and|2811,2814
tone|2815,2819
bilaterally|2820,2831
.|2831,2832
No|2833,2835
abnormal|2836,2844
movements|2845,2854
,|2854,2855
<EOL>|2855,2856
tremors|2856,2863
.|2863,2864
Strength|2865,2873
full|2874,2878
power|2879,2884
_|2885,2886
_|2886,2887
_|2887,2888
on|2889,2891
right|2892,2897
4|2898,2899
+|2899,2900
/|2900,2901
5|2901,2902
on|2903,2905
left|2906,2910
.|2910,2911
No|2912,2914
<EOL>|2914,2915
pronator|2915,2923
drift|2924,2929
<EOL>|2929,2930
<EOL>|2930,2931
Sensation|2931,2940
:|2940,2941
Intact|2942,2948
to|2949,2951
light|2952,2957
touch|2958,2963
bilaterally|2964,2975
.|2975,2976
<EOL>|2976,2977
<EOL>|2977,2978
Toes|2978,2982
downgoing|2983,2992
bilaterally|2993,3004
<EOL>|3004,3005
<EOL>|3005,3006
Coordination|3006,3018
:|3018,3019
normal|3020,3026
on|3027,3029
finger|3030,3036
-|3036,3037
nose|3037,3041
-|3041,3042
finger|3042,3048
,|3048,3049
rapid|3050,3055
alternating|3056,3067
<EOL>|3067,3068
movements|3068,3077
,|3077,3078
heel|3079,3083
to|3084,3086
shin|3087,3091
<EOL>|3091,3092
<EOL>|3092,3093
<EOL>|3094,3095
Pertinent|3095,3104
Results|3105,3112
:|3112,3113
<EOL>|3113,3114
CT|3114,3116
Head|3117,3121
<EOL>|3121,3122
1|3122,3123
.|3123,3124
No|3125,3127
evidence|3128,3136
of|3137,3139
abscess|3140,3147
formation|3148,3157
.|3157,3158
<EOL>|3159,3160
2.|3160,3162
Stable|3163,3169
appearance|3170,3180
of|3181,3183
postoperative|3184,3197
changes|3198,3205
related|3206,3213
to|3214,3216
right|3217,3222
<EOL>|3223,3224
frontal|3224,3231
mass|3232,3236
resection|3237,3246
with|3247,3251
residual|3252,3260
encephalomalacia|3261,3277
and|3278,3281
edema|3282,3287
<EOL>|3288,3289
in|3289,3291
a|3292,3293
similar|3294,3301
distribution|3302,3314
as|3315,3317
_|3318,3319
_|3319,3320
_|3320,3321
MR|3322,3324
exam|3325,3329
.|3329,3330
<EOL>|3331,3332
<EOL>|3332,3333
<EOL>|3334,3335
patient|3358,3365
presented|3366,3375
to|3376,3378
the|3379,3382
ED|3383,3385
at|3386,3388
_|3389,3390
_|3390,3391
_|3391,3392
on|3393,3395
_|3396,3397
_|3397,3398
_|3398,3399
with|3400,3404
complaints|3405,3415
of|3416,3418
<EOL>|3419,3420
itchy|3420,3425
head|3426,3430
and|3431,3434
exposed|3435,3442
hardware|3443,3451
.|3451,3452
She|3454,3457
was|3458,3461
admitted|3462,3470
to|3471,3473
the|3474,3477
floor|3478,3483
<EOL>|3484,3485
for|3485,3488
observation|3489,3500
and|3501,3504
pre-operative|3505,3518
planning|3519,3527
.|3527,3528
On|3530,3532
3.5|3533,3536
she|3537,3540
was|3541,3544
<EOL>|3545,3546
taken|3546,3551
to|3552,3554
the|3555,3558
OR|3559,3561
for|3562,3565
wound|3566,3571
revision|3572,3580
and|3581,3584
removal|3585,3592
of|3593,3595
the|3596,3599
exposed|3600,3607
<EOL>|3608,3609
hardware|3609,3617
.|3617,3618
She|3620,3623
tolerated|3624,3633
the|3634,3637
procedure|3638,3647
well|3648,3652
and|3653,3656
was|3657,3660
transferred|3661,3672
<EOL>|3673,3674
to|3674,3676
the|3677,3680
_|3681,3682
_|3682,3683
_|3683,3684
post-operatively|3685,3701
.|3701,3702
She|3704,3707
was|3708,3711
transferred|3712,3723
to|3724,3726
the|3727,3730
floor|3731,3736
<EOL>|3737,3738
for|3738,3741
further|3742,3749
management|3750,3760
and|3761,3764
remained|3765,3773
stable|3774,3780
.|3780,3781
On|3783,3785
the|3786,3789
morning|3790,3797
of|3798,3800
<EOL>|3801,3802
_|3802,3803
_|3803,3804
_|3804,3805
she|3806,3809
was|3810,3813
deemed|3814,3820
fit|3821,3824
for|3825,3828
discharge|3829,3838
and|3839,3842
was|3843,3846
given|3847,3852
instructions|3853,3865
<EOL>|3866,3867
for|3867,3870
close|3871,3876
follow|3877,3883
-|3883,3884
up|3884,3886
of|3887,3889
her|3890,3893
incision|3894,3902
.|3902,3903
<EOL>|3905,3906
<EOL>|3907,3908
Medications|3908,3919
on|3920,3922
Admission|3923,3932
:|3932,3933
<EOL>|3933,3934
azathioprine|3934,3946
,|3946,3947
Pentasa|3948,3955
,|3955,3956
topiramate|3957,3967
,|3967,3968
<EOL>|3968,3969
alprazolam|3969,3979
,|3979,3980
omeprazole|3981,3991
,|3991,3992
zolpidem|3993,4001
,|4001,4002
venlafaxine|4003,4014
hcl|4015,4018
er|4019,4021
30|4022,4024
,|4024,4025
<EOL>|4025,4026
popylthiouracil|4026,4041
,|4041,4042
promethazine|4043,4055
-|4055,4056
patient|4057,4064
does|4065,4069
not|4070,4073
have|4074,4078
doses|4079,4084
at|4085,4087
<EOL>|4088,4089
the|4089,4092
<EOL>|4092,4093
time|4093,4097
of|4098,4100
the|4101,4104
exam|4105,4109
.|4109,4110
<EOL>|4110,4111
<EOL>|4111,4112
<EOL>|4113,4114
Discharge|4114,4123
Medications|4124,4135
:|4135,4136
<EOL>|4136,4137
1.|4137,4139
acetaminophen|4140,4153
325|4154,4157
mg|4158,4160
Tablet|4161,4167
Sig|4168,4171
:|4171,4172
_|4173,4174
_|4174,4175
_|4175,4176
Tablets|4177,4184
PO|4185,4187
Q6H|4188,4191
(|4192,4193
every|4193,4198
6|4199,4200
<EOL>|4201,4202
hours|4202,4207
)|4207,4208
as|4209,4211
needed|4212,4218
for|4219,4222
pain|4223,4227
.|4227,4228
<EOL>|4230,4231
2.|4231,4233
azathioprine|4234,4246
50|4247,4249
mg|4250,4252
Tablet|4253,4259
Sig|4260,4263
:|4263,4264
One|4265,4268
(|4269,4270
1|4270,4271
)|4271,4272
Tablet|4273,4279
PO|4280,4282
DAILY|4283,4288
<EOL>|4289,4290
(|4290,4291
Daily|4291,4296
)|4296,4297
.|4297,4298
<EOL>|4300,4301
3.|4301,4303
alprazolam|4304,4314
1|4315,4316
mg|4317,4319
Tablet|4320,4326
Sig|4327,4330
:|4330,4331
0.5|4332,4335
Tablet|4336,4342
PO|4343,4345
TID|4346,4349
(|4350,4351
3|4351,4352
times|4353,4358
a|4359,4360
day|4361,4364
)|4364,4365
<EOL>|4366,4367
as|4367,4369
needed|4370,4376
for|4377,4380
anxiety|4381,4388
.|4388,4389
<EOL>|4391,4392
4.|4392,4394
promethazine|4395,4407
25|4408,4410
mg|4411,4413
Tablet|4414,4420
Sig|4421,4424
:|4424,4425
One|4426,4429
(|4430,4431
1|4431,4432
)|4432,4433
Tablet|4434,4440
PO|4441,4443
Q6H|4444,4447
(|4448,4449
every|4449,4454
6|4455,4456
<EOL>|4457,4458
hours|4458,4463
)|4463,4464
as|4465,4467
needed|4468,4474
for|4475,4478
nausea|4479,4485
.|4485,4486
<EOL>|4488,4489
5.|4489,4491
omeprazole|4492,4502
20|4503,4505
mg|4506,4508
Capsule|4509,4516
,|4516,4517
Delayed|4518,4525
Release|4526,4533
(|4533,4534
E.C|4534,4537
.|4537,4538
)|4538,4539
Sig|4540,4543
:|4543,4544
One|4545,4548
(|4549,4550
1|4550,4551
)|4551,4552
<EOL>|4553,4554
Capsule|4554,4561
,|4561,4562
Delayed|4563,4570
Release|4571,4578
(|4578,4579
E.C|4579,4582
.|4582,4583
)|4583,4584
PO|4585,4587
DAILY|4588,4593
(|4594,4595
Daily|4595,4600
)|4600,4601
.|4601,4602
<EOL>|4604,4605
6.|4605,4607
cephalexin|4608,4618
500|4619,4622
mg|4623,4625
Capsule|4626,4633
Sig|4634,4637
:|4637,4638
One|4639,4642
(|4643,4644
1|4644,4645
)|4645,4646
Capsule|4647,4654
PO|4655,4657
Q6H|4658,4661
(|4662,4663
every|4663,4668
<EOL>|4669,4670
6|4670,4671
hours|4672,4677
)|4677,4678
for|4679,4682
13|4683,4685
days|4686,4690
.|4690,4691
<EOL>|4691,4692
Disp|4692,4696
:|4696,4697
*|4697,4698
52|4698,4700
Capsule|4701,4708
(|4708,4709
s|4709,4710
)|4710,4711
*|4711,4712
Refills|4713,4720
:|4720,4721
*|4721,4722
0|4722,4723
*|4723,4724
<EOL>|4724,4725
7.|4725,4727
docusate|4728,4736
sodium|4737,4743
100|4744,4747
mg|4748,4750
Capsule|4751,4758
Sig|4759,4762
:|4762,4763
One|4764,4767
(|4768,4769
1|4769,4770
)|4770,4771
Capsule|4772,4779
PO|4780,4782
BID|4783,4786
(|4787,4788
2|4788,4789
<EOL>|4790,4791
times|4791,4796
a|4797,4798
day|4799,4802
)|4802,4803
.|4803,4804
<EOL>|4806,4807
8.|4807,4809
zolpidem|4810,4818
5|4819,4820
mg|4821,4823
Tablet|4824,4830
Sig|4831,4834
:|4834,4835
Two|4836,4839
(|4840,4841
2|4841,4842
)|4842,4843
Tablet|4844,4850
PO|4851,4853
HS|4854,4856
(|4857,4858
at|4858,4860
bedtime|4861,4868
)|4868,4869
<EOL>|4870,4871
as|4871,4873
needed|4874,4880
for|4881,4884
for|4885,4888
sleep|4889,4894
.|4894,4895
<EOL>|4897,4898
9.|4898,4900
mesalamine|4901,4911
250|4912,4915
mg|4916,4918
Capsule|4919,4926
,|4926,4927
Extended|4928,4936
Release|4937,4944
Sig|4945,4948
:|4948,4949
Two|4950,4953
(|4954,4955
2|4955,4956
)|4956,4957
<EOL>|4958,4959
Capsule|4959,4966
,|4966,4967
Extended|4968,4976
Release|4977,4984
PO|4985,4987
QID|4988,4991
(|4992,4993
4|4993,4994
times|4995,5000
a|5001,5002
day|5003,5006
)|5006,5007
.|5007,5008
<EOL>|5010,5011
10.|5011,5014
topiramate|5015,5025
100|5026,5029
mg|5030,5032
Tablet|5033,5039
Sig|5040,5043
:|5043,5044
Two|5045,5048
(|5049,5050
2|5050,5051
)|5051,5052
Tablet|5053,5059
PO|5060,5062
BID|5063,5066
(|5067,5068
2|5068,5069
times|5070,5075
<EOL>|5076,5077
a|5077,5078
day|5079,5082
)|5082,5083
.|5083,5084
<EOL>|5086,5087
11.|5087,5090
fluticasone|5091,5102
-|5102,5103
salmeterol|5103,5113
250|5114,5117
-|5117,5118
50|5118,5120
mcg|5121,5124
/|5124,5125
dose|5125,5129
Disk|5130,5134
with|5135,5139
Device|5140,5146
Sig|5147,5150
:|5150,5151
<EOL>|5152,5153
One|5153,5156
(|5157,5158
1|5158,5159
)|5159,5160
Disk|5161,5165
with|5166,5170
Device|5171,5177
Inhalation|5178,5188
BID|5189,5192
(|5193,5194
2|5194,5195
times|5196,5201
a|5202,5203
day|5204,5207
)|5207,5208
.|5208,5209
<EOL>|5211,5212
12.|5212,5215
propylthiouracil|5216,5232
50|5233,5235
mg|5236,5238
Tablet|5239,5245
Sig|5246,5249
:|5249,5250
Two|5251,5254
(|5255,5256
2|5256,5257
)|5257,5258
Tablet|5259,5265
PO|5266,5268
Q8H|5269,5272
<EOL>|5273,5274
(|5274,5275
every|5275,5280
8|5281,5282
hours|5283,5288
)|5288,5289
.|5289,5290
<EOL>|5292,5293
13.|5293,5296
venlafaxine|5297,5308
75|5309,5311
mg|5312,5314
Capsule|5315,5322
,|5322,5323
Ext|5324,5327
Release|5328,5335
24|5336,5338
hr|5339,5341
Sig|5342,5345
:|5345,5346
One|5347,5350
(|5351,5352
1|5352,5353
)|5353,5354
<EOL>|5355,5356
Capsule|5356,5363
,|5363,5364
Ext|5365,5368
Release|5369,5376
24|5377,5379
hr|5380,5382
PO|5383,5385
DAILY|5386,5391
(|5392,5393
Daily|5393,5398
)|5398,5399
.|5399,5400
<EOL>|5402,5403
14.|5403,5406
venlafaxine|5407,5418
75|5419,5421
mg|5422,5424
Capsule|5425,5432
,|5432,5433
Ext|5434,5437
Release|5438,5445
24|5446,5448
hr|5449,5451
Sig|5452,5455
:|5455,5456
Two|5457,5460
(|5461,5462
2|5462,5463
)|5463,5464
<EOL>|5465,5466
Capsule|5466,5473
,|5473,5474
Ext|5475,5478
Release|5479,5486
24|5487,5489
hr|5490,5492
PO|5493,5495
DAILY|5496,5501
(|5502,5503
Daily|5503,5508
)|5508,5509
.|5509,5510
<EOL>|5512,5513
15.|5513,5516
hydrocodone|5517,5528
-|5528,5529
acetaminophen|5529,5542
_|5543,5544
_|5544,5545
_|5545,5546
mg|5547,5549
Tablet|5550,5556
Sig|5557,5560
:|5560,5561
_|5562,5563
_|5563,5564
_|5564,5565
Tablets|5566,5573
<EOL>|5574,5575
PO|5575,5577
Q8H|5578,5581
(|5582,5583
every|5583,5588
8|5589,5590
hours|5591,5596
)|5596,5597
as|5598,5600
needed|5601,5607
for|5608,5611
back|5612,5616
pain|5617,5621
.|5621,5622
<EOL>|5622,5623
Disp|5623,5627
:|5627,5628
*|5628,5629
45|5629,5631
Tablet|5632,5638
(|5638,5639
s|5639,5640
)|5640,5641
*|5641,5642
Refills|5643,5650
:|5650,5651
*|5651,5652
0|5652,5653
*|5653,5654
<EOL>|5654,5655
<EOL>|5655,5656
<EOL>|5657,5658
Discharge|5658,5667
Disposition|5668,5679
:|5679,5680
<EOL>|5680,5681
Home|5681,5685
<EOL>|5685,5686
<EOL>|5687,5688
Discharge|5688,5697
Diagnosis|5698,5707
:|5707,5708
<EOL>|5708,5709
exposure|5709,5717
of|5718,5720
craniotomy|5721,5731
hardware|5732,5740
and|5741,5744
infection|5745,5754
<EOL>|5754,5755
<EOL>|5755,5756
<EOL>|5757,5758
Mental|5779,5785
Status|5786,5792
:|5792,5793
Clear|5794,5799
and|5800,5803
coherent|5804,5812
.|5812,5813
<EOL>|5813,5814
Level|5814,5819
of|5820,5822
Consciousness|5823,5836
:|5836,5837
Alert|5838,5843
and|5844,5847
interactive|5848,5859
.|5859,5860
<EOL>|5860,5861
Activity|5861,5869
Status|5870,5876
:|5876,5877
Ambulatory|5878,5888
-|5889,5890
Independent|5891,5902
.|5902,5903
<EOL>|5903,5904
<EOL>|5904,5905
<EOL>|5906,5907
|5931,5932
Have|5932,5936
a|5937,5938
friend|5939,5945
/|5945,5946
family|5946,5952
member|5953,5959
check|5960,5965
your|5966,5970
incision|5971,5979
daily|5980,5985
for|5986,5989
<EOL>|5990,5991
signs|5991,5996
of|5997,5999
infection|6000,6009
.|6009,6010
<EOL>|6010,6011
|6011,6012
Take|6012,6016
your|6017,6021
pain|6022,6026
medicine|6027,6035
as|6036,6038
prescribed|6039,6049
.|6049,6050
<EOL>|6050,6051
|6051,6052
Exercise|6052,6060
should|6061,6067
be|6068,6070
limited|6071,6078
to|6079,6081
walking|6082,6089
;|6089,6090
no|6091,6093
lifting|6094,6101
,|6101,6102
straining|6103,6112
,|6112,6113
<EOL>|6114,6115
or|6115,6117
excessive|6118,6127
bending|6128,6135
.|6135,6136
<EOL>|6136,6137
|6137,6138
You|6138,6141
may|6142,6145
wash|6146,6150
your|6151,6155
hair|6156,6160
only|6161,6165
after|6166,6171
sutures|6172,6179
and|6180,6183
/|6183,6184
or|6184,6186
staples|6187,6194
have|6195,6199
<EOL>|6200,6201
been|6201,6205
removed|6206,6213
.|6213,6214
<EOL>|6215,6216
|6216,6217
Increase|6217,6225
your|6226,6230
intake|6231,6237
of|6238,6240
fluids|6241,6247
and|6248,6251
fiber|6252,6257
,|6257,6258
as|6259,6261
narcotic|6262,6270
pain|6271,6275
<EOL>|6276,6277
medicine|6277,6285
can|6286,6289
cause|6290,6295
constipation|6296,6308
.|6308,6309
We|6310,6312
generally|6313,6322
recommend|6323,6332
taking|6333,6339
<EOL>|6340,6341
an|6341,6343
over|6344,6348
the|6349,6352
counter|6353,6360
stool|6361,6366
softener|6367,6375
,|6375,6376
such|6377,6381
as|6382,6384
Docusate|6385,6393
(|6394,6395
Colace|6395,6401
)|6401,6402
<EOL>|6403,6404
while|6404,6409
taking|6410,6416
narcotic|6417,6425
pain|6426,6430
medication|6431,6441
.|6441,6442
<EOL>|6442,6443
|6443,6444
Unless|6444,6450
directed|6451,6459
by|6460,6462
your|6463,6467
doctor|6468,6474
,|6474,6475
do|6476,6478
not|6479,6482
take|6483,6487
any|6488,6491
<EOL>|6492,6493
anti-inflammatory|6493,6510
medicines|6511,6520
such|6521,6525
as|6526,6528
Motrin|6529,6535
,|6535,6536
Aspirin|6537,6544
,|6544,6545
Advil|6546,6551
,|6551,6552
and|6553,6556
<EOL>|6557,6558
Ibuprofen|6558,6567
etc|6568,6571
.|6571,6572
<EOL>|6573,6574
|6574,6575
Clearance|6575,6584
to|6585,6587
drive|6588,6593
and|6594,6597
return|6598,6604
to|6605,6607
work|6608,6612
will|6613,6617
be|6618,6620
addressed|6621,6630
at|6631,6633
<EOL>|6634,6635
your|6635,6639
post-operative|6640,6654
office|6655,6661
visit|6662,6667
.|6667,6668
<EOL>|6668,6669
|6669,6670
Make|6670,6674
sure|6675,6679
to|6680,6682
continue|6683,6691
to|6692,6694
use|6695,6698
your|6699,6703
incentive|6704,6713
spirometer|6714,6724
while|6725,6730
<EOL>|6731,6732
at|6732,6734
home|6735,6739
,|6739,6740
unless|6741,6747
you|6748,6751
have|6752,6756
been|6757,6761
instructed|6762,6772
not|6773,6776
to|6777,6779
.|6779,6780
<EOL>|6781,6782
<EOL>|6782,6783
CALL|6783,6787
YOUR|6788,6792
SURGEON|6793,6800
IMMEDIATELY|6801,6812
IF|6813,6815
YOU|6816,6819
EXPERIENCE|6820,6830
ANY|6831,6834
OF|6835,6837
THE|6838,6841
<EOL>|6842,6843
FOLLOWING|6843,6852
<EOL>|6852,6853
<EOL>|6853,6854
|6854,6855
New|6855,6858
onset|6859,6864
of|6865,6867
tremors|6868,6875
or|6876,6878
seizures|6879,6887
.|6887,6888
<EOL>|6888,6889
|6889,6890
Any|6890,6893
confusion|6894,6903
or|6904,6906
change|6907,6913
in|6914,6916
mental|6917,6923
status|6924,6930
.|6930,6931
<EOL>|6932,6933
|6933,6934
Any|6934,6937
numbness|6938,6946
,|6946,6947
tingling|6948,6956
,|6956,6957
weakness|6958,6966
in|6967,6969
your|6970,6974
extremities|6975,6986
.|6986,6987
<EOL>|6987,6988
|6988,6989
Pain|6989,6993
or|6994,6996
headache|6997,7005
that|7006,7010
is|7011,7013
continually|7014,7025
increasing|7026,7036
,|7036,7037
or|7038,7040
not|7041,7044
<EOL>|7045,7046
relieved|7046,7054
by|7055,7057
pain|7058,7062
medication|7063,7073
.|7073,7074
<EOL>|7074,7075
|7075,7076
Any|7076,7079
signs|7080,7085
of|7086,7088
infection|7089,7098
at|7099,7101
the|7102,7105
wound|7106,7111
site|7112,7116
:|7116,7117
redness|7118,7125
,|7125,7126
swelling|7127,7135
,|7135,7136
<EOL>|7137,7138
tenderness|7138,7148
,|7148,7149
or|7150,7152
drainage|7153,7161
.|7161,7162
<EOL>|7162,7163
|7163,7164
Fever|7164,7169
greater|7170,7177
than|7178,7182
or|7183,7185
equal|7186,7191
to|7192,7194
101|7195,7198
°|7198,7199
F|7200,7201
.|7201,7202
<EOL>|7202,7203
<EOL>|7203,7204
<EOL>|7205,7206
Followup|7206,7214
Instructions|7215,7227
:|7227,7228
<EOL>|7228,7229
_|7229,7230
_|7230,7231
_|7231,7232
<EOL>|7232,7233

