 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|32,36
No|37,39
:|39,40
_|43,44
_|44,45
_|45,46
<EOL>|46,47
<EOL>|48,49
Admission|49,58
Date|59,63
:|63,64
_|66,67
_|67,68
_|68,69
Discharge|83,92
Date|93,97
:|97,98
_|101,102
_|102,103
_|103,104
<EOL>|104,105
<EOL>|106,107
Date|107,111
of|112,114
Birth|115,120
:|120,121
_|123,124
_|124,125
_|125,126
Sex|139,142
:|142,143
F|146,147
<EOL>|147,148
<EOL>|149,150
Service|150,157
:|157,158
MEDICINE|159,167
<EOL>|167,168
<EOL>|169,170
Penicillins|182,193
/|194,195
Dilantin|196,204
_|205,206
_|206,207
_|207,208
<EOL>|208,209
<EOL>|210,211
Attending|211,220
:|220,221
_|222,223
_|223,224
_|224,225
.|225,226
<EOL>|226,227
<EOL>|228,229
diarrhea|246,254
<EOL>|254,255
<EOL>|256,257
Major|257,262
Surgical|263,271
or|272,274
Invasive|275,283
Procedure|284,293
:|293,294
<EOL>|294,295
none|295,299
<EOL>|299,300
<EOL>|300,301
<EOL>|302,303
Ms.|331,334
_|335,336
_|336,337
_|337,338
is|339,341
an|342,344
_|345,346
_|346,347
_|347,348
F|349,350
with|351,355
a|356,357
medical|358,365
history|366,373
notable|374,381
for|382,385
<EOL>|386,387
irritable|387,396
bowel|397,402
syndrome|403,411
and|412,415
dementia|416,424
.|424,425
<EOL>|426,427
<EOL>|427,428
She|428,431
reports|432,439
no|440,442
problems|443,451
with|452,456
her|457,460
bowels|461,467
for|468,471
many|472,476
years|477,482
until|483,488
the|489,492
<EOL>|493,494
acute|494,499
onset|500,505
of|506,508
diarrhea|509,517
_|518,519
_|519,520
_|520,521
morning|522,529
.|529,530
Prior|531,536
to|537,539
<EOL>|540,541
this|541,545
event|546,551
she|552,555
had|556,559
no|560,562
recent|563,569
travel|570,576
or|577,579
sick|580,584
contacts|585,593
but|594,597
did|598,601
eat|602,605
<EOL>|606,607
corned|607,613
beef|614,618
and|619,622
cabbage|623,630
at|631,633
her|634,637
local|638,643
_|644,645
_|645,646
_|646,647
hall|648,652
(|653,654
last|654,658
_|659,660
_|660,661
_|661,662
was|663,666
<EOL>|667,668
_|668,669
_|669,670
_|670,671
)|671,672
.|672,673
She|674,677
noted|678,683
nausea|684,690
with|691,695
non-bloody|696,706
,|706,707
<EOL>|708,709
non-bilious|709,720
vomitting|721,730
and|731,734
loose|735,740
watery|741,747
diarrhea|748,756
.|756,757
She|758,761
had|762,765
no|766,768
<EOL>|769,770
fever|770,775
,|775,776
abdominal|777,786
cramping|787,795
,|795,796
or|797,799
blood|800,805
in|806,808
her|809,812
stool|813,818
.|818,819
<EOL>|819,820
<EOL>|820,821
Since|821,826
that|827,831
time|832,836
her|837,840
nausea|841,847
/|847,848
vomitting|848,857
have|858,862
improved|863,871
but|872,875
her|876,879
<EOL>|880,881
diarrhea|881,889
has|890,893
not|894,897
improved|898,906
despite|907,914
Imodium|915,922
.|922,923
She|924,927
was|928,931
unable|932,938
to|939,941
<EOL>|942,943
keep|943,947
down|948,952
oral|953,957
foods|958,963
and|964,967
presented|968,977
to|978,980
the|981,984
ED|985,987
today|988,993
.|993,994
<EOL>|995,996
<EOL>|996,997
Vital|997,1002
signs|1003,1008
on|1009,1011
arrival|1012,1019
to|1020,1022
_|1023,1024
_|1024,1025
_|1025,1026
ED|1027,1029
:|1029,1030
T|1031,1032
97.6|1033,1037
,|1037,1038
P|1039,1040
97|1041,1043
,|1043,1044
BP|1045,1047
167|1048,1051
/|1051,1052
81|1052,1054
,|1054,1055
<EOL>|1056,1057
100|1057,1060
%|1060,1061
on|1062,1064
RA|1065,1067
.|1067,1068
Her|1069,1072
evaluation|1073,1083
in|1084,1086
the|1087,1090
ED|1091,1093
was|1094,1097
notable|1098,1105
for|1106,1109
guaiac|1110,1116
<EOL>|1117,1118
positive|1118,1126
stool|1127,1132
,|1132,1133
a|1134,1135
WBC|1136,1139
count|1140,1145
of|1146,1148
4.1|1149,1152
,|1152,1153
and|1154,1157
an|1158,1160
elevated|1161,1169
BUN|1170,1173
to|1174,1176
33|1177,1179
.|1179,1180
<EOL>|1181,1182
In|1182,1184
the|1185,1188
ED|1189,1191
she|1192,1195
received|1196,1204
1|1205,1206
liter|1207,1212
of|1213,1215
normal|1216,1222
saline|1223,1229
.|1229,1230
<EOL>|1230,1231
<EOL>|1231,1232
Review|1232,1238
of|1239,1241
Systems|1242,1249
:|1249,1250
Pain|1251,1255
assessment|1256,1266
on|1267,1269
arrival|1270,1277
to|1278,1280
the|1281,1284
floor|1285,1290
:|1290,1291
_|1292,1293
_|1293,1294
_|1294,1295
<EOL>|1296,1297
(|1297,1298
no|1298,1300
pain|1301,1305
)|1305,1306
.|1306,1307
No|1308,1310
recent|1311,1317
illnesses|1318,1327
.|1327,1328
No|1329,1331
fevers|1332,1338
,|1338,1339
chills|1340,1346
,|1346,1347
or|1348,1350
night|1351,1356
<EOL>|1357,1358
sweats|1358,1364
.|1364,1365
No|1366,1368
SOB|1369,1372
,|1372,1373
cough|1374,1379
,|1379,1380
or|1381,1383
chest|1384,1389
pain|1390,1394
.|1394,1395
No|1396,1398
urinary|1399,1406
symptoms|1407,1415
.|1415,1416
Other|1417,1422
<EOL>|1423,1424
systems|1424,1431
reviewed|1432,1440
in|1441,1443
detail|1444,1450
and|1451,1454
all|1455,1458
otherwise|1459,1468
negative|1469,1477
.|1477,1478
<EOL>|1478,1479
<EOL>|1480,1481
Hypertension|1503,1515
<EOL>|1515,1516
Dementia|1516,1524
<EOL>|1524,1525
Osteoporosis|1525,1537
<EOL>|1537,1538
Irritable|1538,1547
bowel|1548,1553
syndrome|1554,1562
<EOL>|1562,1563
Macrocytosis|1563,1575
of|1576,1578
unclear|1579,1586
etiology|1587,1595
<EOL>|1595,1596
Left|1596,1600
ear|1601,1604
hearing|1605,1612
loss|1613,1617
<EOL>|1617,1618
Status|1618,1624
post|1625,1629
hysterectomy|1630,1642
<EOL>|1642,1643
Status|1643,1649
post|1650,1654
appendectomy|1655,1667
<EOL>|1667,1668
Status|1668,1674
post|1675,1679
ovarian|1680,1687
cyst|1688,1692
removal|1693,1700
<EOL>|1700,1701
Cataract|1701,1709
surgery|1710,1717
<EOL>|1717,1718
Glaucoma|1718,1726
<EOL>|1726,1727
<EOL>|1728,1729
:|1743,1744
<EOL>|1744,1745
_|1745,1746
_|1746,1747
_|1747,1748
<EOL>|1748,1749
:|1763,1764
<EOL>|1764,1765
Not|1765,1768
relevant|1769,1777
to|1778,1780
the|1781,1784
current|1785,1792
admission|1793,1802
.|1802,1803
<EOL>|1803,1804
<EOL>|1805,1806
Vital|1821,1826
Signs|1827,1832
:|1832,1833
T|1834,1835
98.6|1836,1840
,|1840,1841
P|1842,1843
64|1844,1846
,|1846,1847
BP|1848,1850
124|1851,1854
/|1854,1855
72|1855,1857
,|1857,1858
95|1859,1861
%|1861,1862
on|1863,1865
RA|1866,1868
.|1868,1869
<EOL>|1869,1870
<EOL>|1870,1871
-|1893,1894
Gen|1895,1898
:|1898,1899
Elderly|1900,1907
female|1908,1914
sitting|1915,1922
up|1923,1925
in|1926,1928
bed|1929,1932
in|1933,1935
NAD|1936,1939
.|1939,1940
<EOL>|1940,1941
-|1941,1942
HEENT|1943,1948
:|1948,1949
Hard|1950,1954
of|1955,1957
hearing|1958,1965
.|1965,1966
Right|1967,1972
ear|1973,1976
better|1977,1983
than|1984,1988
left|1989,1993
.|1993,1994
<EOL>|1994,1995
-|1995,1996
Chest|1997,2002
:|2002,2003
Normal|2004,2010
respirations|2011,2023
and|2024,2027
breathing|2028,2037
comfortably|2038,2049
on|2050,2052
room|2053,2057
<EOL>|2058,2059
air.|2059,2063
Lungs|2064,2069
clear|2070,2075
to|2076,2078
auscultation|2079,2091
bilaterally|2092,2103
.|2103,2104
<EOL>|2104,2105
-|2105,2106
CV|2107,2109
:|2109,2110
Regular|2111,2118
rhythm|2119,2125
.|2125,2126
Normal|2127,2133
S1|2134,2136
,|2136,2137
S2|2138,2140
.|2140,2141
No|2142,2144
murmurs|2145,2152
or|2153,2155
gallops|2156,2163
.|2163,2164
JVP|2165,2168
<EOL>|2169,2170
<|2170,2171
5|2171,2172
cm|2173,2175
.|2175,2176
<EOL>|2177,2178
-|2178,2179
Abdomen|2180,2187
:|2187,2188
Normal|2189,2195
bowel|2196,2201
sounds|2202,2208
.|2208,2209
Soft|2210,2214
,|2214,2215
nontender|2216,2225
,|2225,2226
nondistended|2227,2239
.|2239,2240
<EOL>|2241,2242
-|2242,2243
Extremities|2244,2255
:|2255,2256
No|2257,2259
ankle|2260,2265
edema|2266,2271
.|2271,2272
<EOL>|2272,2273
-|2273,2274
Neuro|2275,2280
:|2280,2281
Alert|2282,2287
,|2287,2288
oriented|2289,2297
x|2298,2299
_|2300,2301
_|2301,2302
_|2302,2303
.|2303,2304
Most|2305,2309
of|2310,2312
history|2313,2320
aided|2321,2326
by|2327,2329
<EOL>|2330,2331
daughter|2331,2339
.|2339,2340
Does|2341,2345
not|2346,2349
know|2350,2354
home|2355,2359
medications|2360,2371
or|2372,2374
specifics|2375,2384
timing|2385,2391
of|2392,2394
<EOL>|2395,2396
recent|2396,2402
events|2403,2409
.|2409,2410
Has|2411,2414
short|2415,2420
-|2420,2421
term|2421,2425
memory|2426,2432
impairment|2433,2443
.|2443,2444
Speech|2445,2451
and|2452,2455
<EOL>|2456,2457
language|2457,2465
are|2466,2469
normal|2470,2476
.|2476,2477
<EOL>|2478,2479
-|2479,2480
Psych|2481,2486
:|2486,2487
Appearance|2488,2498
,|2498,2499
behavior|2500,2508
,|2508,2509
and|2510,2513
affect|2514,2520
all|2521,2524
normal|2525,2531
.|2531,2532
<EOL>|2532,2533
<EOL>|2533,2534
<EOL>|2535,2536
Pertinent|2536,2545
Results|2546,2553
:|2553,2554
<EOL>|2554,2555
Admission|2555,2564
Labs|2565,2569
:|2569,2570
<EOL>|2570,2571
_|2571,2572
_|2572,2573
_|2573,2574
09|2575,2577
:|2577,2578
35AM|2578,2582
BLOOD|2583,2588
WBC|2589,2592
-|2592,2593
4.1|2593,2596
(|2597,2598
Neuts|2598,2603
-|2603,2604
58|2604,2606
Bands|2607,2612
-|2612,2613
2|2613,2614
Lymphs|2615,2621
-|2621,2622
24|2622,2624
<EOL>|2625,2626
Monos|2626,2631
-|2631,2632
15|2632,2634
*|2634,2635
Eos|2636,2639
-|2639,2640
0|2640,2641
Baso|2642,2646
-|2646,2647
1|2647,2648
_|2649,2650
_|2650,2651
_|2651,2652
Myelos|2653,2659
-|2659,2660
0|2660,2661
)|2661,2662
RBC|2663,2666
-|2666,2667
4|2667,2668
.|2668,2669
40|2669,2671
<EOL>|2672,2673
Hgb|2673,2676
-|2676,2677
14.9|2677,2681
Hct|2682,2685
-|2685,2686
43.5|2686,2690
MCV|2691,2694
-|2694,2695
99|2695,2697
*|2697,2698
MCH|2699,2702
-|2702,2703
33|2703,2705
.|2705,2706
8|2706,2707
*|2707,2708
MCHC|2709,2713
-|2713,2714
34.2|2714,2718
RDW|2719,2722
-|2722,2723
13.2|2723,2727
Plt|2728,2731
<EOL>|2732,2733
_|2733,2734
_|2734,2735
_|2735,2736
<EOL>|2736,2737
_|2737,2738
_|2738,2739
_|2739,2740
09|2741,2743
:|2743,2744
35AM|2744,2748
BLOOD|2749,2754
Glucose|2755,2762
-|2762,2763
118|2763,2766
*|2766,2767
UreaN|2768,2773
-|2773,2774
33|2774,2776
*|2776,2777
Creat|2778,2783
-|2783,2784
1.1|2784,2787
Na|2788,2790
-|2790,2791
144|2791,2794
<EOL>|2795,2796
K|2796,2797
-|2797,2798
3.4|2798,2801
Cl|2802,2804
-|2804,2805
107|2805,2808
HCO3|2809,2813
-|2813,2814
21|2814,2816
*|2816,2817
AnGap|2818,2823
-|2823,2824
19|2824,2826
ALT|2827,2830
-|2830,2831
21|2831,2833
AST|2834,2837
-|2837,2838
22|2838,2840
AlkPhos|2841,2848
-|2848,2849
53|2849,2851
<EOL>|2852,2853
TotBili|2853,2860
-|2860,2861
0.6|2861,2864
Lipase|2865,2871
-|2871,2872
16|2872,2874
Albumin|2875,2882
-|2882,2883
4.6|2883,2886
<EOL>|2886,2887
-|2888,2889
_|2890,2891
_|2891,2892
_|2892,2893
10|2894,2896
:|2896,2897
30AM|2897,2901
URINE|2902,2907
Color|2908,2913
-|2913,2914
Yellow|2914,2920
Appear|2921,2927
-|2927,2928
Hazy|2928,2932
Sp|2933,2935
_|2936,2937
_|2937,2938
_|2938,2939
<EOL>|2940,2941
Blood|2941,2946
-|2946,2947
NEG|2947,2950
Nitrite|2951,2958
-|2958,2959
NEG|2959,2962
Protein|2963,2970
-|2970,2971
30|2971,2973
Glucose|2974,2981
-|2981,2982
NEG|2982,2985
Ketone|2986,2992
-|2992,2993
NEG|2993,2996
<EOL>|2997,2998
Bilirub|2998,3005
-|3005,3006
NEG|3006,3009
Urobiln|3010,3017
-|3017,3018
NEG|3018,3021
pH|3022,3024
-|3024,3025
6.0|3025,3028
Leuks|3029,3034
-|3034,3035
NEG|3035,3038
RBC|3039,3042
-|3042,3043
1|3043,3044
WBC|3045,3048
-|3048,3049
4|3049,3050
Bacteri|3051,3058
-|3058,3059
MOD|3059,3062
<EOL>|3063,3064
Yeast|3064,3069
-|3069,3070
NONE|3070,3074
Epi|3075,3078
-|3078,3079
0|3079,3080
CastGr|3081,3087
-|3087,3088
7|3088,3089
*|3089,3090
CastHy|3091,3097
-|3097,3098
93|3098,3100
*|3100,3101
CastCel|3102,3109
-|3109,3110
1|3110,3111
*|3111,3112
<EOL>|3112,3113
.|3113,3114
<EOL>|3114,3115
Microbiology|3115,3127
:|3127,3128
<EOL>|3128,3129
_|3129,3130
_|3130,3131
_|3131,3132
Stool|3133,3138
Cultures|3139,3147
:|3147,3148
<EOL>|3148,3149
_|3149,3150
_|3150,3151
_|3151,3152
9|3153,3154
:|3154,3155
58|3155,3157
pm|3158,3160
STOOL|3161,3166
CONSISTENCY|3171,3182
:|3182,3183
WATERY|3184,3190
Source|3196,3202
:|3202,3203
<EOL>|3204,3205
Stool|3205,3210
.|3210,3211
<EOL>|3212,3213
FECAL|3216,3221
CULTURE|3222,3229
(|3230,3231
Pending|3231,3238
)|3238,3239
:|3239,3240
<EOL>|3241,3242
CAMPYLOBACTER|3245,3258
CULTURE|3259,3266
(|3267,3268
Pending|3268,3275
)|3275,3276
:|3276,3277
<EOL>|3278,3279
CLOSTRIDIUM|3282,3293
DIFFICILE|3294,3303
TOXIN|3304,3309
A|3310,3311
&|3312,3313
B|3314,3315
TEST|3316,3320
(|3321,3322
Final|3322,3327
_|3328,3329
_|3329,3330
_|3330,3331
:|3331,3332
<EOL>|3333,3334
Feces|3340,3345
negative|3346,3354
for|3355,3358
C|3359,3360
.|3360,3361
difficile|3361,3370
toxin|3371,3376
A|3377,3378
&|3379,3380
B|3381,3382
by|3383,3385
EIA|3386,3389
.|3389,3390
<EOL>|3391,3392
(|3403,3404
Reference|3404,3413
Range|3414,3419
-|3419,3420
Negative|3420,3428
)|3428,3429
.|3429,3430
<EOL>|3431,3432
.|3432,3433
<EOL>|3433,3434
_|3434,3435
_|3435,3436
_|3436,3437
Urine|3438,3443
Cultures|3444,3452
NGTD|3453,3457
<EOL>|3457,3458
_|3458,3459
_|3459,3460
_|3460,3461
06|3462,3464
:|3464,3465
47AM|3465,3469
BLOOD|3470,3475
WBC|3476,3479
-|3479,3480
6|3480,3481
.|3481,3482
6|3482,3483
#|3483,3484
RBC|3485,3488
-|3488,3489
3|3489,3490
.|3490,3491
72|3491,3493
*|3493,3494
Hgb|3495,3498
-|3498,3499
12.3|3499,3503
Hct|3504,3507
-|3507,3508
36.5|3508,3512
<EOL>|3513,3514
MCV|3514,3517
-|3517,3518
98|3518,3520
MCH|3521,3524
-|3524,3525
33|3525,3527
.|3527,3528
2|3528,3529
*|3529,3530
MCHC|3531,3535
-|3535,3536
33.8|3536,3540
RDW|3541,3544
-|3544,3545
12.6|3545,3549
Plt|3550,3553
_|3554,3555
_|3555,3556
_|3556,3557
<EOL>|3557,3558
_|3558,3559
_|3559,3560
_|3560,3561
06|3562,3564
:|3564,3565
47AM|3565,3569
BLOOD|3570,3575
Glucose|3576,3583
-|3583,3584
93|3584,3586
UreaN|3587,3592
-|3592,3593
12|3593,3595
Creat|3596,3601
-|3601,3602
0.7|3602,3605
Na|3606,3608
-|3608,3609
143|3609,3612
<EOL>|3613,3614
K|3614,3615
-|3615,3616
3.7|3616,3619
Cl|3620,3622
-|3622,3623
109|3623,3626
*|3626,3627
HCO3|3628,3632
-|3632,3633
28|3633,3635
AnGap|3636,3641
-|3641,3642
10|3642,3644
<EOL>|3644,3645
_|3645,3646
_|3646,3647
_|3647,3648
09|3649,3651
:|3651,3652
35AM|3652,3656
BLOOD|3657,3662
ALT|3663,3666
-|3666,3667
21|3667,3669
AST|3670,3673
-|3673,3674
22|3674,3676
AlkPhos|3677,3684
-|3684,3685
53|3685,3687
TotBili|3688,3695
-|3695,3696
0.6|3696,3699
<EOL>|3699,3700
_|3700,3701
_|3701,3702
_|3702,3703
09|3704,3706
:|3706,3707
35AM|3707,3711
BLOOD|3712,3717
cTropnT|3718,3725
-|3725,3726
<|3726,3727
0|3727,3728
.|3728,3729
01|3729,3731
<EOL>|3731,3732
_|3732,3733
_|3733,3734
_|3734,3735
06|3736,3738
:|3738,3739
47AM|3739,3743
BLOOD|3744,3749
Calcium|3750,3757
-|3757,3758
8|3758,3759
.|3759,3760
2|3760,3761
*|3761,3762
Phos|3763,3767
-|3767,3768
2|3768,3769
.|3769,3770
4|3770,3771
*|3771,3772
Mg|3773,3775
-|3775,3776
1.|3776,3778
_|3778,3779
_|3779,3780
_|3780,3781
y|3782,3783
/|3783,3784
o|3784,3785
F|3786,3787
with|3788,3792
PMhx|3793,3797
of|3798,3800
IBS|3801,3804
and|3805,3808
Dementia|3809,3817
who|3818,3821
presented|3822,3831
with|3832,3836
_|3837,3838
_|3838,3839
_|3839,3840
<EOL>|3841,3842
days|3842,3846
of|3847,3849
nausea|3850,3856
,|3856,3857
vomiting|3858,3866
and|3867,3870
non-bloody|3871,3881
diarrhea|3882,3890
.|3890,3891
Pt|3892,3894
was|3895,3898
notably|3899,3906
<EOL>|3907,3908
dehydrated|3908,3918
on|3919,3921
admission|3922,3931
with|3932,3936
acute|3937,3942
renal|3943,3948
failure|3949,3956
and|3957,3960
symptomatic|3961,3972
<EOL>|3973,3974
orthostasis|3974,3985
.|3985,3986
She|3987,3990
was|3991,3994
treated|3995,4002
with|4003,4007
IVF|4008,4011
and|4012,4015
bowel|4016,4021
rest|4022,4026
.|4026,4027
<EOL>|4029,4030
Infectious|4030,4040
work|4041,4045
up|4046,4048
including|4049,4058
Cdiff|4059,4064
returned|4065,4073
negative|4074,4082
and|4083,4086
<EOL>|4087,4088
presentation|4088,4100
was|4101,4104
most|4105,4109
consistent|4110,4120
with|4121,4125
norovirus|4126,4135
.|4135,4136
Pt|4138,4140
was|4141,4144
slowly|4145,4151
<EOL>|4152,4153
advanced|4153,4161
a|4162,4163
diet|4164,4168
and|4169,4172
diarrhea|4173,4181
improved|4182,4190
.|4190,4191
Renal|4193,4198
function|4199,4207
returned|4208,4216
<EOL>|4217,4218
to|4218,4220
baseline|4221,4229
with|4230,4234
IVF|4235,4238
and|4239,4242
pt|4243,4245
was|4246,4249
tolerating|4250,4260
a|4261,4262
bland|4263,4268
diet|4269,4273
without|4274,4281
<EOL>|4282,4283
any|4283,4286
evidence|4287,4295
of|4296,4298
orthostasis|4299,4310
by|4311,4313
the|4314,4317
day|4318,4321
of|4322,4324
discharge|4325,4334
.|4334,4335
Pt|4337,4339
was|4340,4343
<EOL>|4344,4345
seen|4345,4349
by|4350,4352
_|4353,4354
_|4354,4355
_|4355,4356
who|4357,4360
felt|4361,4365
that|4366,4370
she|4371,4374
was|4375,4378
safe|4379,4383
for|4384,4387
discharge|4388,4397
home|4398,4402
without|4403,4410
<EOL>|4411,4412
services|4412,4420
.|4420,4421
<EOL>|4423,4424
.|4424,4425
<EOL>|4425,4426
Conjunctivitis|4426,4440
(|4441,4442
left|4442,4446
eye|4447,4450
)|4450,4451
:|4451,4452
At|4453,4455
the|4456,4459
time|4460,4464
of|4465,4467
admission|4468,4477
,|4477,4478
pt|4479,4481
reported|4482,4490
<EOL>|4491,4492
being|4492,4497
treated|4498,4505
with|4506,4510
azithromycin|4511,4523
drops|4524,4529
for|4530,4533
left|4534,4538
eye|4539,4542
<EOL>|4543,4544
conjunctivitis|4544,4558
but|4559,4562
was|4563,4566
having|4567,4573
ongoing|4574,4581
symptoms|4582,4590
.|4590,4591
Pt|4592,4594
was|4595,4598
started|4599,4606
<EOL>|4607,4608
on|4608,4610
erythromycin|4611,4623
opthalmic|4624,4633
ointment|4634,4642
with|4643,4647
some|4648,4652
improvement|4653,4664
in|4665,4667
<EOL>|4668,4669
conjunctival|4669,4681
injection|4682,4691
.|4691,4692
She|4694,4697
was|4698,4701
instructed|4702,4712
to|4713,4715
monitor|4716,4723
for|4724,4727
any|4728,4731
<EOL>|4732,4733
worsening|4733,4742
in|4743,4745
eye|4746,4749
symptoms|4750,4758
and|4759,4762
was|4763,4766
scheduled|4767,4776
for|4777,4780
follow|4781,4787
up|4788,4790
with|4791,4795
<EOL>|4796,4797
her|4797,4800
PCP|4801,4804
.|4804,4805
<EOL>|4805,4806
.|4806,4807
<EOL>|4807,4808
Otherwise|4808,4817
,|4817,4818
there|4819,4824
were|4825,4829
no|4830,4832
changes|4833,4840
made|4841,4845
to|4846,4848
her|4849,4852
chronic|4853,4860
medication|4861,4871
<EOL>|4872,4873
regimen|4873,4880
<EOL>|4881,4882
.|4882,4883
<EOL>|4883,4884
Code|4884,4888
Status|4889,4895
:|4895,4896
DNR|4897,4900
/|4900,4901
DNI|4901,4904
confirmed|4905,4914
on|4915,4917
admission|4918,4927
with|4928,4932
patient|4933,4940
and|4941,4944
her|4945,4948
<EOL>|4949,4950
HCP|4950,4953
.|4953,4954
<EOL>|4954,4955
<EOL>|4955,4956
<EOL>|4957,4958
Medications|4958,4969
on|4970,4972
Admission|4973,4982
:|4982,4983
<EOL>|4983,4984
-|4984,4985
list|4985,4989
confirmed|4990,4999
with|5000,5004
primary|5005,5012
caregiver|5013,5022
on|5023,5025
admission|5026,5035
-|5035,5036
<EOL>|5036,5037
_|5037,5038
_|5038,5039
_|5039,5040
10|5041,5043
mg|5044,5046
daily|5047,5052
<EOL>|5053,5054
Namenda|5054,5061
10|5062,5064
mg|5065,5067
daily|5068,5073
<EOL>|5073,5074
Aspirin|5074,5081
162|5082,5085
.|5085,5086
5|5086,5087
mg|5088,5090
daily|5091,5096
<EOL>|5100,5101
Raloxifene|5101,5111
(|5112,5113
Evista|5113,5119
)|5119,5120
60|5121,5123
mg|5124,5126
daily|5127,5132
<EOL>|5135,5136
Multivitamin|5136,5148
daily|5149,5154
<EOL>|5154,5155
Glucosamine|5155,5166
<EOL>|5170,5171
Calcium|5171,5178
supplement|5179,5189
<EOL>|5189,5190
Cholecalciferol|5190,5205
(|5206,5207
Vitamin|5207,5214
D3|5215,5217
)|5217,5218
1,000|5219,5224
units|5225,5230
daily|5231,5236
<EOL>|5239,5240
Ascorbic|5240,5248
Acid|5249,5253
SR|5254,5256
500|5257,5260
mg|5261,5263
daily|5264,5269
<EOL>|5269,5270
<EOL>|5271,5272
Discharge|5272,5281
Medications|5282,5293
:|5293,5294
<EOL>|5294,5295
1.|5295,5297
donepezil|5298,5307
5|5308,5309
mg|5310,5312
Tablet|5313,5319
Sig|5320,5323
:|5323,5324
Two|5325,5328
(|5329,5330
2|5330,5331
)|5331,5332
Tablet|5333,5339
PO|5340,5342
HS|5343,5345
(|5346,5347
at|5347,5349
bedtime|5350,5357
)|5357,5358
.|5358,5359
<EOL>|5360,5361
<EOL>|5362,5363
2.|5363,5365
Namenda|5366,5373
10|5374,5376
mg|5377,5379
Tablet|5380,5386
Sig|5387,5390
:|5390,5391
One|5392,5395
(|5396,5397
1|5397,5398
)|5398,5399
Tablet|5400,5406
PO|5407,5409
qhs|5410,5413
(|5414,5415
)|5415,5416
.|5416,5417
<EOL>|5419,5420
3.|5420,5422
aspirin|5423,5430
162|5431,5434
mg|5435,5437
Tablet|5438,5444
,|5444,5445
Delayed|5446,5453
Release|5454,5461
(|5462,5463
E.C|5463,5466
.|5466,5467
)|5467,5468
Sig|5469,5472
:|5472,5473
One|5474,5477
(|5478,5479
1|5479,5480
)|5480,5481
<EOL>|5482,5483
Tablet|5483,5489
,|5489,5490
Delayed|5491,5498
Release|5499,5506
(|5507,5508
E.C|5508,5511
.|5511,5512
)|5512,5513
PO|5514,5516
once|5517,5521
a|5522,5523
day|5524,5527
.|5527,5528
<EOL>|5530,5531
4.|5531,5533
raloxifene|5534,5544
60|5545,5547
mg|5548,5550
Tablet|5551,5557
Sig|5558,5561
:|5561,5562
One|5563,5566
(|5567,5568
1|5568,5569
)|5569,5570
Tablet|5571,5577
PO|5578,5580
once|5581,5585
a|5586,5587
week|5588,5592
.|5592,5593
<EOL>|5595,5596
5.|5596,5598
multivitamin|5599,5611
Oral|5613,5617
<EOL>|5617,5618
6.|5618,5620
Glucosamine|5621,5632
Oral|5634,5638
<EOL>|5638,5639
7.|5639,5641
Vitamin|5642,5649
D|5650,5651
Oral|5653,5657
<EOL>|5657,5658
8.|5658,5660
ascorbic|5661,5669
acid|5670,5674
Oral|5676,5680
<EOL>|5680,5681
9.|5681,5683
Calcium|5684,5691
500|5692,5695
Oral|5697,5701
<EOL>|5701,5702
10.|5702,5705
erythromycin|5706,5718
5|5719,5720
mg|5721,5723
/|5723,5724
gram|5724,5728
(|5729,5730
0.5|5730,5733
%|5734,5735
)|5735,5736
Ointment|5737,5745
Sig|5746,5749
:|5749,5750
0.5|5751,5754
inch|5755,5759
<EOL>|5760,5761
Ophthalmic|5761,5771
four|5772,5776
times|5777,5782
a|5783,5784
day|5785,5788
for|5789,5792
5|5793,5794
days|5795,5799
:|5799,5800
apply|5801,5806
to|5807,5809
left|5810,5814
eye|5815,5818
for|5820,5823
<EOL>|5824,5825
another|5825,5832
5|5833,5834
days|5835,5839
.|5840,5841
<EOL>|5841,5842
Disp|5842,5846
:|5846,5847
*|5847,5848
qs|5848,5850
tube|5851,5855
*|5855,5856
Refills|5857,5864
:|5864,5865
*|5865,5866
0|5866,5867
*|5867,5868
<EOL>|5868,5869
<EOL>|5869,5870
<EOL>|5871,5872
Discharge|5872,5881
Disposition|5882,5893
:|5893,5894
<EOL>|5894,5895
Home|5895,5899
<EOL>|5899,5900
<EOL>|5901,5902
Discharge|5902,5911
Diagnosis|5912,5921
:|5921,5922
<EOL>|5922,5923
Primary|5923,5930
:|5930,5931
<EOL>|5932,5933
Gastrointestinal|5933,5949
Virus|5950,5955
<EOL>|5955,5956
Dehydration|5956,5967
<EOL>|5968,5969
Symptomatic|5969,5980
orthostasis|5981,5992
<EOL>|5992,5993
<EOL>|5993,5994
<EOL>|5995,5996
Mental|6017,6023
Status|6024,6030
:|6030,6031
Clear|6032,6037
and|6038,6041
coherent|6042,6050
.|6050,6051
<EOL>|6051,6052
Level|6052,6057
of|6058,6060
Consciousness|6061,6074
:|6074,6075
Alert|6076,6081
and|6082,6085
interactive|6086,6097
.|6097,6098
<EOL>|6098,6099
Activity|6099,6107
Status|6108,6114
:|6114,6115
Ambulatory|6116,6126
-|6127,6128
Independent|6129,6140
.|6140,6141
<EOL>|6141,6142
<EOL>|6142,6143
<EOL>|6144,6145
You|6169,6172
were|6173,6177
admitted|6178,6186
with|6187,6191
an|6192,6194
acute|6195,6200
diarrheal|6201,6210
illness|6211,6218
and|6219,6222
<EOL>|6223,6224
dehydration|6224,6235
.|6235,6236
This|6238,6242
was|6243,6246
likely|6247,6253
due|6254,6257
to|6258,6260
a|6261,6262
virus|6263,6268
which|6269,6274
can|6275,6278
be|6279,6281
very|6282,6286
<EOL>|6287,6288
contagious|6288,6298
.|6298,6299
You|6301,6304
have|6305,6309
been|6310,6314
treated|6315,6322
with|6323,6327
IV|6328,6330
fluids|6331,6337
and|6338,6341
supportive|6342,6352
<EOL>|6353,6354
care|6354,6358
with|6359,6363
improvement|6364,6375
in|6376,6378
your|6379,6383
symptoms|6384,6392
.|6392,6393
You|6395,6398
have|6399,6403
been|6404,6408
seen|6409,6413
by|6414,6416
<EOL>|6417,6418
physical|6418,6426
therapy|6427,6434
who|6435,6438
agree|6439,6444
that|6445,6449
you|6450,6453
are|6454,6457
safe|6458,6462
to|6463,6465
return|6466,6472
home|6473,6477
<EOL>|6478,6479
today|6479,6484
.|6484,6485
We|6487,6489
encourage|6490,6499
you|6500,6503
take|6504,6508
as|6509,6511
much|6512,6516
oral|6517,6521
hydration|6522,6531
as|6532,6534
possible|6535,6543
<EOL>|6544,6545
and|6545,6548
continue|6549,6557
advancing|6558,6567
your|6568,6572
diet|6573,6577
as|6578,6580
tolerated|6581,6590
.|6590,6591
Please|6593,6599
keep|6600,6604
your|6605,6609
<EOL>|6610,6611
appointment|6611,6622
with|6623,6627
Dr.|6628,6631
_|6632,6633
_|6633,6634
_|6634,6635
on|6636,6638
_|6639,6640
_|6640,6641
_|6641,6642
.|6642,6643
<EOL>|6643,6644
.|6644,6645
<EOL>|6645,6646
We|6646,6648
have|6649,6653
given|6654,6659
you|6660,6663
a|6664,6665
new|6666,6669
prescription|6670,6682
to|6683,6685
help|6686,6690
treat|6691,6696
the|6697,6700
left|6701,6705
eye|6706,6709
<EOL>|6710,6711
conjunctivitis|6711,6725
,|6725,6726
please|6727,6733
continue|6734,6742
using|6743,6748
the|6749,6752
erythromycin|6753,6765
ointment|6766,6774
<EOL>|6775,6776
for|6776,6779
another|6780,6787
5|6788,6789
days|6790,6794
.|6794,6795
If|6797,6799
you|6800,6803
develop|6804,6811
any|6812,6815
rash|6816,6820
on|6821,6823
your|6824,6828
face|6829,6833
,|6833,6834
<EOL>|6835,6836
fevers|6836,6842
,|6842,6843
visual|6844,6850
changes|6851,6858
or|6859,6861
worsening|6862,6871
in|6872,6874
eye|6875,6878
symptoms|6879,6887
,|6887,6888
please|6889,6895
call|6896,6900
<EOL>|6901,6902
your|6902,6906
PCP|6907,6910
or|6911,6913
return|6914,6920
for|6921,6924
urgent|6925,6931
evaluation|6932,6942
.|6942,6943
<EOL>|6943,6944
.|6944,6945
<EOL>|6945,6946
Otherwise|6946,6955
,|6955,6956
we|6957,6959
have|6960,6964
not|6965,6968
made|6969,6973
any|6974,6977
changes|6978,6985
to|6986,6988
your|6989,6993
medications|6994,7005
<EOL>|7005,7006
<EOL>|7007,7008
Followup|7008,7016
Instructions|7017,7029
:|7029,7030
<EOL>|7030,7031
_|7031,7032
_|7032,7033
_|7033,7034
<EOL>|7034,7035

