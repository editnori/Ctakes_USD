CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Known|Modifier|false|false||Knownnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Adverse reaction to drug|Finding|true|false||Adverse Drug Reactionsnull|Adverse reaction to drug|Finding|true|false||Drug Reactionsnull|Pharmaceutical Preparations|Drug|false|false||Drug
null|Pharmacologic Substance|Drug|false|false||Drugnull|Drug problem|Finding|false|false||Drugnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Chief complaint (finding)|Finding|false|false||Chief Complaintnull|Complaint (finding)|Finding|false|false||Complaintnull|null|Attribute|false|false||Complaintnull|Atypical chest pain|Finding|false|false|C1527391;C0817096|Atypical chest painnull|atypia morphology|Finding|false|false||Atypicalnull|Atypical|Modifier|false|false||Atypicalnull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0262384;C0008031;C2926613;C1549543;C0030193;C0741025|chest
null|Anterior thoracic region|Anatomy|false|false|C0262384;C0008031;C2926613;C1549543;C0030193;C0741025|chestnull|Administration Method - Pain|Finding|false|false|C1527391;C0817096|pain
null|Pain|Finding|false|false|C1527391;C0817096|painnull|null|Attribute|false|false||painnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|ECHO protocol|Procedure|false|false||Echo
null|Extension for Community Healthcare Outcomes|Procedure|false|false||Echonull|Echo <Calopterygidae>|Entity|false|false||Echonull|History of present illness (finding)|Finding|false|false||History of Present Illnessnull|null|Attribute|false|false||History of Present Illnessnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Present illness|Finding|false|false||Present Illnessnull|Present|Finding|false|false||Present
null|Presentation|Finding|false|false||Presentnull|Illness (finding)|Finding|false|false||Illnessnull|Woman|Subject|false|false||woman
null|Human, Female adult|Subject|false|false||womannull|Intermittent|Time|false|false||intermittentnull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C2926613;C0008031;C0741025|chest
null|Anterior thoracic region|Anatomy|false|false|C2926613;C0008031;C0741025|chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Several|LabModifier|false|false||severalnull|month|Time|false|false||monthsnull|Administration Method - Pain|Finding|false|false|C0037004;C4299050|Pain
null|Pain|Finding|false|false|C0037004;C4299050|Painnull|null|Attribute|false|false||Painnull|Left posterior|Modifier|false|false||left posteriornull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Posterior pituitary disease|Disorder|false|false||posteriornull|Dorsal|Modifier|false|false||posteriornull|Procedures on Shoulder|Procedure|false|false|C0037004;C4299050|shoulder
null|Examination of shoulder(s)|Procedure|false|false|C0037004;C4299050|shouldernull|Upper extremity>Shoulder|Anatomy|false|false|C1549543;C0030193;C0869975;C0221590|shoulder
null|Shoulder|Anatomy|false|false|C1549543;C0030193;C0869975;C0221590|shouldernull|Anorectal Malformations|Disorder|false|false|C0446516;C1140618;C1269078|armnull|AKR1A1 wt Allele|Finding|false|false|C0446516;C1140618;C1269078|arm
null|ARMC9 gene|Finding|false|false|C0446516;C1140618;C1269078|armnull|Protocol Treatment Arm|Procedure|false|false|C0446516;C1140618;C1269078|arm
null|Axillary Reverse Mapping|Procedure|false|false|C0446516;C1140618;C1269078|arm
null|Study Arm|Procedure|false|false|C0446516;C1140618;C1269078|armnull|Upper arm|Anatomy|false|false|C3495676;C1522541;C5400986;C4761640;C1824218;C3715044|arm
null|null|Anatomy|false|false|C3495676;C1522541;C5400986;C4761640;C1824218;C3715044|arm
null|Upper Extremity|Anatomy|false|false|C3495676;C1522541;C5400986;C4761640;C1824218;C3715044|armnull|Fingers|Anatomy|false|false|C1428865|fingersnull|Fingers, unit of measurement|LabModifier|false|false||fingersnull|GPSM2 gene|Finding|false|false|C0016129|pinsnull|Pins - Internal fixators|Device|false|false||pins
null|Pin Device Component|Device|false|false||pins
null|Medical pins|Device|false|false||pinsnull|Needle device|Device|false|false||needlesnull|Symptoms|Finding|false|false||symptomnull|null|Attribute|false|false||symptomnull|Dyspnea|Finding|false|false||SOBnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Minimal|Modifier|false|false||minimal
null|Mild (qualifier value)|Modifier|false|false||minimal
null|Minimum|Modifier|false|false||minimalnull|Increased sweating|Finding|false|false||diaphoresisnull|Gastroesophageal reflux disease|Disorder|false|false||gerdnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Tylenol|Drug|false|false||tylenol
null|Tylenol|Drug|false|false||tylenolnull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Hypertensive disease|Disorder|false|false||HTNnull|Asthma|Disorder|false|false||Asthmanull|Diverticulitis|Disorder|false|false||Diverticulitisnull|Several|LabModifier|false|false||severalnull|year|Time|false|false||yearsnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|Right hip region structure|Anatomy|false|false|C1292890;C1430701;C0529134;C1505163;C1654726;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1555302;C0035139;C0392806;C0559956|R hipnull|Prosthetic arthroplasty of hip (procedure)|Procedure|false|false|C0022122;C0228391;C0019552;C4299095;C0524470|hip replacementnull|heme iron polypeptide|Drug|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|hip
null|ST13 protein, human|Drug|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|hip
null|ST13 protein, human|Drug|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|hip
null|RPL29 protein, human|Drug|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|hip
null|RPL29 protein, human|Drug|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|hip
null|HHIP protein, human|Drug|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|hip
null|HHIP protein, human|Drug|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|hip
null|heme iron polypeptide|Drug|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|hipnull|RPL29 wt Allele|Finding|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|hip
null|REG3A gene|Finding|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|hip
null|RPL29 gene|Finding|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|hip
null|ST13 wt Allele|Finding|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|hip
null|ST13 gene|Finding|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|hip
null|HHIP gene|Finding|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|hip
null|HHIP wt Allele|Finding|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|hip
null|REG3A wt Allele|Finding|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|hipnull|Procedure on hip|Procedure|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|hipnull|Lower extremity>Hip|Anatomy|false|false|C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1430701;C0529134;C1505163;C1654726;C0392806;C1555302;C0035139;C0559956;C1292890|hip
null|Hip structure|Anatomy|false|false|C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1430701;C0529134;C1505163;C1654726;C0392806;C1555302;C0035139;C0559956;C1292890|hip
null|Structure of habenulopeduncular tract|Anatomy|false|false|C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1430701;C0529134;C1505163;C1654726;C0392806;C1555302;C0035139;C0559956;C1292890|hip
null|Bone structure of ischium|Anatomy|false|false|C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1430701;C0529134;C1505163;C1654726;C0392806;C1555302;C0035139;C0559956;C1292890|hipnull|Replacement|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C0524470|replacementnull|Replacement - supply|Procedure|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|replacement
null|Surgical Replantation|Procedure|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|replacementnull|Social and personal history|Finding|false|false||Social History
null|Social History|Finding|false|false||Social Historynull|Social|Finding|false|false||Socialnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Family Medical History|Finding|false|false||Family Historynull|Entity Name Part Type - family|Finding|false|false||Family
null|Last Name|Finding|false|false||Family
null|Living Arrangement - Family|Finding|false|false||Family
null|Family (taxonomic)|Finding|false|false||Family
null|Family Collection|Finding|false|false||Familynull|Family|Subject|false|false||Familynull|History of present illness (finding)|Finding|false|true||History
null|History of previous events|Finding|false|true||History
null|Historical aspects qualifier|Finding|false|true||History
null|Medical History|Finding|false|true||History
null|Concept History|Finding|false|true||Historynull|History|Subject|false|false||Historynull|Relationship - Mother|Finding|false|false||Mothernull|Mother (person)|Subject|false|false||Mothernull|Hypertensive disease|Disorder|false|false||HTNnull|Indirect exposure mechanism - Father|Finding|false|false||Father
null|Relationship - Father|Finding|false|false||Father
null|Father - courtesy title|Finding|false|false||Fathernull|Father (person)|Subject|false|false||Fathernull|Brother - courtesy title|Finding|false|false||Brother
null|Relationship - Brother|Finding|false|false||Brothernull|Brothers|Subject|false|false||Brothernull|Brother - courtesy title|Finding|false|false||Brother
null|Relationship - Brother|Finding|false|false||Brothernull|Brothers|Subject|false|false||Brothernull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Generalnull|General medical service|Procedure|false|false||Generalnull|Generalized|Modifier|false|false||Generalnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|false|false||acutenull|Emotional distress|Finding|true|false||distress
null|Distress|Finding|true|false||distressnull|HEENT|Anatomy|false|false||HEENTnull|Scleral Diseases|Disorder|false|false|C0036410;C0521367|Scleranull|examination of sclera|Procedure|false|false|C0036410;C0521367|Scleranull|Sclera|Anatomy|false|false|C2228481;C0026987;C0036412;C0205180|Scleranull|Anicteric|Finding|false|false|C0036410|anictericnull|Myelofibrosis|Disorder|false|false|C0694605;C0036410|MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false|C0026987|MMMnull|Oropharyngeal|Anatomy|false|false|C2228481;C1550016;C0036412|oropharynxnull|Remote control command - Clear|Finding|false|false|C0521367|clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|Neck
null|Neck problem|Finding|false|false|C0027530;C3159206|Necknull|dendritic spine neck|Anatomy|false|false|C0332254;C0812434;C0684335;C0428897|Neck
null|Neck|Anatomy|false|false|C0332254;C0812434;C0684335;C0428897|Necknull|Supple|Finding|false|false|C0027530;C3159206|supplenull|Jugular venous pressure|Finding|false|false|C0027530;C3159206|JVPnull|Elevated|Modifier|false|false||elevated
null|High|Modifier|false|false||elevatednull|Leukocyte adhesion deficiency type 1|Disorder|true|false|C0226032|LAD
null|Leukocyte adhesion deficiency|Disorder|true|false|C0226032|LADnull|ITGB2 wt Allele|Finding|true|false|C0226032|LAD
null|DLD gene|Finding|true|false|C0226032|LADnull|Anterior descending branch of left coronary artery|Anatomy|true|false|C1414063;C1706333;C5550999;C0398738|LADnull|Ladino Language|Entity|true|false||LADnull|Lung|Anatomy|false|false||Lungsnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Auscultation|Procedure|false|false||auscultationnull|Wheezing|Finding|true|false||wheezesnull|Basilar Rales|Finding|false|false||rales
null|Rales|Finding|false|false||ralesnull|Regular|Modifier|false|false||Regularnull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Rhythm|Finding|false|false||rhythm
null|rhythmic process (biological)|Finding|false|false||rhythmnull|Heart murmur|Finding|true|false||murmursnull|Pericardial friction rub|Finding|true|false||rubsnull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|Abdomennull|Abdomen problem|Finding|false|false|C0230168;C0000726|Abdomennull|Abdomen|Anatomy|false|false|C0153662;C0941288|Abdomen
null|Abdominal Cavity|Anatomy|false|false|C0153662;C0941288|Abdomennull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|Bowel sounds|Finding|false|false|C0021853|bowel soundsnull|Intestines|Anatomy|false|false|C0232693|bowelnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Rebound tenderness|Finding|true|false||rebound tendernessnull|Emotional tenderness|Finding|true|false||tenderness
null|Sore to touch|Finding|true|false||tendernessnull|Protective muscle spasm|Finding|true|false||guardingnull|Organomegaly|Finding|true|false||organomegalynull|Hereditary Multiple Exostoses|Disorder|false|false||Extnull|EXT1 wt Allele|Finding|false|false||Ext
null|EXT1 gene|Finding|false|false||Extnull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Clubbing|Disorder|true|false||clubbingnull|Cyanosis|Finding|true|false||cyanosisnull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0851353;C0005768;C0229664;C0005767|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0005768;C0229664;C0005767;C0851353|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C0014792;C1114281|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0005768;C0229664;C0005767;C0851353|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C0014792;C1114281|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MB
null|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MBnull|creatine kinase activity|Finding|false|false||CK-MBnull|Serum creatine phosphokinase MB isoenzyme measurement|Procedure|false|false||CK-MB
null|Creatine kinase MB measurement|Procedure|false|false||CK-MBnull|MB 3|Drug|false|false||MB-3null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MB
null|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MBnull|creatine kinase activity|Finding|false|false||CK-MBnull|Serum creatine phosphokinase MB isoenzyme measurement|Procedure|false|false||CK-MB
null|Creatine kinase MB measurement|Procedure|false|false||CK-MBnull|Cardiovascular system|Anatomy|false|false|C0809864;C1718621;C1705923;C0038435;C0684224;C0947630;C2603343;C0008972;C0700287;C0723460;C4255046|Cardiologynull|cardiology (field)|Title|false|false||Cardiologynull|Cardiology service|Entity|false|false||Cardiologynull|Report (document)|Finding|false|false|C0007226|Reportnull|Reporting|Procedure|false|false|C0007226|Reportnull|null|Attribute|false|false|C0007226|Reportnull|stress study|Procedure|false|false|C0007226|Stress Studynull|Stress bismuth subsalicylate|Drug|false|false|C0007226|Stress
null|Stress bismuth subsalicylate|Drug|false|false|C0007226|Stressnull|Stress|Finding|false|false|C0007226|Stressnull|W stress|Attribute|false|false|C0007226|Stressnull|Study Object|Finding|false|false|C0007226|Studynull|Scientific Study|Procedure|false|false|C0007226|Study
null|Study|Procedure|false|false|C0007226|Study
null|Clinical Research|Procedure|false|false|C0007226|Studynull|Room of building - Study|Device|false|false||Studynull|Exercise|Finding|false|false||EXERCISEnull|Exercise Pain Management|Procedure|false|false||EXERCISEnull|Rest|Finding|false|false||RESTINGnull|Data|Finding|false|false||DATAnull|Data call receiving device|Device|false|false||DATAnull|Data <Amphipyrinae>|Entity|false|false||DATAnull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false|C1305231;C0030471|SINUS
null|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false|C1305231;C0030471|SINUSnull|pathologic fistula|Disorder|false|false|C1305231;C0030471|SINUSnull|Sinus - general anatomical term|Anatomy|false|false|C5676667;C0016169;C0023211;C0723346|SINUS
null|Nasal sinus|Anatomy|false|false|C5676667;C0016169;C0023211;C0723346|SINUSnull|Anti-enterocyte antibody positivity|Finding|false|false|C1305231;C0030471|AEAnull|Left Bundle-Branch Block|Disorder|false|false|C1305231;C0030471|LBBBnull|null|Lab|false|false||LBBBnull|null|Finding|false|false|C4037974;C0018787|HEART RATEnull|examination of heart rate|Procedure|false|false|C4037974;C0018787|HEART RATEnull|heart rate|Attribute|false|false|C4037974;C0018787|HEART RATE
null|null|Attribute|false|false|C4037974;C0018787|HEART RATEnull|Mean Heart Rate|LabModifier|false|false||HEART RATEnull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|HEART
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|HEARTnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|HEARTnull|Chest>Heart|Anatomy|false|false|C2197023;C2041121;C0018810;C0488794;C0153957;C0153500;C0795691;C0871208;C1549480|HEART
null|Heart|Anatomy|false|false|C2197023;C2041121;C0018810;C0488794;C0153957;C0153500;C0795691;C0871208;C1549480|HEARTnull|Amount type - Rate|Finding|false|false|C4037974;C0018787|RATEnull|Rating (action)|Event|false|false|C4037974;C0018787|RATEnull|Rate|LabModifier|false|false||RATEnull|Blood pressure finding|Finding|false|false||BLOOD PRESSURE
null|Systemic arterial pressure|Finding|false|false||BLOOD PRESSURE
null|Blood Pressure|Finding|false|false||BLOOD PRESSUREnull|Blood pressure determination|Procedure|false|false||BLOOD PRESSUREnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Pressure (finding)|Finding|false|false||PRESSURE
null|null|Finding|false|false||PRESSURE
null|Baresthesia|Finding|false|false||PRESSUREnull|null|Phenomenon|false|false||PRESSUREnull|Pressure (property)|LabModifier|false|false||PRESSUREnull|Clinical trial protocol document|Finding|false|false||PROTOCOL
null|Study Protocol|Finding|false|false||PROTOCOL
null|Protocols documentation|Finding|false|false||PROTOCOL
null|Protocol - answer to question|Finding|false|false||PROTOCOL
null|Library Protocol|Finding|false|false||PROTOCOLnull|Tumor stage|Attribute|false|false||STAGEnull|Stage|Time|false|false||STAGE
null|Phase|Time|false|false||STAGEnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||TIME
null|Time (foundation metadata concept)|Finding|false|false||TIME
null|Value type - Time|Finding|false|false||TIME
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||TIME
null|Data types - Time|Finding|false|false||TIME
null|null|Finding|false|false||TIMEnull|Time|Time|false|false||TIMEnull|methamphetamine|Drug|false|false||SPEED
null|amphetamine|Drug|false|false||SPEED
null|amphetamine|Drug|false|false||SPEED
null|methamphetamine|Drug|false|false||SPEED
null|methamphetamine|Drug|false|false||SPEEDnull|Speed (motion)|LabModifier|false|false||SPEEDnull|Elevation procedure|Procedure|false|false|C4037974;C0018787|ELEVATIONnull|Elevation|Modifier|false|false||ELEVATIONnull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|HEART
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|HEARTnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|HEARTnull|Chest>Heart|Anatomy|false|false|C0153957;C0153500;C0795691;C0439775|HEART
null|Heart|Anatomy|false|false|C0153957;C0153500;C0795691;C0439775|HEARTnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Minangkabau Language|Entity|false|false||MINnull|Minute of time|Time|false|false||MINnull|Minimum|Modifier|false|false||MINnull|Minute Unit of Plane Angle|LabModifier|false|false||MIN
null|minim|LabModifier|false|false||MINnull|5,10-dihydro-5-methylphenazine|Drug|false|false||MPH
null|methylphenidate|Drug|false|false||MPH
null|methylphenidate|Drug|false|false||MPHnull|Master of Public Health|Finding|false|false||MPHnull|Miles per hour|LabModifier|false|false||MPHnull|Amount type - Rate|Finding|false|false||RATEnull|Rating (action)|Event|false|false||RATEnull|Rate|LabModifier|false|false||RATEnull|Pressure (finding)|Finding|false|false||PRESSURE
null|null|Finding|false|false||PRESSURE
null|Baresthesia|Finding|false|false||PRESSUREnull|null|Phenomenon|false|false||PRESSUREnull|Pressure (property)|LabModifier|false|false||PRESSUREnull|Total exercise time|Time|false|false||TOTAL EXERCISE TIMEnull|Total|Modifier|false|false||TOTALnull|Exercise time|Time|false|false||EXERCISE TIMEnull|Exercise|Finding|false|false||EXERCISEnull|Exercise Pain Management|Procedure|false|false||EXERCISEnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||TIME
null|Time (foundation metadata concept)|Finding|false|false||TIME
null|Value type - Time|Finding|false|false||TIME
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||TIME
null|Data types - Time|Finding|false|false||TIME
null|null|Finding|false|false||TIMEnull|Time|Time|false|false||TIMEnull|MAX protein, human|Drug|false|false||MAX
null|MAX protein, human|Drug|false|false||MAXnull|Max (cigarettes)|Finding|false|false||MAX
null|Oncogene MAX|Finding|false|false||MAX
null|MAX gene|Finding|false|false||MAXnull|Maximum|LabModifier|false|false||MAXnull|Hormone replacement therapy|Procedure|false|false||HRTnull|null|Attribute|false|false||HRT
null|null|Attribute|false|false||HRTnull|Amount type - Rate|Finding|false|false||RATEnull|Rating (action)|Event|false|false||RATEnull|Rate|LabModifier|false|false||RATEnull|Achieved|Finding|false|false||ACHIEVEDnull|Symptoms aspect|Finding|false|false||SYMPTOMS
null|Symptoms|Finding|false|false||SYMPTOMSnull|atypia morphology|Finding|false|false||ATYPICALnull|Atypical|Modifier|false|false||ATYPICALnull|Peak level|Modifier|false|false||PEAKnull|With intensity|Modifier|false|false||INTENSITYnull|Interpretation Process|Finding|false|false||INTERPRETATIONnull|null|Attribute|false|false||INTERPRETATIONnull|Woman|Subject|false|false||woman
null|Human, Female adult|Subject|false|false||womannull|atypia morphology|Finding|false|false||atypicalnull|Atypical|Modifier|false|false||atypicalnull|Chest discomfort|Finding|false|false|C1527391;C0817096|chest discomfortnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C2364135;C0741025;C0235710|chest
null|Anterior thoracic region|Anatomy|false|false|C2364135;C0741025;C0235710|chestnull|Discomfort|Finding|false|false|C1527391;C0817096|discomfortnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Minute of time|Time|false|false||minutesnull|Minute Unit of Plane Angle|LabModifier|false|false||minutes
null|Minute (diminutive)|LabModifier|false|false||minutes
null|Small|LabModifier|false|false||minutesnull|Clinical trial protocol document|Finding|false|false||protocol
null|Study Protocol|Finding|false|false||protocol
null|Protocols documentation|Finding|false|false||protocol
null|Protocol - answer to question|Finding|false|false||protocol
null|Library Protocol|Finding|false|false||protocolnull|Fair - language proficiency|Modifier|false|false||fair
null|Fair (qualifier value)|Modifier|false|false||fair
null|Fair Specimen Quality|Modifier|false|false||fairnull|null|Finding|false|false||exercise tolerancenull|null|Attribute|false|false||exercise tolerance
null|Exercise Tolerance|Attribute|false|false||exercise tolerancenull|Exercise|Finding|false|false||exercisenull|Exercise Pain Management|Procedure|false|false||exercisenull|Physiologic tolerance|Finding|false|false||tolerance
null|Mental tolerance|Finding|false|false||tolerance
null|Immune Tolerance|Finding|false|false||tolerance
null|Drug Tolerance|Finding|false|false||tolerancenull|Tolerance|Modifier|false|false||tolerancenull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|ETV3 wt Allele|Finding|false|false||METS
null|ETV3 gene|Finding|false|false||METSnull|Exercise stress test|Procedure|false|false|C4318744|exercise testnull|Exercise|Finding|false|false|C4318744|exercisenull|Exercise Pain Management|Procedure|false|false|C4318744|exercisenull|Tests (qualifier value)|Finding|false|false|C4318744|test
null|Testing|Finding|false|false|C4318744|testnull|Laboratory Procedures|Procedure|false|false|C4318744|testnull|Test - temporal region|Anatomy|false|false|C0015259;C0015260;C0039593;C0392366;C0022885;C0456984;C1522704;C1578483;C1550655;C1578481;C1578486;C1578484;C1578485;C1553888;C1522634;C1553397|testnull|Test Result|Lab|false|false|C4318744|testnull|Test Dosing Unit|LabModifier|false|false||testnull|Relationship modifier - Patient|Finding|false|false|C4318744|patient
null|Specimen Type - Patient|Finding|false|false|C4318744|patient
null|Mail Claim Party - Patient|Finding|false|false|C4318744|patient
null|Report source - Patient|Finding|false|false|C4318744|patient
null|null|Finding|false|false|C4318744|patient
null|Disabled Person Code - Patient|Finding|false|false|C4318744|patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Request - ActReason|Finding|false|false|C4318744|request
null|request - ActMood|Finding|false|false|C4318744|request
null|Question (inquiry)|Finding|false|false|C4318744|requestnull|null|Event|false|false||requestnull|Secondary to|Modifier|false|false||secondary tonull|Neoplasm Metastasis|Disorder|false|false||secondarynull|metastatic qualifier|Finding|false|false||secondarynull|Secondary to|Modifier|false|false||secondarynull|second (number)|LabModifier|false|false||secondarynull|Fatigue|Finding|false|false||fatiguenull|During exercise|Time|false|false||During exercisenull|Exercise|Finding|false|false||exercisenull|Exercise Pain Management|Procedure|false|false||exercisenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Bed Status - Isolated|Finding|false|false||isolated
null|Isolated|Finding|false|false||isolatednull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Left sided|Modifier|false|false||left-sidednull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Chest discomfort|Finding|false|false|C1527391;C0817096|chest discomfortnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C2364135;C0741025;C0235710|chest
null|Anterior thoracic region|Anatomy|false|false|C2364135;C0741025;C0235710|chestnull|Discomfort|Finding|false|false|C1527391;C0817096|discomfortnull|Academic Research Enhancement Awards|Event|false|false||areanull|Geographic Locations|Entity|false|false||areanull|Area|Modifier|false|false||areanull|Discomfort|Finding|false|false||discomfortnull|Tender|Modifier|false|false||tendernull|Palpation|Procedure|false|false||palpationnull|Discomfort|Finding|false|false||discomfortnull|REST protein, human|Drug|false|false||rest
null|REST protein, human|Drug|false|false||restnull|REST gene|Finding|false|false||rest
null|site-specific telomere resolvase activity|Finding|false|false||rest
null|Rest|Finding|false|false||restnull|Absent|Finding|false|false||absentnull|Expression Negative|Lab|false|false||absentnull|Minute of time|Time|false|false||minutesnull|Minute Unit of Plane Angle|LabModifier|false|false||minutes
null|Minute (diminutive)|LabModifier|false|false||minutes
null|Small|LabModifier|false|false||minutesnull|Present|Finding|false|false||presence ofnull|Providing presence (regime/therapy)|Procedure|false|false||presencenull|Presence (property)|Modifier|false|false||presencenull|Left Bundle-Branch Block|Disorder|false|false||LBBBnull|null|Lab|false|false||LBBBnull|Uninterpretable|Modifier|false|false||uninterpretablenull|Ischemia|Finding|false|false||ischemianull|Ischemia Procedure|Procedure|false|false||ischemianull|Rhythm|Finding|false|false||rhythm
null|rhythmic process (biological)|Finding|false|false||rhythmnull|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false|C1305231;C0030471|sinus
null|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false|C1305231;C0030471|sinusnull|pathologic fistula|Disorder|false|false|C1305231;C0030471|sinusnull|Sinus - general anatomical term|Anatomy|false|false|C0016169;C0723346|sinus
null|Nasal sinus|Anatomy|false|false|C0016169;C0723346|sinusnull|Frequently|Time|false|false||frequentnull|Bed Status - Isolated|Finding|false|false||isolated
null|Isolated|Finding|false|false||isolatednull|pamidronate|Drug|false|false||APDs
null|pamidronate|Drug|false|false||APDsnull|ACTIVATED PI3K-DELTA SYNDROME|Disorder|false|false||APDsnull|PIK3CD wt Allele|Finding|false|false||APDsnull|Infrequent|Time|false|false||occasionalnull|Heart Atrium|Anatomy|false|false|C0429001|atrialnull|Paired ventricular premature complexes|Finding|false|false|C0018792;C0018792|coupletsnull|Heart Atrium|Anatomy|false|false|C0429001|atrialnull|Triplet Multiple Birth|Subject|false|false||tripletsnull|Rest|Finding|false|false||Restingnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Systolic Hypertension|Disorder|false|false||systolic hypertensionnull|Systole|Finding|false|false||systolicnull|Hypertensive disease|Disorder|false|false||hypertensionnull|Blood pressure finding|Finding|false|false||blood pressure
null|Systemic arterial pressure|Finding|false|false||blood pressure
null|Blood Pressure|Finding|false|false||blood pressurenull|Blood pressure determination|Procedure|false|false||blood pressurenull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Communication Response|Finding|false|false||response
null|Disease Response|Finding|false|false||response
null|Answer (statement)|Finding|false|false||responsenull|Response process|Subject|false|false||responsenull|Exercise|Finding|false|false||exercisenull|Exercise Pain Management|Procedure|false|false||exercisenull|Heart rate response (observable entity)|Attribute|false|false|C4037974;C0018787|heart rate responsenull|null|Finding|false|false|C4037974;C0018787|heart ratenull|examination of heart rate|Procedure|false|false|C4037974;C0018787|heart ratenull|heart rate|Attribute|false|false|C4037974;C0018787|heart rate
null|null|Attribute|false|false|C4037974;C0018787|heart ratenull|Mean Heart Rate|LabModifier|false|false||heart ratenull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C2197023;C0795691;C2911692;C1706817;C1704632;C1549480;C0153957;C0153500;C0018810;C0488794;C1997754;C2041121;C0871208|heart
null|Heart|Anatomy|false|false|C2197023;C0795691;C2911692;C1706817;C1704632;C1549480;C0153957;C0153500;C0018810;C0488794;C1997754;C2041121;C0871208|heartnull|Response Frequency|Time|false|false||rate responsenull|Amount type - Rate|Finding|false|false|C4037974;C0018787|ratenull|Rating (action)|Event|false|false|C4037974;C0018787|ratenull|Rate|LabModifier|false|false||ratenull|response to exercise|Finding|false|false||response to exercisenull|Communication Response|Finding|false|false|C4037974;C0018787|response
null|Disease Response|Finding|false|false|C4037974;C0018787|response
null|Answer (statement)|Finding|false|false|C4037974;C0018787|responsenull|Response process|Subject|false|false||responsenull|Exercise|Finding|false|false||exercisenull|Exercise Pain Management|Procedure|false|false||exercisenull|MILDLY|Modifier|false|false||mildly
null|Mild (qualifier value)|Modifier|false|false||mildlynull|Blunted|Modifier|false|false||bluntednull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Fair - language proficiency|Modifier|false|false||Fair
null|Fair (qualifier value)|Modifier|false|false||Fair
null|Fair Specimen Quality|Modifier|false|false||Fairnull|null|Finding|false|false||exercise tolerancenull|null|Attribute|false|false||exercise tolerance
null|Exercise Tolerance|Attribute|false|false||exercise tolerancenull|Exercise|Finding|false|false||exercisenull|Exercise Pain Management|Procedure|false|false||exercisenull|Physiologic tolerance|Finding|false|false||tolerance
null|Mental tolerance|Finding|false|false||tolerance
null|Immune Tolerance|Finding|false|false||tolerance
null|Drug Tolerance|Finding|false|false||tolerancenull|Tolerance|Modifier|false|false||tolerancenull|Symptoms aspect|Finding|true|false||symptoms
null|Symptoms|Finding|true|false||symptomsnull|Uninterpretable|Modifier|false|false||uninterpretablenull|Equine Gonadotropins|Drug|false|false||ECG
null|Equine Gonadotropins|Drug|false|false||ECG
null|Equine Gonadotropins|Drug|false|false||ECGnull|Electrocardiogram image|Finding|false|false||ECG
null|Electrocardiogram|Finding|false|false||ECGnull|Electrocardiography|Procedure|false|false||ECGnull|Workload|LabModifier|false|false||workloadnull|Rest|Finding|false|false||Restingnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Systole|Finding|false|false||systolicnull|Hypertensive disease|Disorder|false|false||hypertensionnull|Appropriate|Modifier|false|false||appropriatenull|Speed of blood pressure response|Attribute|false|false||blood pressure responsenull|Blood pressure finding|Finding|false|false||blood pressure
null|Systemic arterial pressure|Finding|false|false||blood pressure
null|Blood Pressure|Finding|false|false||blood pressurenull|Blood pressure determination|Procedure|false|false||blood pressurenull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Communication Response|Finding|false|false||response
null|Disease Response|Finding|false|false||response
null|Answer (statement)|Finding|false|false||responsenull|Response process|Subject|false|false||responsenull|Exercise|Finding|false|false||exercisenull|Exercise Pain Management|Procedure|false|false||exercisenull|Suboptimal|Modifier|false|false||Suboptimalnull|Study Object|Finding|false|false||studynull|Scientific Study|Procedure|false|false||study
null|Study|Procedure|false|false||study
null|Clinical Research|Procedure|false|false||studynull|Room of building - Study|Device|false|false||studynull|Target heart rate|Procedure|false|false|C4037974;C0018787|target heart ratenull|Target|Finding|false|false||targetnull|Therapeutically Applicable Research to Generate Effective Treatments|Procedure|false|false|C4037974;C0018787|targetnull|null|Finding|false|false|C4037974;C0018787|heart ratenull|examination of heart rate|Procedure|false|false|C4037974;C0018787|heart ratenull|heart rate|Attribute|false|false|C4037974;C0018787|heart rate
null|null|Attribute|false|false|C4037974;C0018787|heart ratenull|Mean Heart Rate|LabModifier|false|false||heart ratenull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C1549480;C5575831;C0744682;C0795691;C0153957;C0153500;C0018810;C0488794;C0871208;C2197023;C2041121|heart
null|Heart|Anatomy|false|false|C1549480;C5575831;C0744682;C0795691;C0153957;C0153500;C0018810;C0488794;C0871208;C2197023;C2041121|heartnull|Amount type - Rate|Finding|false|false|C4037974;C0018787|ratenull|Rating (action)|Event|false|false|C4037974;C0018787|ratenull|Rate|LabModifier|false|false||ratenull|BRIEF Health Literacy Screening Tool|Finding|false|false||Brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||Briefnull|Brief|Time|false|false||Briefnull|Shortened|Modifier|false|false||Briefnull|Hospital course|Finding|false|false||Hospital Coursenull|null|Attribute|false|false||Hospital Coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||Coursenull|Several|LabModifier|false|false||severalnull|Transaction counts and value totals - month|Finding|false|false||month
null|Precision - month|Finding|false|false||monthnull|month|Time|false|false||month
null|Monthly (qualifier value)|Time|false|false||monthnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Left sided|Modifier|false|false||left sided
null|Left|Modifier|false|false||left sidednull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Anorectal Malformations|Disorder|false|false|C0446516;C1140618;C1269078|armnull|AKR1A1 wt Allele|Finding|false|false|C0446516;C1140618;C1269078|arm
null|ARMC9 gene|Finding|false|false|C0446516;C1140618;C1269078|armnull|Protocol Treatment Arm|Procedure|false|false|C0446516;C1140618;C1269078|arm
null|Axillary Reverse Mapping|Procedure|false|false|C0446516;C1140618;C1269078|arm
null|Study Arm|Procedure|false|false|C0446516;C1140618;C1269078|armnull|Upper arm|Anatomy|false|false|C1824218;C3715044;C3495676;C1522541;C5400986;C4761640|arm
null|null|Anatomy|false|false|C1824218;C3715044;C3495676;C1522541;C5400986;C4761640|arm
null|Upper Extremity|Anatomy|false|false|C1824218;C3715044;C3495676;C1522541;C5400986;C4761640|armnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0741025|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025|chestnull|Walls of a building|Device|false|false||wallnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Left Bundle-Branch Block|Disorder|false|false||LBBBnull|null|Lab|false|false||LBBBnull|Chest Pain|Finding|false|false|C1527391;C0817096|Chest Painnull|null|Attribute|false|false|C1527391;C0817096|Chest Painnull|Chest problem|Finding|false|false|C1527391;C0817096|Chestnull|Chest|Anatomy|false|false|C1549543;C0030193;C0008031;C2926613;C0741025|Chest
null|Anterior thoracic region|Anatomy|false|false|C1549543;C0030193;C0008031;C2926613;C0741025|Chestnull|Administration Method - Pain|Finding|false|false|C1527391;C0817096|Pain
null|Pain|Finding|false|false|C1527391;C0817096|Painnull|null|Attribute|false|false||Painnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Nature|Finding|false|false|C0262187|nature
null|Natures|Finding|false|false|C0262187|naturenull|ACSS2 protein, human|Drug|false|false|C0262187|ACS
null|ACSS2 protein, human|Drug|false|false|C0262187|ACSnull|Acrocallosal Syndrome|Disorder|false|false|C0262187|ACS
null|Acute Chest Syndrome|Disorder|false|false|C0262187|ACSnull|ACS - Activity Card Sort|Finding|false|false|C0262187|ACS
null|American Community Survey|Finding|false|false|C0262187|ACS
null|ACCS gene|Finding|false|false|C0262187|ACS
null|CO-methylating acetyl-CoA synthase activity|Finding|false|false|C0262187|ACS
null|PLA2G15 gene|Finding|false|false|C0262187|ACS
null|ACSS2 wt Allele|Finding|false|false|C0262187|ACS
null|ACSS2 gene|Finding|false|false|C0262187|ACS
null|acetate-CoA ligase activity|Finding|false|false|C0262187|ACSnull|anterior calcarine sulcus (human only)|Anatomy|false|false|C1825842;C5400867;C4318612;C1842089;C1424787;C1150760;C2266615;C5551036;C1262865;C0349590;C0742343;C0796147;C4042561|ACSnull|Alternate Care Site|Device|false|false||ACSnull|American College of Surgeons|Entity|false|false||ACS
null|American Cancer Society|Entity|false|false||ACS
null|Alternate Care Site|Entity|false|false||ACSnull|Several|LabModifier|false|false||severalnull|Cardiac attachment|Finding|false|false|C0018787|cardiacnull|Heart|Anatomy|false|false|C1314974|cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||cardiacnull|risk factors - observation list|Finding|false|false||risk factors
null|risk factors|Finding|false|false||risk factors
null|History of - risk factor|Finding|false|false||risk factorsnull|null|Attribute|false|false||risk factorsnull|Risk|Finding|false|false||risknull|Left Bundle-Branch Block|Disorder|false|false||LBBBnull|null|Lab|false|false||LBBBnull|Physicians|Subject|false|false||physiciansnull|HTRA2 gene|Finding|false|false||oMInull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|Living Alone|Finding|false|false||alonenull|alone - group size|Subject|false|false||alonenull|Singular|LabModifier|false|false||alonenull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Echocardiography, Stress|Procedure|false|false||Stress Echonull|Stress bismuth subsalicylate|Drug|false|false||Stress
null|Stress bismuth subsalicylate|Drug|false|false||Stressnull|Stress|Finding|false|false||Stressnull|W stress|Attribute|false|false||Stressnull|ECHO protocol|Procedure|false|false||Echo
null|Extension for Community Healthcare Outcomes|Procedure|false|false||Echonull|Echo <Calopterygidae>|Entity|false|false||Echonull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|regional|Modifier|false|false||regional
null|Local|Modifier|false|false||regionalnull|DYSFUNCTION - SKIN DISORDERS|Disorder|false|false||dysfunctionnull|Dysfunction|Finding|false|false||dysfunction
null|physiopathological|Finding|false|false||dysfunction
null|Functional disorder|Finding|false|false||dysfunctionnull|Hypokinesia|Finding|false|false||hypokinesisnull|inferiority|Finding|false|false||inferiornull|Inferior|Modifier|false|false||inferiornull|Inferolateral|Modifier|false|false||inferolateralnull|Walls of a building|Device|false|false||wallsnull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|Single vessel disease|Disorder|false|false||single vessel diseasenull|Marital Status - Single|Finding|false|false||single
null|Unmarried|Finding|false|false||singlenull|Singular|LabModifier|false|false||singlenull|Vessel Positions|Anatomy|false|false||vessel
null|Blood Vessel|Anatomy|false|false||vesselnull|Vessel (unit of presentation)|LabModifier|false|false||vesselnull|Disease|Disorder|false|false||diseasenull|Pancreatic Ductal Adenocarcinoma|Disorder|false|false|C0226047|PDA
null|PATENT DUCTUS ARTERIOSUS 1|Disorder|false|false|C0226047|PDA
null|Patent ductus arteriosus|Disorder|false|false|C0226047|PDAnull|Posterior interventricular branch of right coronary artery|Anatomy|false|false|C1335302;C0013274;C4282128;C5779816;C1704711|PDAnull|Distribution [PK]|Finding|false|false|C0226047|distribution
null|Distribution|Finding|false|false|C0226047|distributionnull|Spatial Distribution|Modifier|false|false||distributionnull|Cardiovascular system|Anatomy|false|false|C0009818|cardiologynull|cardiology (field)|Title|false|false||cardiologynull|Cardiology service|Entity|false|false||cardiologynull|Consultation|Procedure|false|false|C0007226|consultnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|aspirin|Drug|false|false||aspirin
null|aspirin|Drug|false|false||aspirinnull|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Drug|false|false||statin
null|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Drug|false|false||statinnull|EEF1A2 gene|Finding|false|false||statinnull|3-hydroxy-3-methylglutaryl-coenzyme A reductase inhibitor (disposition)|Modifier|false|false||statinnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Asthma|Disorder|false|false||asthmanull|Release - action (qualifier value)|Finding|false|false|C0007226|release
null|Released (action)|Finding|false|false|C0007226|releasenull|Discharge (release)|Procedure|false|false|C0007226|release
null|Release (procedure)|Procedure|false|false|C0007226|release
null|Patient Discharge|Procedure|false|false|C0007226|releasenull|diltiazem|Drug|false|false||diltiazem
null|diltiazem|Drug|false|false||diltiazemnull|Instructions|Finding|false|false|C0007226|instructions
null|Instruction [Publication Type]|Finding|false|false|C0007226|instructionsnull|null|Attribute|false|false|C0007226|instructionsnull|Cardiovascular system|Anatomy|false|false|C1283071;C0391871;C3263700;C0030685;C0680255;C1963578;C1442085;C0302828|cardiologynull|cardiology (field)|Title|false|false||cardiologynull|Cardiology service|Entity|false|false||cardiologynull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Supraventricular tachycardia|Disorder|false|false||Supraventricular tachycardianull|Supraventricular Tachycardia by ECG Finding|Finding|false|false||Supraventricular tachycardianull|Tachycardia by ECG Finding|Finding|false|false||tachycardia
null|Tachycardia|Finding|false|false||tachycardianull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Numerous|LabModifier|false|false||multiplenull|Does run (finding)|Finding|false|false||runsnull|Supraventricular tachycardia|Disorder|false|false||SVTnull|Supraventricular Tachycardia by ECG Finding|Finding|false|false||SVTnull|Multinational Association of Supportive Care in Cancer Antiemesis Tool|Finding|false|false||MAT
null|MAT1A wt Allele|Finding|false|false||MAT
null|[acyl-carrier-protein] S-malonyltransferase activity|Finding|false|false||MAT
null|Multifocal atrial tachycardia|Finding|false|false||MAT
null|ACAT1 wt Allele|Finding|false|false||MAT
null|ACAT1 gene|Finding|false|false||MAT
null|MAT1A gene|Finding|false|false||MATnull|Mats|Device|false|false||MATnull|MAT Format|Modifier|false|false||MATnull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Obstructed|Finding|false|false||obstructivenull|Lung diseases|Disorder|false|false|C4037972;C0024109|lung diseasenull|Lung diseases|Disorder|false|false|C4037972;C0024109|lungnull|Lung Problem|Finding|false|false|C4037972;C0024109|lungnull|Chest>Lung|Anatomy|false|false|C0012634;C0024115;C0740941;C1947944;C0042153;C0457083;C0241361;C1547296;C0039773;C1555457;C0024115|lung
null|Lung|Anatomy|false|false|C0012634;C0024115;C0740941;C1947944;C0042153;C0457083;C0241361;C1547296;C0039773;C1555457;C0024115|lungnull|Disease|Disorder|false|false|C4037972;C0024109|diseasenull|Chronic - Admission Level of Care Code|Finding|false|false|C4037972;C0024109|chronicnull|Provision of recurring care for chronic illness|Procedure|false|false|C4037972;C0024109|chronicnull|chronic|Time|false|false||chronicnull|theophylline use|Finding|false|false|C4037972;C0024109|theophylline usenull|theophylline|Drug|false|false||theophylline
null|theophylline|Drug|false|false||theophyllinenull|Assay of theophylline|Procedure|false|false|C4037972;C0024109|theophyllinenull|Use - dosing instruction imperative|Finding|false|false|C4037972;C0024109|use
null|utilization qualifier|Finding|false|false|C4037972;C0024109|use
null|Usage|Finding|false|false|C4037972;C0024109|usenull|Cardiovascular system|Anatomy|false|false||Cardiologynull|cardiology (field)|Title|false|false||Cardiologynull|Cardiology service|Entity|false|false||Cardiologynull|theophylline|Drug|false|false||theophylline
null|theophylline|Drug|false|false||theophyllinenull|Assay of theophylline|Procedure|false|false||theophyllinenull|Pulmonologists|Subject|false|false||pulmonologistnull|Vitelliform Macular Dystrophy|Disorder|false|false||bestnull|BEST1 wt Allele|Finding|false|false||best
null|BEST1 gene|Finding|false|false||bestnull|best (quality)|Modifier|false|false||bestnull|Course|Time|false|false||coursenull|Clinical action|Finding|false|false||action
null|null|Finding|false|false||actionnull|Action|Event|false|false||actionnull|Instructions|Finding|false|false||instructions
null|Instruction [Publication Type]|Finding|false|false||instructionsnull|null|Attribute|false|false||instructionsnull|Use of|Finding|false|false||use ofnull|Use - dosing instruction imperative|Finding|false|false||use
null|utilization qualifier|Finding|false|false||use
null|Usage|Finding|false|false||usenull|theophylline|Drug|false|false||theophylline
null|theophylline|Drug|false|false||theophyllinenull|Assay of theophylline|Procedure|false|false||theophyllinenull|Pulmonologists|Subject|false|false||pulmonologistnull|Cardiovascular system|Anatomy|false|false||cardiologynull|cardiology (field)|Title|false|false||cardiologynull|Cardiology service|Entity|false|false||cardiologynull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|Tylenol|Drug|false|false||Tylenol
null|Tylenol|Drug|false|false||Tylenolnull|Every four hours|Time|false|false||Q4hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|albuterol sulfate|Drug|false|false||Albuterol Sulfate
null|albuterol sulfate|Drug|false|false||Albuterol Sulfatenull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||Sulfate
null|Sulfates, Inorganic|Drug|false|false||Sulfate
null|sulfate ion|Drug|false|false||Sulfate
null|sulfate ion|Drug|false|false||Sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||Sulfatenull|Puff Dosing Unit|LabModifier|false|false||puffsnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Dyspnea|Finding|false|false||SOBnull|fluticasone|Drug|false|false||Fluticasone
null|fluticasone|Drug|false|false||Fluticasonenull|microgram|LabModifier|false|false||mcgnull|Spray Dosage Form|Drug|false|false||spraynull|Spray (administration method)|Finding|false|false||spraynull|Spray (action)|Event|false|false||spraynull|Spray Dosing Unit|LabModifier|false|false||spraynull|Suspension substance|Drug|false|false||suspension
null|Suspensions|Drug|false|false||suspensionnull|Suspension (action)|Finding|false|false||suspensionnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Hypersensitivity|Finding|false|false||allergiesnull|null|Attribute|false|false||allergiesnull|Inhalant dose form|Drug|false|false||INH
null|isoniazid|Drug|false|false||INH
null|isoniazid|Drug|false|false||INHnull|Inhalation Route of Administration|Finding|false|false||INHnull|Ingush language|Entity|false|false||INHnull|Inhalation Dosing Unit|LabModifier|false|false||INHnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|hydrochlorothiazide|Drug|false|false||HCTZ
null|hydrochlorothiazide|Drug|false|false||HCTZnull|Daily|Time|false|false||dailynull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|omeprazole|Drug|false|false||omeprazole
null|omeprazole|Drug|false|false||omeprazolenull|simvastatin|Drug|false|false||simvastatin
null|simvastatin|Drug|false|false||simvastatinnull|theophylline|Drug|false|false||theophylline
null|theophylline|Drug|false|false||theophyllinenull|Assay of theophylline|Procedure|false|false||theophyllinenull|Sustained Release Dosage Form|Drug|false|false||sustained releasenull|Sustained|Finding|false|false||sustainednull|Release - action (qualifier value)|Finding|false|false||release
null|Released (action)|Finding|false|false||releasenull|Discharge (release)|Procedure|false|false||release
null|Release (procedure)|Procedure|false|false||release
null|Patient Discharge|Procedure|false|false||releasenull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|Spiriva|Drug|false|false||spiriva
null|Spiriva|Drug|false|false||spirivanull|microgram|LabModifier|false|false||mcgnull|Inhalation Route of Administration|Finding|false|false||inhalation
null|Inspiration (function)|Finding|false|false||inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||inhalationnull|Arylsulfatase A, human|Drug|false|false||ASA
null|Arylsulfatase A, human|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASAnull|ARSA gene|Finding|false|false||ASAnull|CALCIUM SUPPLEMENTS|Drug|false|false|C0262329|Calcium
null|calcium|Drug|false|false|C0262329|Calcium
null|calcium|Drug|false|false|C0262329|Calcium
null|calcium|Drug|false|false|C0262329|Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false|C0262329|Calcium
null|Calcium, Dietary|Drug|false|false|C0262329|Calcium
null|Calcium [EPC]|Drug|false|false|C0262329|Calcium
null|Calcium Drug Class|Drug|false|false|C0262329|Calciumnull|Calcium metabolic function|Finding|false|false|C0262329|Calciumnull|Calcium measurement|Procedure|false|false|C0262329|Calciumnull|Receptors, Antigen, B-Cell|Drug|false|false|C0262329|sig
null|Receptors, Antigen, B-Cell|Drug|false|false|C0262329|signull|Receptors, Antigen, B-Cell|Finding|false|false|C0262329|signull|Short insular gyrus|Anatomy|false|false|C0201925;C0006726;C3540037;C0006675;C2936886;C3714611;C0034789;C1549115;C1547294;C1556129;C1546841;C1547312;C1548543;C1556120;C1556126;C3244284;C1556125;C1561529;C1556128;C1556127;C1556122;C1556121;C1556124;C1556123;C1548550;C1549105;C1609613;C1547283;C1547306;C1549064;C1556131;C1556130;C1546837;C1556137;C1556136;C1556133;C1556132;C1556135;C1556134;C0034789;C4553026|signull|Surveillance Implementation Group|Entity|false|false||sig
null|Staphylococcus intermedius group|Entity|false|false||signull|unknown vaccine or immune globulin|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|unknown vaccine or immune globulin|Drug|false|false||unknownnull|Unknown - Patient_s Relationship to Insured|Finding|false|false|C0262329|unknown
null|Unknown - Special Program Code|Finding|false|false|C0262329|unknown
null|Unknown - Production Class Code|Finding|false|false|C0262329|unknown
null|Unknown - Patient Outcome|Finding|false|false|C0262329|unknown
null|Unknown - Recreational Drug Use Code|Finding|false|false|C0262329|unknown
null|Unknown - Escort Required|Finding|false|false|C0262329|unknown
null|Unknown - Transport Arranged|Finding|false|false|C0262329|unknown
null|Unknown - Living Arrangement|Finding|false|false|C0262329|unknown
null|Unknown - Employment Status|Finding|false|false|C0262329|unknown
null|Unknown - Relationship|Finding|false|false|C0262329|unknown
null|Unknown - publishing section|Finding|false|false|C0262329|unknown
null|Unknown Publicity Code|Finding|false|false|C0262329|unknown
null|Unknown - Event reason|Finding|false|false|C0262329|unknown
null|Unknown - Religion|Finding|false|false|C0262329|unknown
null|Unknown - Organ Donor Code|Finding|false|false|C0262329|unknown
null|unknown - NullFlavor|Finding|false|false|C0262329|unknown
null|Unknown - Notify Clergy Code|Finding|false|false|C0262329|unknown
null|Unknown - Administrative Gender|Finding|false|false|C0262329|unknown
null|Unknown - Patient Condition Code|Finding|false|false|C0262329|unknown
null|Unknown - Living Will Code|Finding|false|false|C0262329|unknown
null|Marital Status - Unknown|Finding|false|false|C0262329|unknown
null|Unknown - mode of arrival code|Finding|false|false|C0262329|unknown
null|Unknown - Patient Class|Finding|false|false|C0262329|unknown
null|Unknown - Event Expected|Finding|false|false|C0262329|unknown
null|Unknown - Expanded yes/no indicator|Finding|false|false|C0262329|unknown
null|Unknown - Immunization Registry Status|Finding|false|false|C0262329|unknown
null|Unknown - Container status|Finding|false|false|C0262329|unknown
null|Unknown - CWE statuses|Finding|false|false|C0262329|unknown
null|Unknown - Job Status|Finding|false|false|C0262329|unknown
null|Unknown - Precaution Code|Finding|false|false|C0262329|unknown
null|Unknown - Contact Role|Finding|false|false|C0262329|unknown
null|Unknown - Living Dependency|Finding|false|false|C0262329|unknownnull|Ethnic group unknown|Subject|false|false||unknownnull|Unknown - Allergy Severity|Modifier|false|false||unknown
null|Unknown - HL7 update mode|Modifier|false|false||unknown
null|Unknown|Modifier|false|false||unknownnull|cod liver oil|Drug|false|false|C4037986;C1278929;C0023884|Cod liver oil
null|cod liver oil|Drug|false|false|C4037986;C1278929;C0023884|Cod liver oil
null|cod liver oil|Drug|false|false|C4037986;C1278929;C0023884|Cod liver oilnull|cod, unspecified preparation|Drug|false|false|C4037986;C1278929;C0023884|Cod
null|null|Drug|false|false|C4037986;C1278929;C0023884|Cod
null|Cyclophosphamide/Dacarbazine/Vincristine|Drug|false|false|C4037986;C1278929;C0023884|Cod
null|cod, unspecified preparation|Drug|false|false|C4037986;C1278929;C0023884|Cod
null|codfish allergenic extract|Drug|false|false|C4037986;C1278929;C0023884|Cod
null|codfish allergenic extract|Drug|false|false|C4037986;C1278929;C0023884|Codnull|Cancerization of Pancreatic Ducts|Finding|false|false|C4037986;C1278929;C0023884|Cod
null|Cemento-osseous dysplasia|Finding|false|false|C4037986;C1278929;C0023884|Cod
null|SNRPB gene|Finding|false|false|C4037986;C1278929;C0023884|Cod
null|Cause of Death|Finding|false|false|C4037986;C1278929;C0023884|Codnull|Cod|Entity|false|false||Codnull|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|false|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|false|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|livernull|Benign neoplasm of liver|Disorder|false|false|C4037986;C1278929;C0023884|liver
null|Liver diseases|Disorder|false|false|C4037986;C1278929;C0023884|livernull|Liver problem|Finding|false|false|C4037986;C1278929;C0023884|livernull|Procedures on liver|Procedure|false|false|C4037986;C1278929;C0023884|livernull|Abdomen>Liver|Anatomy|false|false|C3488428;C0459207;C0056632;C2702357;C5444130;C0457523;C1420285;C0007465;C0009213;C0028908;C1517288;C1947940;C3541397;C0872387;C0577060;C0023895;C0496870;C0721399;C0023899|liver
null|null|Anatomy|false|false|C3488428;C0459207;C0056632;C2702357;C5444130;C0457523;C1420285;C0007465;C0009213;C0028908;C1517288;C1947940;C3541397;C0872387;C0577060;C0023895;C0496870;C0721399;C0023899|liver
null|Liver|Anatomy|false|false|C3488428;C0459207;C0056632;C2702357;C5444130;C0457523;C1420285;C0007465;C0009213;C0028908;C1517288;C1947940;C3541397;C0872387;C0577060;C0023895;C0496870;C0721399;C0023899|livernull|oil ingredients|Drug|false|false|C4037986;C1278929;C0023884|oil
null|oil ingredients|Drug|false|false|C4037986;C1278929;C0023884|oil
null|Oil Dosage Form|Drug|false|false|C4037986;C1278929;C0023884|oil
null|Oils|Drug|false|false|C4037986;C1278929;C0023884|oil
null|Food Oil|Drug|false|false|C4037986;C1278929;C0023884|oilnull|UNK gene|Finding|false|false||unknull|Unknown|Modifier|false|false||unknull|Multivitamin preparation|Drug|false|false||Multivitamin
null|Multivitamin preparation|Drug|false|false||Multivitamin
null|Multivitamin preparation|Drug|false|false||Multivitaminnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|Acetaminophen [EPC]|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophennull|Acetaminophen measurement|Procedure|false|false||acetaminophennull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Every four hours|Time|false|false||Q4Hnull|Every - dosing instruction fragment|Finding|false|false||everynull|Every (qualifier)|Modifier|false|false||everynull|4 Hours|Time|false|false||4 hoursnull|Hour|Time|false|false||hoursnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|albuterol sulfate|Drug|false|false||albuterol sulfate
null|albuterol sulfate|Drug|false|false||albuterol sulfatenull|albuterol|Drug|false|false||albuterol
null|albuterol|Drug|false|false||albuterolnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfate
null|Sulfates, Inorganic|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfatenull|mcg/actuation|LabModifier|false|false||mcg/Actuationnull|microgram|LabModifier|false|false||mcgnull|Actuation (unit of presentation)|LabModifier|false|false||Actuationnull|Facial Hemiatrophy|Disorder|false|false||HFAnull|High frequency audiometry|Procedure|false|false||HFAnull|Inhalers, Aerosol|Device|false|false||Aerosol Inhalernull|Aerosol Dose Form|Drug|false|false||Aerosolnull|Aerosols|Device|false|false||Aerosolnull|Inhaler (unit of presentation)|Finding|false|false||Inhalernull|Inhaler|Device|false|false||Inhalernull|Inhaler Dosing Unit|LabModifier|false|false||Inhalernull|Puff Dosing Unit|LabModifier|false|false||Puff
null|Picofarad|LabModifier|false|false||Puffnull|Inhalation Route of Administration|Finding|false|false||Inhalation
null|Inspiration (function)|Finding|false|false||Inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||Inhalationnull|Every six hours|Time|false|false||Q6Hnull|6 Hours|Time|false|false||6 hoursnull|Hour|Time|false|false||hoursnull|Dyspnea|Finding|false|false||SOBnull|Wheezing|Finding|false|false||wheezenull|fluticasone / salmeterol|Drug|false|false||fluticasone-salmeterolnull|fluticasone|Drug|false|false||fluticasone
null|fluticasone|Drug|false|false||fluticasonenull|salmeterol|Drug|false|false||salmeterol
null|salmeterol|Drug|false|false||salmeterolnull|microgram|LabModifier|false|false||mcgnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Disk Drug Form|Drug|false|false|C1556138|Disknull|Disc - Body Part|Anatomy|false|false|C1550509;C0993608;C0034789|Disknull|Disk Device|Device|false|false||Disk
null|Disk - package|Device|false|false||Disknull|Disk Shape|Modifier|false|false||Disknull|Disk Dosing Unit|LabModifier|false|false||Disknull|Participation Type - device|Finding|false|false|C1556138|Devicenull|Medical Devices|Device|false|false||Device
null|Devices|Device|false|false||Devicenull|Kind of quantity - Device|LabModifier|false|false||Devicenull|Receptors, Antigen, B-Cell|Drug|false|false|C0262329|Sig
null|Receptors, Antigen, B-Cell|Drug|false|false|C0262329|Signull|Receptors, Antigen, B-Cell|Finding|false|false|C0262329;C1556138|Signull|Short insular gyrus|Anatomy|false|false|C0034789;C0034789|Signull|Surveillance Implementation Group|Entity|false|false||Sig
null|Staphylococcus intermedius group|Entity|false|false||Signull|Disk Drug Form|Drug|false|false|C1556138|Disknull|Disc - Body Part|Anatomy|false|false|C1550509;C4035627;C0004048;C0205535;C1332410;C0993608;C4546282;C1561538;C1561539|Disknull|Disk Device|Device|false|false||Disk
null|Disk - package|Device|false|false||Disknull|Disk Shape|Modifier|false|false||Disknull|Disk Dosing Unit|LabModifier|false|false||Disknull|Participation Type - device|Finding|false|false|C1556138|Devicenull|Medical Devices|Device|false|false||Device
null|Devices|Device|false|false||Devicenull|Kind of quantity - Device|LabModifier|false|false||Devicenull|Inhalation Route of Administration|Finding|false|false|C1556138|Inhalation
null|Inspiration (function)|Finding|false|false|C1556138|Inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||Inhalationnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false|C1556138|BIDnull|BID gene|Finding|false|false|C1556138|BIDnull|Twice a day|Time|false|false||BIDnull|2 times|Finding|false|false|C1556138|2 timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false|C1556138|day
null|Precision - day|Finding|false|false|C1556138|daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|fluticasone|Drug|false|false||fluticasone
null|fluticasone|Drug|false|false||fluticasonenull|mcg/actuation|LabModifier|false|false||mcg/Actuationnull|microgram|LabModifier|false|false||mcgnull|Actuation (unit of presentation)|LabModifier|false|false||Actuationnull|SPRAY, SUSPENSION|Drug|false|false||Spray, Suspensionnull|Spray Dosage Form|Drug|false|false||Spraynull|Spray (administration method)|Finding|false|false||Spraynull|Spray (action)|Event|false|false||Spraynull|Spray Dosing Unit|LabModifier|false|false||Spraynull|Suspension substance|Drug|false|false||Suspension
null|Suspensions|Drug|false|false||Suspensionnull|Suspension (action)|Finding|false|false||Suspensionnull|Nasal brand of oxymetazoline|Drug|false|false|C0028429|Nasal
null|Nasal brand of oxymetazoline|Drug|false|false|C0028429|Nasal
null|Nasal dosage form|Drug|false|false|C0028429|Nasalnull|Nasal Route of Administration|Finding|false|false|C0028429|Nasal
null|Nasal (intended site)|Finding|false|false|C0028429|Nasalnull|null|Anatomy|false|false|C4520890;C1522019;C1527304;C3539909;C0020517;C1547542;C0489531;C1314973;C0683368;C1457887;C1720092;C1272939;C0721966;C1561538;C1561539|Nasalnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false|C0028429|oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false|C0028429|day
null|Precision - day|Finding|false|false|C0028429|daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Allergy - Charge Type Reason|Finding|false|false|C0028429|allergy
null|Allergic disposition|Finding|false|false|C0028429|allergy
null|Hypersensitivity|Finding|false|false|C0028429|allergy
null|Response to antigens|Finding|false|false|C0028429|allergy
null|History of allergies|Finding|false|false|C0028429|allergy
null|Allergic Reaction|Finding|false|false|C0028429|allergynull|Allergy Specialty|Title|false|false||allergynull|Symptoms aspect|Finding|false|false|C0028429|symptoms
null|Symptoms|Finding|false|false|C0028429|symptomsnull|hydrochlorothiazide|Drug|false|false||hydrochlorothiazide
null|hydrochlorothiazide|Drug|false|false||hydrochlorothiazidenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|omeprazole|Drug|false|false||omeprazole
null|omeprazole|Drug|false|false||omeprazolenull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0030685;C0680255;C1963578;C0006935;C1283071;C0391871|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0030685;C0680255;C1963578;C0006935;C1283071;C0391871|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Delayed Release Dosage Form|Drug|false|false||Delayed Releasenull|Views delayed|Attribute|false|false||Delayednull|Deferred|Time|false|false||Delayednull|Release - action (qualifier value)|Finding|false|false|C0524463;C1325531|Release
null|Released (action)|Finding|false|false|C0524463;C1325531|Releasenull|Discharge (release)|Procedure|false|false|C0524463;C1325531|Release
null|Release (procedure)|Procedure|false|false|C0524463;C1325531|Release
null|Patient Discharge|Procedure|false|false|C0524463;C1325531|Releasenull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935;C1283071;C0391871;C0030685;C0680255;C1963578|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935;C1283071;C0391871;C0030685;C0680255;C1963578|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Delayed Release Dosage Form|Drug|false|false||Delayed Releasenull|Views delayed|Attribute|false|false||Delayednull|Deferred|Time|false|false||Delayednull|Release - action (qualifier value)|Finding|false|false|C0524463;C1325531|Release
null|Released (action)|Finding|false|false|C0524463;C1325531|Releasenull|Discharge (release)|Procedure|false|false|C0524463;C1325531|Release
null|Release (procedure)|Procedure|false|false|C0524463;C1325531|Release
null|Patient Discharge|Procedure|false|false|C0524463;C1325531|Releasenull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|simvastatin|Drug|false|false||simvastatin
null|simvastatin|Drug|false|false||simvastatinnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|tiotropium bromide|Drug|false|false||tiotropium bromide
null|tiotropium bromide|Drug|false|false||tiotropium bromidenull|tiotropium|Drug|false|false||tiotropium
null|tiotropium|Drug|false|false||tiotropiumnull|Bromides|Drug|false|false||bromidenull|Bromides measurement|Procedure|false|false|C0524463;C1325531|bromidenull|microgram|LabModifier|false|false||mcgnull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935;C0004048;C0205535;C0202341|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935;C0004048;C0205535;C0202341|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Inhalation Devices|Device|false|false||Inhalation Devicenull|Inhalation Route of Administration|Finding|false|false|C0524463;C1325531|Inhalation
null|Inspiration (function)|Finding|false|false|C0524463;C1325531|Inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||Inhalationnull|Participation Type - device|Finding|false|false||Devicenull|Medical Devices|Device|false|false||Device
null|Devices|Device|false|false||Devicenull|Kind of quantity - Device|LabModifier|false|false||Devicenull|capsule (pharmacologic)|Drug|false|false||Capnull|CATARACT, ANTERIOR POLAR|Disorder|false|false||Capnull|BRD4 wt Allele|Finding|false|false||Cap
null|HACD1 gene|Finding|false|false||Cap
null|SERPINB6 gene|Finding|false|false||Cap
null|BRD4 gene|Finding|false|false||Cap
null|CAP1 gene|Finding|false|false||Cap
null|SORBS1 gene|Finding|false|false||Cap
null|LNPEP gene|Finding|false|false||Capnull|CAP Regimen|Procedure|false|false||Cap
null|cisplatin/cyclophosphamide/doxorubicin protocol|Procedure|false|false||Cap
null|cyclophosphamide/doxorubicin/prednisone protocol|Procedure|false|false||Capnull|Cap (physical object)|Device|false|false||Cap
null|Syringe Caps|Device|false|false||Cap
null|Cap device|Device|false|false||Capnull|College of American Pathologists|Subject|false|false||Capnull|Controlled Attenuation Parameter|Modifier|false|false||Capnull|Capsule Dosing Unit|LabModifier|false|false||Capnull|Inhalation Route of Administration|Finding|false|false||Inhalation
null|Inspiration (function)|Finding|false|false||Inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||Inhalationnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|aspirin|Drug|false|false||aspirin
null|aspirin|Drug|false|false||aspirinnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Multivitamin tablet|Drug|false|false||multivitamin     Tabletnull|Multivitamin preparation|Drug|false|false||multivitamin
null|Multivitamin preparation|Drug|false|false||multivitamin
null|Multivitamin preparation|Drug|false|false||multivitaminnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|diltiazem hydrochloride|Drug|false|false||diltiazem HCl
null|diltiazem hydrochloride|Drug|false|false||diltiazem HClnull|diltiazem|Drug|false|false||diltiazem
null|diltiazem|Drug|false|false||diltiazemnull|Flinders medical centre-7 marker|Drug|false|false||HCl
null|hydrochloride|Drug|false|false||HCl
null|hydrochloride|Drug|false|false||HClnull|Hairy Cell Leukemia|Disorder|false|false||HClnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|refill|Finding|false|false||Refillsnull|nitroglycerin|Drug|false|false||nitroglycerin
null|nitroglycerin|Drug|false|false||nitroglycerinnull|Sublingual Tablet|Drug|false|false||Tablet, Sublingualnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Sublingual Route of Administration|Finding|false|false||Sublingual
null|Sublingual (intended site)|Finding|false|false||Sublingualnull|Sublingual location|Modifier|false|false||Sublingualnull|Receptors, Antigen, B-Cell|Drug|false|false|C0262329|Sig
null|Receptors, Antigen, B-Cell|Drug|false|false|C0262329|Signull|Receptors, Antigen, B-Cell|Finding|false|false|C0262329|Signull|Short insular gyrus|Anatomy|false|false|C0034789;C0034789|Signull|Surveillance Implementation Group|Entity|false|false||Sig
null|Staphylococcus intermedius group|Entity|false|false||Signull|Sublingual Route of Administration|Finding|false|false||Sublingual
null|Sublingual (intended site)|Finding|false|false||Sublingualnull|Sublingual location|Modifier|false|false||Sublingualnull|Minangkabau Language|Entity|false|false||minnull|Minute of time|Time|false|false||minnull|Minimum|Modifier|false|false||minnull|Minute Unit of Plane Angle|LabModifier|false|false||min
null|minim|LabModifier|false|false||minnull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C2926613;C0008031;C0741025|chest
null|Anterior thoracic region|Anatomy|false|false|C2926613;C0008031;C0741025|chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Onset of (contextual qualifier)|Modifier|false|false||onset ofnull|Onset of (contextual qualifier)|Modifier|false|false||onsetnull|Age of Onset|LabModifier|false|false||onsetnull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0008031;C2926613;C0741025;C1549543;C0030193|chest
null|Anterior thoracic region|Anatomy|false|false|C0008031;C2926613;C0741025;C1549543;C0030193|chestnull|Administration Method - Pain|Finding|false|false|C1527391;C0817096|pain
null|Pain|Finding|false|false|C1527391;C0817096|painnull|null|Attribute|false|false||painnull|Repeat Object|Finding|false|false||repeat
null|Repeat|Finding|false|false||repeatnull|Repeat Pattern|Time|false|false||repeatnull|Minangkabau Language|Entity|false|false||minnull|Minute of time|Time|false|false||minnull|Minimum|Modifier|false|false||minnull|Minute Unit of Plane Angle|LabModifier|false|false||min
null|minim|LabModifier|false|false||minnull|Continuous|Finding|false|false||continuednull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0741025;C2926613;C1549543;C0030193;C0008031|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025;C2926613;C1549543;C0030193;C0008031|chestnull|Administration Method - Pain|Finding|false|false|C1527391;C0817096|pain
null|Pain|Finding|false|false|C1527391;C0817096|painnull|null|Attribute|false|false||painnull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C1549543;C0030193;C0008031;C2926613;C0741025|chest
null|Anterior thoracic region|Anatomy|false|false|C1549543;C0030193;C0008031;C2926613;C0741025|chestnull|Administration Method - Pain|Finding|false|false|C1527391;C0817096|pain
null|Pain|Finding|false|false|C1527391;C0817096|painnull|null|Attribute|false|false||painnull|refill|Finding|false|false||Refillsnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Coronary Artery Disease|Disorder|false|false|C0226004;C0003842;C0205042;C0018787|Coronary Artery Disease
null|Coronary Arteriosclerosis|Disorder|false|false|C0226004;C0003842;C0205042;C0018787|Coronary Artery Diseasenull|Coronary artery|Anatomy|false|false|C1956346;C0010054;C0852949;C0012634|Coronary Arterynull|Heart|Anatomy|false|false|C0012634;C1956346;C0010054;C0852949|Coronarynull|Coronary|Modifier|false|false||Coronarynull|Arteriopathic disease|Disorder|false|false|C0226004;C0003842;C0205042;C0018787|Artery Diseasenull|Arterial system|Anatomy|false|false|C0852949;C1956346;C0010054;C0012634|Artery
null|Arteries|Anatomy|false|false|C0852949;C1956346;C0010054;C0012634|Arterynull|Disease|Disorder|false|false|C0018787;C0226004;C0003842;C0205042|Diseasenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Disease|Disorder|false|false||Conditionnull|Logical Condition|Finding|false|false||Conditionnull|null|Attribute|false|false||Conditionnull|Condition|Modifier|false|false||Conditionnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|Discharge instructions|Finding|false|false||Discharge Instructionsnull|hospital discharge instructions (treatment)|Procedure|false|false||Discharge Instructionsnull|null|Attribute|false|false||Discharge Instructionsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|Arm Pain|Finding|false|false|C0446516;C1140618;C1269078|arm painnull|Anorectal Malformations|Disorder|false|false|C0446516;C1140618;C1269078|armnull|AKR1A1 wt Allele|Finding|false|false|C0446516;C1140618;C1269078|arm
null|ARMC9 gene|Finding|false|false|C0446516;C1140618;C1269078|armnull|Protocol Treatment Arm|Procedure|false|false|C0446516;C1140618;C1269078|arm
null|Axillary Reverse Mapping|Procedure|false|false|C0446516;C1140618;C1269078|arm
null|Study Arm|Procedure|false|false|C0446516;C1140618;C1269078|armnull|Upper arm|Anatomy|false|false|C1549543;C0030193;C1522541;C5400986;C4761640;C1824218;C3715044;C0239377;C3495676|arm
null|null|Anatomy|false|false|C1549543;C0030193;C1522541;C5400986;C4761640;C1824218;C3715044;C0239377;C3495676|arm
null|Upper Extremity|Anatomy|false|false|C1549543;C0030193;C1522541;C5400986;C4761640;C1824218;C3715044;C0239377;C3495676|armnull|Administration Method - Pain|Finding|false|false|C0446516;C1140618;C1269078|pain
null|Pain|Finding|false|false|C0446516;C1140618;C1269078|painnull|null|Attribute|false|false||painnull|Heart Diseases|Disorder|false|false|C4037974;C0018787|heart diseasenull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C0018799;C0153957;C0153500;C0795691;C0012634|heart
null|Heart|Anatomy|false|false|C0018799;C0153957;C0153500;C0795691;C0012634|heartnull|Disease|Disorder|false|false|C4037974;C0018787|diseasenull|Tests (qualifier value)|Finding|false|false|C4318744|test
null|Testing|Finding|false|false|C4318744|testnull|Laboratory Procedures|Procedure|false|false|C4318744|testnull|Test - temporal region|Anatomy|false|false|C0456984;C0022885;C0039593;C0392366|testnull|Test Result|Lab|false|false|C4318744|testnull|Test Dosing Unit|LabModifier|false|false||testnull|Coronary Artery Disease|Disorder|false|false|C0226004;C0003842;C0205042;C0018787|coronary artery disease
null|Coronary Arteriosclerosis|Disorder|false|false|C0226004;C0003842;C0205042;C0018787|coronary artery diseasenull|Coronary artery|Anatomy|false|false|C1956346;C0010054;C0012634;C0852949|coronary arterynull|Heart|Anatomy|false|false|C0012634;C1956346;C0010054;C0852949|coronarynull|Coronary|Modifier|false|false||coronarynull|Arteriopathic disease|Disorder|false|false|C0205042;C0226004;C0003842;C0018787|artery diseasenull|Arterial system|Anatomy|false|false|C1956346;C0010054;C0012634;C0852949|artery
null|Arteries|Anatomy|false|false|C1956346;C0010054;C0012634;C0852949|arterynull|Disease|Disorder|false|false|C0226004;C0003842;C0205042;C0018787|diseasenull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Blood pressure finding|Finding|false|false||blood pressure
null|Systemic arterial pressure|Finding|false|false||blood pressure
null|Blood Pressure|Finding|false|false||blood pressurenull|Blood pressure determination|Procedure|false|false||blood pressurenull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Appointments|Event|false|false||appointmentsnull|Following|Time|false|false||following
null|Status post|Time|false|false||followingnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|diltiazem|Drug|false|false||Diltiazem
null|diltiazem|Drug|false|false||Diltiazemnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|To be stopped|Modifier|false|false||STOPPEDnull|theophylline|Drug|false|false||theophylline
null|theophylline|Drug|false|false||theophyllinenull|Assay of theophylline|Procedure|false|false||theophyllinenull|Started|Modifier|false|false||STARTEDnull|nitroglycerin|Drug|false|false||nitroglycerine
null|nitroglycerin|Drug|false|false||nitroglycerinenull|Have Chest Pain|Finding|false|false|C1527391;C0817096|have chest painnull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C2926613;C4054856;C0741025;C1549543;C0030193;C0008031|chest
null|Anterior thoracic region|Anatomy|false|false|C2926613;C4054856;C0741025;C1549543;C0030193;C0008031|chestnull|Administration Method - Pain|Finding|false|false|C1527391;C0817096|pain
null|Pain|Finding|false|false|C1527391;C0817096|painnull|null|Attribute|false|false||painnull|Stop brand of fluoride|Drug|false|false||STOP
null|Stop brand of fluoride|Drug|false|false||STOPnull|MAP6 gene|Finding|false|false||STOPnull|Stop (Instruction Imperative)|Event|false|false||STOPnull|Stop (qualifier value)|Time|false|false||STOPnull|Location characteristic ID - Smoking|Finding|false|false||SMOKING
null|Smoking|Finding|false|false||SMOKING
null|Tobacco smoking behavior|Finding|false|false||SMOKINGnull|kill - ActRelationshipJoin|Finding|false|false||KILL
null|Killing|Finding|false|false||KILL
null|Sacrifice|Finding|false|false||KILLnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions