 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|42,51|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|42,51|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|42,56|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|76,85|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|76,85|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|76,90|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|132,135|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|143,150|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|143,150|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Indicator, Reagent, or Diagnostic Aid|Allergies|184,187|false|false|false|C0013343|Dyes|Dye
Event|Event|Allergies|184,187|false|false|false|||Dye
Drug|Biologically Active Substance|Allergies|189,195|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Drug|Element, Ion, or Isotope|Allergies|189,195|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Drug|Pharmacologic Substance|Allergies|189,195|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Event|Activity|Allergies|196,206|false|false|false|C2700400|Contain (action)|Containing
Finding|Functional Concept|Allergies|196,206|false|false|false|C0332256|Containing (qualifier value)|Containing
Drug|Indicator, Reagent, or Diagnostic Aid|Allergies|207,215|false|false|false|C0009924|Contrast Media|Contrast
Drug|Indicator, Reagent, or Diagnostic Aid|Allergies|207,221|false|false|false|C0009924|Contrast Media|Contrast Media
Anatomy|Tissue|Allergies|216,221|false|false|false|C0162867;C1254021|Media layer;Tunica Media|Media
Finding|Intellectual Product|Allergies|216,221|false|false|false|C0009458;C0677540|Communications Media;PAMS Media|Media
Drug|Organic Chemical|Allergies|224,233|false|false|false|C0030049|oxycodone|Oxycodone
Drug|Pharmacologic Substance|Allergies|224,233|false|false|false|C0030049|oxycodone|Oxycodone
Event|Event|Allergies|224,233|false|false|false|||Oxycodone
Procedure|Laboratory Procedure|Allergies|224,233|false|false|false|C0524222|Oxycodone measurement|Oxycodone
Drug|Organic Chemical|Allergies|237,247|false|false|false|C0055729|cilostazol|cilostazol
Drug|Pharmacologic Substance|Allergies|237,247|false|false|false|C0055729|cilostazol|cilostazol
Event|Event|Allergies|237,247|false|false|false|||cilostazol
Drug|Organic Chemical|Allergies|250,261|false|false|false|C1569608|varenicline|Varenicline
Drug|Pharmacologic Substance|Allergies|250,261|false|false|false|C1569608|varenicline|Varenicline
Event|Event|Allergies|250,261|false|false|false|||Varenicline
Event|Event|Allergies|264,273|false|false|false|||Attending
Finding|Functional Concept|Allergies|264,273|false|false|false|C1999232|Attending (action)|Attending
Event|Event|Chief Complaint|299,308|false|false|false|||Shortness
Attribute|Clinical Attribute|Chief Complaint|299,318|false|false|false|C2707305||Shortness of breath
Finding|Sign or Symptom|Chief Complaint|299,318|false|false|false|C0013404|Dyspnea|Shortness of breath
Finding|Body Substance|Chief Complaint|312,318|false|false|false|C0225386|Breath|breath
Finding|Classification|Chief Complaint|321,326|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|327,335|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|327,335|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|339,357|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|348,357|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|348,357|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|348,357|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|348,357|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|348,357|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|Chief Complaint|359,369|false|false|false|||Intubation
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|359,369|false|false|false|C0021925|Intubation (procedure)|Intubation
Finding|Functional Concept|Chief Complaint|372,382|false|false|false|C0443254|mechanical method|Mechanical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|372,382|false|false|false|C0699886|Mechanical Treatments|Mechanical
Finding|Finding|Chief Complaint|372,394|false|false|false|C4760388|Mechanical ventilation finding|Mechanical Ventilation
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|372,394|false|false|false|C0199470|Mechanical ventilation|Mechanical Ventilation
Event|Event|Chief Complaint|383,394|false|false|false|||Ventilation
Finding|Physiologic Function|Chief Complaint|383,394|false|false|false|C0035203;C2945579|Respiration;Ventilation, function (observable entity)|Ventilation
Phenomenon|Phenomenon or Process|Chief Complaint|383,394|false|false|false|C0042491|Environmental air flow|Ventilation
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|383,394|false|false|false|C0554804|Assisted breathing|Ventilation
Event|Event|Chief Complaint|396,405|false|false|false|||Extubated
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|396,405|false|false|false|C0553891|Tracheal Extubation|Extubated
Finding|Idea or Concept|Chief Complaint|407,416|false|false|false|C1548539;C3245481|EntityNameUseR2 - temporary;Job Status - Temporary|Temporary
Finding|Intellectual Product|Chief Complaint|407,416|false|false|false|C1548539;C3245481|EntityNameUseR2 - temporary;Job Status - Temporary|Temporary
Finding|Gene or Genome|Chief Complaint|417,422|false|false|false|C3470541;C3890506|PACERR gene;RUBCNL gene|Pacer
Event|Event|Chief Complaint|423,432|false|false|false|||Placement
Procedure|Health Care Activity|Chief Complaint|423,432|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|Placement
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|423,432|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|Placement
Finding|Gene or Genome|Chief Complaint|433,436|false|false|false|C1421450;C2349087|EZR gene;EZR wt Allele|CVL
Event|Event|Chief Complaint|437,446|false|false|false|||Insertion
Finding|Functional Concept|Chief Complaint|437,446|false|false|false|C1512796;C1883719|Insert (object);Insertion Mutation|Insertion
Finding|Genetic Function|Chief Complaint|437,446|false|false|false|C1512796;C1883719|Insert (object);Insertion Mutation|Insertion
Procedure|Health Care Activity|Chief Complaint|437,446|false|false|false|C0021107;C0441587|Clinical act of insertion;Implantation procedure|Insertion
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|437,446|false|false|false|C0021107;C0441587|Clinical act of insertion;Implantation procedure|Insertion
Disorder|Disease or Syndrome|History of Present Illness|487,491|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|History of Present Illness|487,491|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|History of Present Illness|487,491|false|false|false|||COPD
Finding|Gene or Genome|History of Present Illness|487,491|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|History of Present Illness|505,513|false|false|false|||admitted
Disorder|Disease or Syndrome|History of Present Illness|516,521|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Event|Event|History of Present Illness|516,521|false|false|false|||times
Event|Event|History of Present Illness|537,544|false|false|false|||dyspnea
Finding|Finding|History of Present Illness|537,544|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|History of Present Illness|537,544|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Disorder|Disease or Syndrome|History of Present Illness|546,549|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|546,549|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|History of Present Illness|546,549|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|History of Present Illness|546,549|false|false|false|||CAD
Finding|Gene or Genome|History of Present Illness|546,549|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|History of Present Illness|546,549|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|History of Present Illness|546,549|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|546,549|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|551,557|false|false|false|C0018792|Heart Atrium|atrial
Attribute|Clinical Attribute|History of Present Illness|551,570|false|false|false|C2926591||atrial fibrillation
Disorder|Disease or Syndrome|History of Present Illness|551,570|false|false|false|C0004238|Atrial Fibrillation|atrial fibrillation
Lab|Laboratory or Test Result|History of Present Illness|551,570|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|atrial fibrillation
Disorder|Disease or Syndrome|History of Present Illness|558,570|false|false|false|C0232197|Fibrillation|fibrillation
Event|Event|History of Present Illness|558,570|false|false|false|||fibrillation
Drug|Organic Chemical|History of Present Illness|574,582|false|false|false|C1831808|apixaban|apixaban
Drug|Pharmacologic Substance|History of Present Illness|574,582|false|false|false|C1831808|apixaban|apixaban
Event|Event|History of Present Illness|574,582|false|false|false|||apixaban
Event|Event|History of Present Illness|587,596|false|false|false|||presented
Event|Event|History of Present Illness|603,612|false|false|false|||shortness
Attribute|Clinical Attribute|History of Present Illness|603,622|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|History of Present Illness|603,622|false|false|false|C0013404|Dyspnea|shortness of breath
Event|Event|History of Present Illness|616,622|false|false|false|||breath
Finding|Body Substance|History of Present Illness|616,622|false|false|false|C0225386|Breath|breath
Event|Event|History of Present Illness|635,645|false|false|false|||discharged
Event|Event|History of Present Illness|663,673|false|false|false|||discharged
Event|Event|History of Present Illness|674,678|false|false|false|||home
Finding|Idea or Concept|History of Present Illness|674,678|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|History of Present Illness|674,678|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|History of Present Illness|674,678|false|false|false|C1553498|home health encounter|home
Finding|Finding|History of Present Illness|674,692|false|false|false|C4534324|Home with services|home with services
Event|Event|History of Present Illness|684,692|false|false|false|||services
Event|Occupational Activity|History of Present Illness|684,692|false|false|false|C0557854|Services|services
Procedure|Health Care Activity|History of Present Illness|684,692|false|false|false|C1704289|Clinical Service|services
Finding|Idea or Concept|History of Present Illness|711,722|false|false|false|C0750502|Significant|significant
Disorder|Disease or Syndrome|History of Present Illness|723,727|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|History of Present Illness|723,727|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|History of Present Illness|723,727|false|false|false|||COPD
Finding|Gene or Genome|History of Present Illness|723,727|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|History of Present Illness|741,745|false|false|false|||PFTs
Event|Event|History of Present Illness|754,761|false|false|false|||showing
Finding|Finding|History of Present Illness|762,770|false|false|false|C0205082|Severe (severity modifier)|severely
Event|Event|History of Present Illness|771,778|false|false|false|||reduced
Finding|Finding|History of Present Illness|771,783|false|false|false|C5139283|Reduced forced expiratory volume in one second|reduced FEV1
Attribute|Clinical Attribute|History of Present Illness|779,783|false|false|false|C0802965||FEV1
Event|Event|History of Present Illness|779,783|false|false|false|||FEV1
Procedure|Diagnostic Procedure|History of Present Illness|779,783|false|false|false|C0849974|Pulmonary Function Test/Forced Expiratory Volume 1|FEV1
Finding|Finding|History of Present Illness|788,798|false|false|false|C4085643;C5201148;C5962468|Moderate;Moderate Effect;Moderate Response|moderately
Event|Event|History of Present Illness|799,806|false|false|false|||reduced
Finding|Finding|History of Present Illness|799,811|false|false|false|C5139283|Reduced forced expiratory volume in one second|reduced FEV1
Attribute|Clinical Attribute|History of Present Illness|807,811|false|false|false|C0802965||FEV1
Procedure|Diagnostic Procedure|History of Present Illness|807,811|false|false|false|C0849974|Pulmonary Function Test/Forced Expiratory Volume 1|FEV1
Attribute|Clinical Attribute|History of Present Illness|807,815|false|false|false|C0802741||FEV1/FVC
Procedure|Diagnostic Procedure|History of Present Illness|807,815|false|false|false|C3815113|Forced Expiratory Volume in 1 Second to Forced Vital Capacity Ratio Measurement|FEV1/FVC
Lab|Laboratory or Test Result|History of Present Illness|812,815|false|false|false|C3714541|Forced Vital Capacity|FVC
Event|Event|History of Present Illness|836,843|false|false|false|||feeling
Finding|Finding|History of Present Illness|836,850|false|false|false|C0424578|Psychological Well Being|feeling better
Event|Event|History of Present Illness|844,850|false|false|false|||better
Finding|Idea or Concept|History of Present Illness|844,850|false|false|false|C1550462|Observation Interpretation - better|better
Event|Event|History of Present Illness|857,867|false|false|false|||discharged
Event|Event|History of Present Illness|877,887|false|false|false|||continuing
Drug|Hormone|History of Present Illness|892,902|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|History of Present Illness|892,902|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|History of Present Illness|892,902|false|false|false|C0032952|prednisone|prednisone
Event|Event|History of Present Illness|892,902|false|false|false|||prednisone
Finding|Idea or Concept|History of Present Illness|929,932|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|History of Present Illness|929,932|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|History of Present Illness|943,955|false|false|false|||presentation
Finding|Idea or Concept|History of Present Illness|943,955|false|false|false|C0449450|Presentation|presentation
Event|Event|History of Present Illness|974,979|false|false|false|||began
Event|Event|History of Present Illness|983,989|false|false|false|||become
Event|Event|History of Present Illness|990,995|false|false|false|||short
Finding|Sign or Symptom|History of Present Illness|990,1005|false|false|false|C0013404|Dyspnea|short of breath
Finding|Body Substance|History of Present Illness|999,1005|false|false|false|C0225386|Breath|breath
Event|Event|History of Present Illness|1024,1032|false|false|false|||exertion
Finding|Organism Function|History of Present Illness|1024,1032|false|false|false|C0015264|Exertion|exertion
Event|Event|History of Present Illness|1038,1047|false|false|false|||developed
Drug|Organic Chemical|History of Present Illness|1050,1055|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|1050,1055|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|History of Present Illness|1050,1055|false|false|false|||cough
Finding|Sign or Symptom|History of Present Illness|1050,1055|false|false|false|C0010200|Coughing|cough
Finding|Finding|History of Present Illness|1050,1066|false|false|false|C0239134|Productive Cough|cough productive
Event|Event|History of Present Illness|1056,1066|false|false|false|||productive
Disorder|Disease or Syndrome|History of Present Illness|1071,1076|false|false|false|C0155339|Brown Tendon Sheath Syndrome|brown
Finding|Finding|History of Present Illness|1071,1083|false|false|false|C0457099|Brown sputum|brown sputum
Event|Event|History of Present Illness|1077,1083|false|false|false|||sputum
Finding|Body Substance|History of Present Illness|1077,1083|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Finding|Intellectual Product|History of Present Illness|1077,1083|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Event|Event|History of Present Illness|1088,1093|false|false|false|||fever
Finding|Finding|History of Present Illness|1088,1093|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|History of Present Illness|1088,1093|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|History of Present Illness|1095,1101|false|false|false|||chills
Finding|Sign or Symptom|History of Present Illness|1095,1101|true|false|false|C0085593|Chills|chills
Attribute|Clinical Attribute|History of Present Illness|1103,1109|false|false|false|C4255480||nausea
Event|Event|History of Present Illness|1103,1109|false|false|false|||nausea
Finding|Sign or Symptom|History of Present Illness|1103,1109|false|false|false|C0027497|Nausea|nausea
Event|Event|History of Present Illness|1111,1119|false|false|false|||vomiting
Finding|Sign or Symptom|History of Present Illness|1111,1119|false|false|false|C0042963|Vomiting|vomiting
Event|Event|History of Present Illness|1121,1129|false|false|false|||diarrhea
Finding|Finding|History of Present Illness|1121,1129|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|History of Present Illness|1121,1129|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Event|Event|History of Present Illness|1136,1142|false|false|false|||sleeps
Event|Event|History of Present Illness|1191,1197|false|false|false|||stable
Finding|Intellectual Product|History of Present Illness|1191,1197|false|false|false|C1547311|Patient Condition Code - Stable|stable
Disorder|Neoplastic Process|History of Present Illness|1204,1213|false|false|false|C0027627|Neoplasm Metastasis|secondary
Event|Event|History of Present Illness|1204,1213|false|false|false|||secondary
Finding|Functional Concept|History of Present Illness|1204,1213|false|false|false|C1522484|metastatic qualifier|secondary
Event|Event|History of Present Illness|1214,1221|false|false|false|||concern
Finding|Idea or Concept|History of Present Illness|1214,1221|false|false|false|C2699424|Concern|concern
Event|Event|History of Present Illness|1244,1251|false|false|false|||trouble
Event|Event|History of Present Illness|1252,1259|false|false|false|||walking
Finding|Functional Concept|History of Present Illness|1260,1263|false|false|false|C0678226;C3146286|Due;Due to|due
Finding|Idea or Concept|History of Present Illness|1260,1263|false|false|false|C0678226;C3146286|Due;Due to|due
Attribute|Clinical Attribute|History of Present Illness|1268,1272|false|false|false|C2598155||pain
Event|Event|History of Present Illness|1268,1272|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|1268,1272|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1268,1272|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1282,1285|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1282,1285|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|History of Present Illness|1282,1285|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|History of Present Illness|1282,1285|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Event|Event|History of Present Illness|1282,1285|false|false|false|||hip
Finding|Gene or Genome|History of Present Illness|1282,1285|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1282,1285|false|false|false|C1292890|Procedure on hip|hip
Anatomy|Body Location or Region|History of Present Illness|1291,1296|false|false|false|C0039866;C4299091|Lower extremity>Thigh;Thigh structure|thigh
Attribute|Clinical Attribute|History of Present Illness|1302,1308|false|false|false|C0944911||weight
Event|Event|History of Present Illness|1302,1308|false|false|false|||weight
Finding|Finding|History of Present Illness|1302,1308|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|History of Present Illness|1302,1308|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|History of Present Illness|1302,1308|false|false|false|C1305866|Weighing patient|weight
Event|Event|History of Present Illness|1309,1316|false|false|false|||bearing
Event|Event|History of Present Illness|1328,1331|false|false|false|||new
Finding|Finding|History of Present Illness|1328,1331|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|History of Present Illness|1328,1331|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Disorder|Injury or Poisoning|History of Present Illness|1336,1341|true|false|false|C0000921|Accidental Falls|falls
Event|Event|History of Present Illness|1336,1341|false|false|false|||falls
Finding|Finding|History of Present Illness|1336,1341|true|false|false|C0085639|Falls|falls
Disorder|Injury or Poisoning|History of Present Illness|1345,1351|true|false|false|C1368081;C3263723;C3714660|Physical trauma;Trauma;Traumatic injury|trauma
Event|Event|History of Present Illness|1345,1351|false|false|false|||trauma
Procedure|Health Care Activity|History of Present Illness|1345,1351|true|false|false|C0548346|Trauma assessment and care|trauma
Event|Event|History of Present Illness|1356,1360|false|false|false|||loss
Finding|Finding|History of Present Illness|1356,1360|true|false|false|C5890125|Loss (adaptation)|loss
Finding|Sign or Symptom|History of Present Illness|1356,1373|true|false|false|C0028643|Numbness|loss of sensation
Event|Event|History of Present Illness|1364,1373|false|false|false|||sensation
Finding|Finding|History of Present Illness|1364,1373|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|History of Present Illness|1364,1373|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|History of Present Illness|1364,1373|false|false|false|C2229507|sensory exam|sensation
Event|Event|History of Present Illness|1375,1383|false|false|false|||numbness
Finding|Finding|History of Present Illness|1375,1383|true|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|History of Present Illness|1375,1383|true|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Event|Event|History of Present Illness|1386,1394|false|false|false|||weakness
Finding|Sign or Symptom|History of Present Illness|1386,1394|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1396,1403|false|false|false|C0042027|Urinary tract|urinary
Finding|Body Substance|History of Present Illness|1407,1412|false|false|false|C0015733|Feces|fecal
Disorder|Disease or Syndrome|History of Present Illness|1407,1425|false|false|false|C0015732|Fecal Incontinence|fecal incontinence
Disorder|Disease or Syndrome|History of Present Illness|1413,1425|false|false|false|C0021167|Incontinence|incontinence
Event|Event|History of Present Illness|1413,1425|false|false|false|||incontinence
Event|Event|History of Present Illness|1429,1439|false|false|false|||difficulty
Finding|Finding|History of Present Illness|1429,1439|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Event|Event|History of Present Illness|1440,1449|false|false|false|||urinating
Finding|Idea or Concept|History of Present Illness|1467,1474|false|false|false|C1555582|Initial (abbreviation)|initial
Drug|Food|History of Present Illness|1475,1480|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|vital
Attribute|Clinical Attribute|History of Present Illness|1475,1486|false|false|false|C0488614;C0518766|Vital signs|vital signs
Procedure|Health Care Activity|History of Present Illness|1475,1486|false|false|false|C0150404|Taking vital signs|vital signs
Event|Event|History of Present Illness|1481,1486|false|false|false|||signs
Finding|Finding|History of Present Illness|1481,1486|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|History of Present Illness|1481,1486|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1515,1520|false|false|false|C0028429||Nasal
Drug|Biomedical or Dental Material|History of Present Illness|1515,1520|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Organic Chemical|History of Present Illness|1515,1520|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Pharmacologic Substance|History of Present Illness|1515,1520|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Finding|Finding|History of Present Illness|1515,1520|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Functional Concept|History of Present Illness|1515,1520|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1522,1529|false|false|false|C1550232|Body Parts - Cannula|Cannula
Finding|Body Substance|History of Present Illness|1522,1529|false|false|false|C1546577;C1550622|Specimen Type - Cannula|Cannula
Finding|Intellectual Product|History of Present Illness|1522,1529|false|false|false|C1546577;C1550622|Specimen Type - Cannula|Cannula
Event|Event|History of Present Illness|1535,1539|false|false|false|||Exam
Finding|Functional Concept|History of Present Illness|1535,1539|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|History of Present Illness|1535,1539|false|false|false|C0582103|Medical Examination|Exam
Event|Event|History of Present Illness|1544,1551|false|false|false|||notable
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1585,1588|false|false|false|C1261075|Structure of right lower lobe of lung|RLL
Finding|Finding|History of Present Illness|1585,1588|false|false|false|C5703311|Radiolucent Lines|RLL
Event|Event|History of Present Illness|1606,1610|false|false|false|||Labs
Lab|Laboratory or Test Result|History of Present Illness|1606,1610|false|false|false|C0587081|Laboratory test finding|Labs
Event|Event|History of Present Illness|1616,1623|false|false|false|||notable
Disorder|Disease or Syndrome|History of Present Illness|1629,1632|false|false|false|C0021400|Influenza|flu
Event|Event|History of Present Illness|1629,1632|false|false|false|||flu
Finding|Gene or Genome|History of Present Illness|1629,1632|false|false|false|C3811318|ZMYND10 wt Allele|flu
Drug|Biomedical or Dental Material|History of Present Illness|1633,1637|false|false|false|C0183753;C1706069|Swab Dosage Form;Swab specimen|swab
Drug|Substance|History of Present Illness|1633,1637|false|false|false|C0183753;C1706069|Swab Dosage Form;Swab specimen|swab
Event|Event|History of Present Illness|1633,1637|false|false|false|||swab
Procedure|Diagnostic Procedure|History of Present Illness|1633,1637|false|false|false|C0563454|Taking of swab|swab
Event|Event|History of Present Illness|1638,1646|false|false|false|||negative
Finding|Classification|History of Present Illness|1638,1646|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|History of Present Illness|1638,1646|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|History of Present Illness|1638,1646|false|false|false|C5237010|Expression Negative|negative
Anatomy|Cell|History of Present Illness|1648,1651|false|false|false|C0023516|Leukocytes|WBC
Finding|Functional Concept|History of Present Illness|1661,1665|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Functional Concept|History of Present Illness|1667,1672|false|false|false|C0333051|shift displacement|shift
Phenomenon|Phenomenon or Process|History of Present Illness|1667,1672|false|false|false|C2347509|Physical Shift|shift
Anatomy|Cell Component|History of Present Illness|1674,1677|false|false|false|C2263086|Nuclear cap binding complex location|CBC
Procedure|Laboratory Procedure|History of Present Illness|1674,1677|false|false|false|C0009555|Complete Blood Count|CBC
Event|Event|History of Present Illness|1688,1691|false|false|false|||WNL
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1693,1696|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Hormone|History of Present Illness|1693,1696|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Pharmacologic Substance|History of Present Illness|1693,1696|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Event|Event|History of Present Illness|1693,1696|false|false|false|||BNP
Finding|Gene or Genome|History of Present Illness|1693,1696|false|false|false|C1417808;C2982014|NPPB gene;NPPB wt Allele|BNP
Procedure|Laboratory Procedure|History of Present Illness|1693,1696|false|false|false|C1095989|Brain natriuretic peptide measurement|BNP
Drug|Organic Chemical|History of Present Illness|1702,1709|false|false|false|C0022924;C0376261|Lactates;lactate|lactate
Drug|Pharmacologic Substance|History of Present Illness|1702,1709|false|false|false|C0022924;C0376261|Lactates;lactate|lactate
Event|Event|History of Present Illness|1702,1709|false|false|false|||lactate
Procedure|Laboratory Procedure|History of Present Illness|1702,1709|false|false|false|C0202115|Lactic acid measurement|lactate
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1735,1742|false|false|false|C0033684|Proteins|protein
Drug|Biologically Active Substance|History of Present Illness|1735,1742|false|false|false|C0033684|Proteins|protein
Event|Event|History of Present Illness|1735,1742|false|false|false|||protein
Finding|Conceptual Entity|History of Present Illness|1735,1742|false|false|false|C1521746|Protein Info|protein
Procedure|Laboratory Procedure|History of Present Illness|1735,1742|false|false|false|C0202202|Protein measurement|protein
Event|Event|History of Present Illness|1757,1765|false|false|false|||negative
Finding|Classification|History of Present Illness|1757,1765|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|History of Present Illness|1757,1765|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|History of Present Illness|1757,1765|false|false|false|C5237010|Expression Negative|negative
Drug|Biologically Active Substance|History of Present Illness|1767,1770|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Drug|Inorganic Chemical|History of Present Illness|1767,1770|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Event|Event|History of Present Illness|1767,1770|false|false|false|||BUN
Procedure|Laboratory Procedure|History of Present Illness|1767,1770|false|false|false|C0005845|Blood urea nitrogen measurement|BUN
Event|Event|History of Present Illness|1783,1790|false|false|false|||Imaging
Finding|Finding|History of Present Illness|1783,1790|false|false|false|C0740845|Imaging problem|Imaging
Procedure|Diagnostic Procedure|History of Present Illness|1783,1790|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|Imaging
Event|Event|History of Present Illness|1792,1795|false|false|false|||CXR
Procedure|Diagnostic Procedure|History of Present Illness|1792,1795|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Intellectual Product|History of Present Illness|1801,1805|false|false|false|C1547225|Mild Severity of Illness Code|mild
Event|Event|History of Present Illness|1816,1827|false|false|false|||atelectasis
Finding|Pathologic Function|History of Present Illness|1816,1827|false|false|false|C0004144|Atelectasis|atelectasis
Event|Event|History of Present Illness|1851,1860|false|false|false|||concerned
Disorder|Disease or Syndrome|History of Present Illness|1865,1874|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|History of Present Illness|1865,1874|false|false|false|||pneumonia
Event|Event|History of Present Illness|1886,1890|false|false|false|||view
Finding|Body Substance|History of Present Illness|1900,1907|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1900,1907|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1900,1907|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1922,1932|false|false|false|C0042313|vancomycin|Vancomycin
Drug|Antibiotic|History of Present Illness|1922,1932|false|false|false|C0042313|vancomycin|Vancomycin
Event|Event|History of Present Illness|1922,1932|false|false|false|||Vancomycin
Procedure|Laboratory Procedure|History of Present Illness|1922,1932|false|false|false|C0489941|Vancomycin measurement|Vancomycin
Drug|Antibiotic|History of Present Illness|1937,1945|false|false|false|C0055003|cefepime|cefepime
Drug|Organic Chemical|History of Present Illness|1937,1945|false|false|false|C0055003|cefepime|cefepime
Event|Event|History of Present Illness|1937,1945|false|false|false|||cefepime
Drug|Antibiotic|History of Present Illness|1958,1970|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|History of Present Illness|1958,1970|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|History of Present Illness|1958,1970|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Event|Event|History of Present Illness|1958,1970|false|false|false|||azithromycin
Drug|Organic Chemical|History of Present Illness|1974,1980|false|false|false|C0939692|DuoNeb|duoneb
Drug|Pharmacologic Substance|History of Present Illness|1974,1980|false|false|false|C0939692|DuoNeb|duoneb
Event|Event|History of Present Illness|1974,1980|false|false|false|||duoneb
Drug|Hormone|History of Present Illness|1988,1998|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|History of Present Illness|1988,1998|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|History of Present Illness|1988,1998|false|false|false|C0032952|prednisone|prednisone
Finding|Idea or Concept|History of Present Illness|2017,2020|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|History of Present Illness|2017,2020|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|History of Present Illness|2028,2036|false|false|false|||Consults
Procedure|Health Care Activity|History of Present Illness|2028,2036|false|false|false|C0009818|Consultation|Consults
Event|Event|History of Present Illness|2046,2052|false|false|false|||Vitals
Event|Event|History of Present Illness|2062,2070|false|false|false|||transfer
Finding|Functional Concept|History of Present Illness|2062,2070|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|History of Present Illness|2062,2070|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|History of Present Illness|2062,2070|false|false|false|C4706767|Transfer (immobility management)|transfer
Event|Activity|History of Present Illness|2111,2118|false|false|false|C1706079||arrival
Event|Event|History of Present Illness|2111,2118|false|false|false|||arrival
Finding|Functional Concept|History of Present Illness|2111,2118|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Anatomy|Anatomical Structure|History of Present Illness|2126,2131|false|false|false|C3714591|Floor (anatomic)|floor
Event|Event|History of Present Illness|2142,2148|false|false|false|||stated
Attribute|Clinical Attribute|History of Present Illness|2153,2162|false|false|false|C5885990||breathing
Event|Event|History of Present Illness|2153,2162|false|false|false|||breathing
Finding|Finding|History of Present Illness|2153,2162|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|History of Present Illness|2153,2162|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|History of Present Illness|2153,2162|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|History of Present Illness|2153,2162|false|false|false|C1160636|respiratory system process|breathing
Event|Event|History of Present Illness|2177,2183|false|false|false|||better
Finding|Idea or Concept|History of Present Illness|2177,2183|false|false|false|C1550462|Observation Interpretation - better|better
Event|Event|History of Present Illness|2193,2202|false|false|false|||continued
Event|Event|History of Present Illness|2211,2220|false|false|false|||shortness
Event|Event|History of Present Illness|2225,2231|false|false|false|||breath
Finding|Body Substance|History of Present Illness|2225,2231|false|false|false|C0225386|Breath|breath
Event|Event|History of Present Illness|2237,2241|false|false|false|||felt
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2256,2260|false|false|false|C0013443;C0521421|Ear structure|ears
Finding|Gene or Genome|History of Present Illness|2256,2260|false|false|false|C1414437|EPRS1 gene|ears
Event|Event|History of Present Illness|2265,2272|false|false|false|||clogged
Finding|Finding|History of Present Illness|2298,2302|false|false|false|C5575035|Well (answer to question)|well
Event|Event|History of Present Illness|2308,2314|false|false|false|||stated
Event|Event|History of Present Illness|2328,2334|false|false|false|||taking
Attribute|Clinical Attribute|History of Present Illness|2343,2354|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|History of Present Illness|2343,2354|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|History of Present Illness|2343,2354|false|false|false|||medications
Finding|Intellectual Product|History of Present Illness|2343,2354|false|false|false|C4284232|Medications|medications
Event|Event|History of Present Illness|2359,2369|false|false|false|||prescribed
Disorder|Disease or Syndrome|Past Medical History|2399,2403|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Past Medical History|2399,2403|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Past Medical History|2399,2403|false|false|false|||COPD
Finding|Gene or Genome|Past Medical History|2399,2403|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|Past Medical History|2404,2410|false|false|false|C0004096|Asthma|Asthma
Event|Event|Past Medical History|2404,2410|false|false|false|||Asthma
Event|Event|Past Medical History|2414,2418|false|false|false|||home
Finding|Idea or Concept|Past Medical History|2414,2418|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Past Medical History|2414,2418|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Past Medical History|2414,2418|false|false|false|C1553498|home health encounter|home
Finding|Finding|Past Medical History|2427,2435|false|false|false|C0741302|atypia morphology|Atypical
Finding|Sign or Symptom|Past Medical History|2427,2446|false|false|false|C0262384|Atypical chest pain|Atypical Chest Pain
Anatomy|Body Location or Region|Past Medical History|2436,2441|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|Past Medical History|2436,2441|false|false|false|C0741025|Chest problem|Chest
Attribute|Clinical Attribute|Past Medical History|2436,2446|false|false|false|C2926613||Chest Pain
Finding|Sign or Symptom|Past Medical History|2436,2446|false|false|false|C0008031|Chest Pain|Chest Pain
Attribute|Clinical Attribute|Past Medical History|2442,2446|false|true|false|C2598155||Pain
Event|Event|Past Medical History|2442,2446|false|false|false|||Pain
Finding|Functional Concept|Past Medical History|2442,2446|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Past Medical History|2442,2446|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Disorder|Disease or Syndrome|Past Medical History|2449,2461|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|Past Medical History|2449,2461|false|false|false|||Hypertension
Disorder|Disease or Syndrome|Past Medical History|2464,2478|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|Hyperlipidemia
Event|Event|Past Medical History|2464,2478|false|false|false|||Hyperlipidemia
Finding|Finding|Past Medical History|2464,2478|false|false|false|C0428465|Serum lipids high (finding)|Hyperlipidemia
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2499,2505|false|false|false|C0018792|Heart Atrium|Atrial
Attribute|Clinical Attribute|Past Medical History|2499,2518|false|false|false|C2926591||Atrial Fibrillation
Disorder|Disease or Syndrome|Past Medical History|2499,2518|false|false|false|C0004238|Atrial Fibrillation|Atrial Fibrillation
Lab|Laboratory or Test Result|Past Medical History|2499,2518|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Atrial Fibrillation
Disorder|Disease or Syndrome|Past Medical History|2506,2518|false|false|false|C0232197|Fibrillation|Fibrillation
Event|Event|Past Medical History|2506,2518|false|false|false|||Fibrillation
Drug|Organic Chemical|Past Medical History|2522,2530|false|false|false|C1831808|apixaban|Apixaban
Drug|Pharmacologic Substance|Past Medical History|2522,2530|false|false|false|C1831808|apixaban|Apixaban
Disorder|Mental or Behavioral Dysfunction|Past Medical History|2533,2540|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|Anxiety
Event|Event|Past Medical History|2533,2540|false|false|false|||Anxiety
Finding|Sign or Symptom|Past Medical History|2533,2540|false|false|false|C0860603|Anxiety symptoms|Anxiety
Anatomy|Body Location or Region|Past Medical History|2543,2551|false|false|false|C0027530|Neck|Cervical
Disorder|Disease or Syndrome|Past Medical History|2543,2563|false|false|false|C0263884|Cervical radiculitis|Cervical Radiculitis
Disorder|Disease or Syndrome|Past Medical History|2552,2563|false|false|false|C0034544|Radiculitis|Radiculitis
Event|Event|Past Medical History|2552,2563|false|false|false|||Radiculitis
Anatomy|Body Location or Region|Past Medical History|2566,2574|false|false|false|C0027530|Neck|Cervical
Disorder|Disease or Syndrome|Past Medical History|2566,2586|false|false|false|C0158241;C1384641|Cervical spondylosis;Cervical spondylosis without myelopathy|Cervical Spondylosis
Disorder|Disease or Syndrome|Past Medical History|2575,2586|false|false|false|C0038019|Spondylosis|Spondylosis
Event|Event|Past Medical History|2575,2586|false|false|false|||Spondylosis
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2589,2597|false|false|false|C0018787|Heart|Coronary
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2589,2604|false|false|false|C0205042|Coronary artery|Coronary Artery
Disorder|Disease or Syndrome|Past Medical History|2589,2612|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|Coronary Artery Disease
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2598,2604|false|false|false|C0003842;C0226004|Arterial system;Arteries|Artery
Anatomy|Body System|Past Medical History|2598,2604|false|false|false|C0003842;C0226004|Arterial system;Arteries|Artery
Disorder|Disease or Syndrome|Past Medical History|2598,2612|false|false|false|C0852949|Arteriopathic disease|Artery Disease
Disorder|Disease or Syndrome|Past Medical History|2605,2612|false|false|false|C0012634|Disease|Disease
Event|Event|Past Medical History|2605,2612|false|false|false|||Disease
Finding|Sign or Symptom|Past Medical History|2615,2623|false|false|false|C0018681|Headache|Headache
Disorder|Disease or Syndrome|Past Medical History|2626,2632|false|false|false|C0019340;C0854331|Herpes simplex dermatitis|Herpes
Disorder|Disease or Syndrome|Past Medical History|2626,2639|false|false|false|C0019360;C0042338|Herpes zoster (disorder);herpesvirus 3, human|Herpes Zoster
Disorder|Virus|Past Medical History|2626,2639|false|false|false|C0019360;C0042338|Herpes zoster (disorder);herpesvirus 3, human|Herpes Zoster
Disorder|Disease or Syndrome|Past Medical History|2633,2639|false|false|false|C0019360|Herpes zoster (disorder)|Zoster
Event|Event|Past Medical History|2633,2639|false|false|false|||Zoster
Finding|Pathologic Function|Past Medical History|2642,2653|false|false|false|C0017181|Gastrointestinal Hemorrhage|GI Bleeding
Event|Event|Past Medical History|2645,2653|false|false|false|||Bleeding
Finding|Pathologic Function|Past Medical History|2645,2653|false|false|false|C0019080|Hemorrhage|Bleeding
Disorder|Disease or Syndrome|Past Medical History|2656,2683|false|false|false|C0085096|Peripheral Vascular Diseases|Peripheral Vascular Disease
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2667,2675|false|false|false|C0005847|Blood Vessel|Vascular
Disorder|Disease or Syndrome|Past Medical History|2667,2683|false|false|false|C0042373|Vascular Diseases|Vascular Disease
Disorder|Disease or Syndrome|Past Medical History|2676,2683|false|false|false|C0012634|Disease|Disease
Event|Event|Past Medical History|2676,2683|false|false|false|||Disease
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2698,2703|false|false|false|C0020889|Bone structure of ilium|iliac
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2698,2710|false|false|false|C0850459|iliac stents|iliac stents
Event|Event|Past Medical History|2704,2710|false|false|false|||stents
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2717,2720|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|Past Medical History|2717,2720|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|Past Medical History|2717,2720|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|Past Medical History|2717,2720|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|Past Medical History|2717,2720|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2717,2720|false|false|false|C1292890|Procedure on hip|hip
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2717,2732|false|false|false|C0392806|Prosthetic arthroplasty of hip (procedure)|hip replacement
Event|Event|Past Medical History|2721,2732|false|false|false|||replacement
Finding|Functional Concept|Past Medical History|2721,2732|false|false|false|C0559956|Replacement|replacement
Procedure|Health Care Activity|Past Medical History|2721,2732|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2721,2732|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Event|Event|Family Medical History|2771,2777|false|false|false|||Mother
Finding|Idea or Concept|Family Medical History|2771,2777|false|false|false|C1546508|Relationship - Mother|Mother
Disorder|Disease or Syndrome|Family Medical History|2783,2789|false|false|false|C0004096|Asthma|asthma
Event|Event|Family Medical History|2783,2789|false|false|false|||asthma
Disorder|Disease or Syndrome|Family Medical History|2794,2806|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|Family Medical History|2794,2806|false|false|false|||hypertension
Finding|Conceptual Entity|Family Medical History|2808,2814|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|Family Medical History|2808,2814|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2820,2825|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|Family Medical History|2820,2825|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|Family Medical History|2820,2825|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Finding|Finding|Family Medical History|2820,2825|false|false|false|C0750873|COLON PROBLEM|colon
Disorder|Neoplastic Process|Family Medical History|2820,2832|false|false|false|C0007102;C0346629;C0699790|Colon Carcinoma;Malignant neoplasm of large intestine;Malignant tumor of colon|colon cancer
Disorder|Neoplastic Process|Family Medical History|2826,2832|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Family Medical History|2826,2832|false|false|false|||cancer
Event|Event|Family Medical History|2835,2842|false|false|false|||Brother
Finding|Conceptual Entity|Family Medical History|2835,2842|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Idea or Concept|Family Medical History|2835,2842|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Disorder|Neoplastic Process|Family Medical History|2848,2856|false|false|false|C0023418|leukemia|leukemia
Event|Event|Family Medical History|2848,2856|false|false|false|||leukemia
Finding|Finding|General Exam|2876,2884|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|General Exam|2876,2884|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|General Exam|2876,2884|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|General Exam|2876,2896|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAMINATION
Procedure|Health Care Activity|General Exam|2876,2896|false|false|false|C0031809|Physical Examination|PHYSICAL EXAMINATION
Event|Activity|General Exam|2885,2896|false|false|false|C4321457|Examination|EXAMINATION
Event|Event|General Exam|2885,2896|false|false|false|||EXAMINATION
Procedure|Health Care Activity|General Exam|2885,2896|false|false|false|C0031809;C0582103|Medical Examination;Physical Examination|EXAMINATION
Procedure|Health Care Activity|General Exam|2900,2909|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|General Exam|2947,2953|false|false|false|||VITALS
Event|Event|General Exam|2983,2990|false|false|false|||GENERAL
Finding|Classification|General Exam|2983,2990|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|General Exam|2983,2990|false|false|false|C3812897|General medical service|GENERAL
Event|Event|General Exam|2992,3001|false|false|false|||breathing
Finding|Finding|General Exam|3002,3010|false|false|false|C2984079|Somewhat|somewhat
Event|Event|General Exam|3032,3038|false|false|false|||wheeze
Finding|Sign or Symptom|General Exam|3032,3038|false|false|false|C0043144|Wheezing|wheeze
Anatomy|Body Location or Region|General Exam|3042,3047|false|false|false|C1512338|HEENT|HEENT
Event|Event|General Exam|3053,3059|false|false|false|||pallor
Finding|Finding|General Exam|3053,3059|true|false|false|C0241137|Pallor of skin|pallor
Event|Event|General Exam|3063,3070|false|false|false|||icterus
Finding|Sign or Symptom|General Exam|3063,3070|true|false|false|C0022346|Icterus|icterus
Anatomy|Body Location or Region|General Exam|3075,3088|false|false|false|C0521367|Oropharyngeal|oropharyngeal
Disorder|Disease or Syndrome|General Exam|3075,3088|false|false|false|C0553694|Disorder of oropharynx|oropharyngeal
Finding|Functional Concept|General Exam|3075,3088|false|false|false|C1522409|Oropharyngeal Route of Administration|oropharyngeal
Disorder|Disease or Syndrome|General Exam|3075,3095|true|false|false|C4039409|Oropharyngeal lesion|oropharyngeal lesion
Event|Event|General Exam|3089,3095|false|false|false|||lesion
Finding|Finding|General Exam|3089,3095|true|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|General Exam|3089,3095|true|false|false|C0221198;C1546698|Lesion|lesion
Anatomy|Body Space or Junction|General Exam|3100,3105|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|General Exam|3100,3105|true|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|General Exam|3100,3105|true|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|General Exam|3100,3105|true|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Event|Event|General Exam|3107,3117|false|false|false|||tenderness
Finding|Mental Process|General Exam|3107,3117|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|General Exam|3107,3117|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Anatomy|Body Location or Region|General Exam|3121,3125|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|General Exam|3121,3125|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|General Exam|3121,3125|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|General Exam|3127,3133|false|false|false|||Supple
Finding|Functional Concept|General Exam|3127,3133|false|false|false|C0332254|Supple|Supple
Event|Event|General Exam|3135,3138|false|false|false|||JVP
Finding|Finding|General Exam|3135,3138|false|false|false|C0428897|Jugular venous pressure|JVP
Anatomy|Body Part, Organ, or Organ Component|General Exam|3147,3154|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|General Exam|3147,3154|false|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Event|General Exam|3156,3159|false|false|false|||RRR
Event|Event|General Exam|3161,3167|false|false|false|||unable
Finding|Finding|General Exam|3161,3167|false|false|false|C1299582|Unable|unable
Event|Event|General Exam|3171,3181|false|false|false|||appreciate
Event|Event|General Exam|3188,3189|false|false|false|||r
Event|Event|General Exam|3190,3191|false|false|false|||g
Attribute|Clinical Attribute|General Exam|3199,3208|false|false|false|C5885990||breathing
Event|Event|General Exam|3199,3208|false|false|false|||breathing
Finding|Finding|General Exam|3199,3208|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|General Exam|3199,3208|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|General Exam|3199,3208|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|General Exam|3199,3208|false|false|false|C1160636|respiratory system process|breathing
Anatomy|Body Part, Organ, or Organ Component|General Exam|3212,3221|false|false|false|C0024109|Lung|PULMONARY
Attribute|Clinical Attribute|General Exam|3212,3221|false|false|false|C2707265||PULMONARY
Finding|Finding|General Exam|3212,3221|false|false|false|C4522268|Pulmonary (intended site)|PULMONARY
Event|Event|General Exam|3231,3238|false|false|false|||wheezes
Finding|Sign or Symptom|General Exam|3231,3238|false|false|false|C0043144|Wheezing|wheezes
Event|Event|General Exam|3243,3249|false|false|false|||ronchi
Anatomy|Body Location or Region|General Exam|3253,3260|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|General Exam|3253,3260|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|General Exam|3253,3260|false|false|false|||ABDOMEN
Finding|Finding|General Exam|3253,3260|false|false|false|C0941288|Abdomen problem|ABDOMEN
Anatomy|Body Part, Organ, or Organ Component|General Exam|3276,3287|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Anatomy|Body Location or Region|General Exam|3292,3297|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|3292,3297|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|General Exam|3292,3307|false|false|false|C0023216|Lower Extremity|lower extremity
Finding|Pathologic Function|General Exam|3292,3313|false|false|false|C0239340|Edema of lower extremity|lower extremity edema
Anatomy|Body Part, Organ, or Organ Component|General Exam|3298,3307|false|false|false|C0015385|Limb structure|extremity
Finding|Pathologic Function|General Exam|3298,3313|false|false|false|C0085649|Peripheral edema|extremity edema
Attribute|Clinical Attribute|General Exam|3308,3313|false|false|false|C1717255||edema
Event|Event|General Exam|3308,3313|false|false|false|||edema
Finding|Pathologic Function|General Exam|3308,3313|false|false|false|C0013604|Edema|edema
Anatomy|Body Location or Region|General Exam|3317,3322|false|false|false|C0230444|Shin|shins
Finding|Body Substance|General Exam|3324,3331|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|General Exam|3324,3331|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|General Exam|3324,3331|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|General Exam|3336,3343|false|false|false|||sitting
Event|Event|General Exam|3348,3353|false|false|false|||style
Event|Event|General Exam|3367,3377|false|false|false|||appreciate
Event|Event|General Exam|3378,3388|false|false|false|||tenderness
Finding|Mental Process|General Exam|3378,3388|false|true|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|General Exam|3378,3388|false|true|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Anatomy|Body Part, Organ, or Organ Component|General Exam|3399,3402|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|General Exam|3399,3402|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|General Exam|3399,3402|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|General Exam|3399,3402|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|General Exam|3399,3402|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|General Exam|3399,3402|false|false|false|C1292890|Procedure on hip|hip
Anatomy|Body System|General Exam|3406,3410|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|General Exam|3406,3410|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|General Exam|3406,3410|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|General Exam|3406,3410|false|false|false|||SKIN
Finding|Body Substance|General Exam|3406,3410|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|General Exam|3406,3410|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Disorder|Disease or Syndrome|General Exam|3420,3424|false|false|false|C5779629|Eruption of skin (disorder)|rash
Event|Event|General Exam|3420,3424|false|false|false|||rash
Finding|Pathologic Function|General Exam|3420,3424|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|General Exam|3420,3424|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Event|Event|General Exam|3429,3439|false|false|false|||NEUROLOGIC
Event|Event|General Exam|3448,3454|false|false|false|||moving
Anatomy|Body Part, Organ, or Organ Component|General Exam|3455,3470|false|false|false|C0278454|All extremities|all extremities
Anatomy|Body Part, Organ, or Organ Component|General Exam|3459,3470|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Drug|Organic Chemical|General Exam|3476,3483|false|false|false|C1995603|PURPOSE (pharmacologic preparation)|purpose
Drug|Pharmacologic Substance|General Exam|3476,3483|false|false|false|C1995603|PURPOSE (pharmacologic preparation)|purpose
Event|Event|General Exam|3476,3483|false|false|false|||purpose
Finding|Functional Concept|General Exam|3476,3483|false|false|false|C1285529|Purpose|purpose
Finding|Finding|General Exam|3488,3496|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|General Exam|3488,3496|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|General Exam|3488,3496|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|General Exam|3488,3508|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAMINATION
Procedure|Health Care Activity|General Exam|3488,3508|false|false|false|C0031809|Physical Examination|PHYSICAL EXAMINATION
Event|Activity|General Exam|3497,3508|false|false|false|C4321457|Examination|EXAMINATION
Event|Event|General Exam|3497,3508|false|false|false|||EXAMINATION
Procedure|Health Care Activity|General Exam|3497,3508|false|false|false|C0031809;C0582103|Medical Examination;Physical Examination|EXAMINATION
Finding|Body Substance|General Exam|3512,3521|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|3512,3521|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|3512,3521|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|3512,3521|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|General Exam|3559,3561|false|false|false|||HR
Event|Event|General Exam|3569,3573|false|false|false|||went
Finding|Idea or Concept|General Exam|3585,3595|false|false|false|C0549178|Continuous|continuous
Event|Event|General Exam|3596,3605|false|false|false|||telemetry
Procedure|Diagnostic Procedure|General Exam|3596,3605|false|false|false|C0039451|Telemetry|telemetry
Finding|Body Substance|General Exam|3607,3614|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|General Exam|3607,3614|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|General Exam|3607,3614|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|General Exam|3624,3631|false|false|false|||respond
Event|Event|General Exam|3635,3640|false|false|false|||vocal
Finding|Functional Concept|General Exam|3635,3640|false|false|false|C0205382|vocal|vocal
Finding|Gene or Genome|General Exam|3644,3651|false|false|false|C1424619;C4761434|CD96 gene;CD96 wt Allele|tactile
Event|Event|General Exam|3652,3659|false|false|false|||stimuli
Phenomenon|Phenomenon or Process|General Exam|3652,3659|false|false|false|C0234402|Stimulus|stimuli
Anatomy|Body Part, Organ, or Organ Component|General Exam|3661,3667|false|false|false|C0034121|Pupil|Pupils
Event|Event|General Exam|3673,3685|false|false|false|||non-reactive
Drug|Amino Acid, Peptide, or Protein|General Exam|3690,3695|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|General Exam|3690,3695|false|false|false|C1570446|TNFSF14 protein, human|light
Event|Event|General Exam|3690,3695|false|false|false|||light
Finding|Finding|General Exam|3690,3695|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|General Exam|3690,3695|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|General Exam|3690,3695|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|General Exam|3690,3695|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|General Exam|3690,3695|false|false|false|C0031765|Phototherapy|light
Anatomy|Body Part, Organ, or Organ Component|General Exam|3708,3713|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|General Exam|3708,3713|true|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|General Exam|3708,3713|true|false|false|C0795691|HEART PROBLEM|heart
Anatomy|Body Location or Region|General Exam|3717,3721|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|General Exam|3717,3721|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|General Exam|3717,3721|true|false|false|C0024115|Lung diseases|lung
Finding|Finding|General Exam|3717,3721|true|false|false|C0740941|Lung Problem|lung
Attribute|Clinical Attribute|General Exam|3717,3728|true|false|false|C0035234|Respiratory Sounds|lung sounds
Event|Event|General Exam|3722,3728|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|General Exam|3722,3728|true|false|false|C0037709||sounds
Event|Event|General Exam|3748,3760|false|false|false|||auscultation
Procedure|Diagnostic Procedure|General Exam|3748,3760|false|false|false|C0004339|Auscultation|auscultation
Finding|Finding|General Exam|3770,3785|false|false|false|C3274944|Pronounced Dead|pronounced dead
Event|Event|General Exam|3781,3785|false|false|false|||dead
Finding|Finding|General Exam|3781,3785|false|false|false|C0011065;C1306577;C1546956|Cessation of life;Dead (finding);Death (finding)|dead
Finding|Organism Function|General Exam|3781,3785|false|false|false|C0011065;C1306577;C1546956|Cessation of life;Dead (finding);Death (finding)|dead
Event|Event|General Exam|3795,3801|false|false|false|||Family
Finding|Classification|General Exam|3795,3801|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|General Exam|3795,3801|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|General Exam|3795,3801|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|General Exam|3795,3801|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Event|Event|General Exam|3807,3815|false|false|false|||notified
Event|Event|General Exam|3837,3845|false|false|false|||declined
Procedure|Diagnostic Procedure|General Exam|3846,3856|false|false|false|C0004398|Autopsy|an autopsy
Event|Event|General Exam|3849,3856|false|false|false|||autopsy
Finding|Intellectual Product|General Exam|3849,3856|false|false|false|C1546546||autopsy
Procedure|Diagnostic Procedure|General Exam|3849,3856|false|false|false|C0004398;C1548821|Autopsy;Autopsy - Consent type|autopsy
Procedure|Health Care Activity|General Exam|3849,3856|false|false|false|C0004398;C1548821|Autopsy;Autopsy - Consent type|autopsy
Event|Event|General Exam|3880,3884|false|false|false|||LABS
Lab|Laboratory or Test Result|General Exam|3880,3884|false|false|false|C0587081|Laboratory test finding|LABS
Procedure|Health Care Activity|General Exam|3888,3897|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Disorder|Disease or Syndrome|General Exam|3930,3935|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3930,3935|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3930,3935|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|3936,3939|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|3944,3947|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|3944,3947|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|3944,3947|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|3953,3956|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|3953,3956|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|3953,3956|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|3953,3956|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|3962,3965|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|3962,3965|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|3971,3974|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|3971,3974|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|3971,3974|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|3971,3974|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|3971,3974|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|3979,3982|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|3979,3982|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|3979,3982|false|false|false|||MCH
Finding|Gene or Genome|General Exam|3979,3982|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|3979,3982|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|3979,3982|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|3988,3992|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|3988,3992|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|4021,4024|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|4041,4046|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4041,4046|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4041,4046|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Body Substance|General Exam|4059,4065|false|false|false|C0024202|Lymph|Lymphs
Drug|Antibiotic|General Exam|4071,4076|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|General Exam|4071,4076|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|General Exam|4071,4076|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|General Exam|4083,4086|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Event|Event|General Exam|4083,4086|false|false|false|||Eos
Finding|Gene or Genome|General Exam|4083,4086|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|General Exam|4189,4194|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4189,4194|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4189,4194|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|4195,4198|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|4215,4220|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4215,4220|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4215,4220|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|4215,4228|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|4215,4228|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|4215,4228|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|4221,4228|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|4221,4228|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|4221,4228|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|4221,4228|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|4221,4228|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|4221,4228|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|4274,4278|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|4274,4278|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|4274,4278|false|false|false|C0202059|Bicarbonate measurement|HCO3
Event|Event|General Exam|4278,4279|false|false|false|||-
Disorder|Disease or Syndrome|General Exam|4303,4308|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4303,4308|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4303,4308|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|4309,4312|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|4309,4312|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|General Exam|4309,4312|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|General Exam|4309,4312|false|false|false|||ALT
Finding|Gene or Genome|General Exam|4309,4312|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|General Exam|4309,4312|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|General Exam|4309,4312|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|General Exam|4309,4312|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|General Exam|4317,4320|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|General Exam|4317,4320|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|4317,4320|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|General Exam|4317,4320|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|General Exam|4317,4320|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Finding|Gene or Genome|General Exam|4317,4320|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|4325,4332|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|General Exam|4325,4332|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|General Exam|4360,4365|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4360,4365|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4360,4365|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|4366,4372|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Drug|Hormone|General Exam|4366,4372|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Disorder|Disease or Syndrome|General Exam|4389,4394|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4389,4394|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4389,4394|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|4389,4402|false|false|false|C0853248|Blood albumin|BLOOD Albumin
Drug|Amino Acid, Peptide, or Protein|General Exam|4395,4402|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Biologically Active Substance|General Exam|4395,4402|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Pharmacologic Substance|General Exam|4395,4402|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Event|Event|General Exam|4395,4402|false|false|false|||Albumin
Finding|Gene or Genome|General Exam|4395,4402|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Finding|Physiologic Function|General Exam|4395,4402|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Procedure|Laboratory Procedure|General Exam|4395,4402|false|false|false|C0201838|Albumin measurement|Albumin
Drug|Biologically Active Substance|General Exam|4407,4414|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|4407,4414|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|4407,4414|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|4407,4414|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|4407,4414|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|General Exam|4407,4414|false|false|false|||Calcium
Finding|Physiologic Function|General Exam|4407,4414|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|4407,4414|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|General Exam|4448,4453|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4448,4453|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4448,4453|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Event|General Exam|4458,4461|false|false|false|||pO2
Finding|Classification|General Exam|4458,4461|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|pO2
Finding|Molecular Function|General Exam|4458,4461|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|pO2
Procedure|Laboratory Procedure|General Exam|4458,4461|false|false|false|C1283004|PO2 measurement|pO2
Lab|Laboratory or Test Result|General Exam|4467,4471|false|false|false|C0391839|Carbon dioxide, partial pressure|pCO2
Procedure|Laboratory Procedure|General Exam|4467,4471|false|false|false|C0201931|Carbon dioxide measurement, partial pressure|pCO2
Anatomy|Body Location or Region|General Exam|4495,4499|false|false|false|C2987514|Anatomical base|Base
Drug|Biomedical or Dental Material|General Exam|4495,4499|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Drug|Chemical Viewed Functionally|General Exam|4495,4499|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|4495,4499|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Finding|Gene or Genome|General Exam|4495,4499|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|Base
Finding|Idea or Concept|General Exam|4495,4499|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|Base
Finding|Intellectual Product|General Exam|4505,4512|false|false|false|C0282411;C0947611|Comment;Published Comment|Comment
Event|Event|General Exam|4519,4522|false|false|false|||TOP
Disorder|Disease or Syndrome|General Exam|4535,4540|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4535,4540|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4535,4540|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|4535,4548|false|false|false|C3824990|lactate in blood (lab test)|BLOOD Lactate
Drug|Organic Chemical|General Exam|4541,4548|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Drug|Pharmacologic Substance|General Exam|4541,4548|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Event|Event|General Exam|4541,4548|false|false|false|||Lactate
Procedure|Laboratory Procedure|General Exam|4541,4548|false|false|false|C0202115|Lactic acid measurement|Lactate
Event|Event|General Exam|4555,4559|false|false|false|||LABS
Lab|Laboratory or Test Result|General Exam|4555,4559|false|false|false|C0587081|Laboratory test finding|LABS
Finding|Body Substance|General Exam|4563,4572|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|4563,4572|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|4563,4572|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|4563,4572|false|false|false|C0030685|Patient Discharge|DISCHARGE
Disorder|Disease or Syndrome|General Exam|4605,4610|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4605,4610|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4605,4610|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|4611,4614|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|4621,4624|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|4621,4624|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|4621,4624|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|4631,4634|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|4631,4634|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|4631,4634|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|4631,4634|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|4640,4643|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|4640,4643|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|4651,4654|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|4651,4654|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|4651,4654|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|4651,4654|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|4651,4654|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|4658,4661|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|4658,4661|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|4658,4661|false|false|false|||MCH
Finding|Gene or Genome|General Exam|4658,4661|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|4658,4661|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|4658,4661|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|4667,4671|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|4667,4671|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|4700,4703|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|4720,4725|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4720,4725|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4720,4725|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|4720,4733|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|4720,4733|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|4720,4733|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|4726,4733|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|4726,4733|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|4726,4733|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|4726,4733|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|4726,4733|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|4726,4733|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|4776,4780|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|4776,4780|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|4776,4780|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|4805,4810|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4805,4810|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4805,4810|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|4805,4818|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|General Exam|4811,4818|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|4811,4818|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|4811,4818|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|4811,4818|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|4811,4818|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|General Exam|4811,4818|false|false|false|||Calcium
Finding|Physiologic Function|General Exam|4811,4818|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|4811,4818|false|false|false|C0201925|Calcium measurement|Calcium
Event|Activity|General Exam|4841,4847|false|false|false|C1707391|Choose (action)|SELECT
Event|Event|General Exam|4841,4847|false|false|false|||SELECT
Procedure|Research Activity|General Exam|4841,4847|false|false|false|C1519229|Selenium and Vitamin E Efficacy Trial|SELECT
Event|Event|General Exam|4848,4855|false|false|false|||IMAGING
Finding|Finding|General Exam|4848,4855|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|General Exam|4848,4855|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Event|Event|General Exam|4877,4880|false|false|false|||CXR
Procedure|Diagnostic Procedure|General Exam|4877,4880|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Activity|General Exam|4884,4894|false|false|false|C1707455|Comparison|COMPARISON
Event|Event|General Exam|4884,4894|false|false|false|||COMPARISON
Anatomy|Body Part, Organ, or Organ Component|Findings|4915,4920|false|false|false|C0018787;C4037974|Chest>Heart;Heart|Heart
Disorder|Neoplastic Process|Findings|4915,4920|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|Heart
Finding|Sign or Symptom|Findings|4915,4920|false|false|false|C0795691|HEART PROBLEM|Heart
Finding|Finding|Findings|4915,4925|false|false|false|C0744689|heart size|Heart size
Event|Event|Findings|4921,4925|false|false|false|||size
Finding|Finding|Findings|4929,4944|false|false|false|C5425894|Mildly enlarged|mildly enlarged
Event|Event|Findings|4936,4944|false|false|false|||enlarged
Finding|Intellectual Product|Findings|4955,4959|false|false|false|C1547225|Mild Severity of Illness Code|mild
Event|Event|Findings|4960,4969|false|false|false|||unfolding
Anatomy|Body Location or Region|Findings|4978,4986|false|false|false|C0817096|Chest|thoracic
Disorder|Disease or Syndrome|Findings|4978,4986|false|false|false|C5779551|Dissecting Thoracic Aortic Aneurysm|thoracic
Anatomy|Body Part, Organ, or Organ Component|Findings|4978,4992|false|false|false|C1522460;C4037977|Chest>Aorta.thoracic;Thoracic aorta|thoracic aorta
Anatomy|Body Part, Organ, or Organ Component|Findings|4987,4992|false|false|false|C0003483;C4037978|Aorta;Chest+Abdomen>Aorta|aorta
Event|Event|Findings|4987,4992|false|false|false|||aorta
Procedure|Health Care Activity|Findings|4987,4992|false|false|false|C0869784|Procedure on aorta|aorta
Event|Event|Findings|5012,5022|false|false|false|||silhouette
Event|Event|Findings|5033,5041|false|false|false|||contours
Event|Event|Findings|5057,5069|false|false|false|||unremarkable
Finding|Intellectual Product|Findings|5080,5084|false|false|false|C1547225|Mild Severity of Illness Code|mild
Event|Event|Findings|5095,5106|false|false|false|||atelectasis
Finding|Pathologic Function|Findings|5095,5106|false|false|false|C0004144|Atelectasis|atelectasis
Anatomy|Body Part, Organ, or Organ Component|Findings|5109,5114|false|false|false|C0024109|Lung|Lungs
Event|Event|Findings|5129,5134|false|false|false|||clear
Finding|Idea or Concept|Findings|5129,5134|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Tissue|Findings|5136,5143|false|false|false|C0032225|Pleura|Pleural
Disorder|Disease or Syndrome|Findings|5136,5143|false|false|false|C0032226|Pleural Diseases|Pleural
Event|Event|Findings|5144,5152|false|false|false|||surfaces
Event|Event|Findings|5157,5162|false|false|false|||clear
Finding|Idea or Concept|Findings|5157,5162|false|false|false|C1550016|Remote control command - Clear|clear
Event|Event|Findings|5172,5180|false|false|false|||effusion
Finding|Body Substance|Findings|5172,5180|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|Findings|5172,5180|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|Findings|5172,5180|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Disorder|Disease or Syndrome|Findings|5184,5196|false|false|false|C0032326|Pneumothorax|pneumothorax
Event|Event|Findings|5184,5196|false|false|false|||pneumothorax
Event|Event|Findings|5198,5203|false|false|false|||Focus
Finding|Functional Concept|Findings|5198,5203|false|false|false|C1285542|Has focus|Focus
Drug|Inorganic Chemical|Findings|5207,5210|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|Findings|5207,5210|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|Findings|5207,5210|false|false|false|C0001861;C3536832|Air (substance);air|air
Event|Event|Findings|5207,5210|false|false|false|||air
Finding|Finding|Findings|5207,5210|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|Findings|5207,5210|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|Findings|5207,5210|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Event|Event|Findings|5211,5215|false|false|false|||seen
Finding|Functional Concept|Findings|5226,5231|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|Findings|5233,5246|false|false|false|C1269845|Structure of hemidiaphragm|hemidiaphragm
Finding|Finding|Findings|5248,5254|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Findings|5248,5254|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|Findings|5255,5265|false|false|false|||represents
Anatomy|Body Part, Organ, or Organ Component|Findings|5266,5273|false|false|false|C0009368|Colon structure (body structure)|colonic
Procedure|Therapeutic or Preventive Procedure|Findings|5266,5287|false|true|false|C0399644|Excision of large intestine for interposition|colonic interposition
Event|Event|Findings|5274,5287|false|false|false|||interposition
Event|Event|Findings|5291,5301|false|false|false|||IMPRESSION
Finding|Intellectual Product|Findings|5291,5301|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|Findings|5291,5301|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Intellectual Product|Findings|5305,5310|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Location or Region|Findings|5311,5326|false|false|false|C0553534|Cardiopulmonary|cardiopulmonary
Disorder|Disease or Syndrome|Findings|5311,5326|false|false|false|C4072686|Cardiovascular disease+Pulmonary disease|cardiopulmonary
Disorder|Congenital Abnormality|Findings|5327,5338|true|false|false|C0000768|Congenital Abnormality|abnormality
Event|Event|Findings|5327,5338|false|false|false|||abnormality
Finding|Finding|Findings|5327,5338|true|false|false|C1704258|Abnormality|abnormality
Drug|Organic Chemical|Findings|5347,5350|false|false|false|C0939812|Ruta graveolens preparation|RUE
Drug|Pharmacologic Substance|Findings|5347,5350|false|false|false|C0939812|Ruta graveolens preparation|RUE
Event|Event|Findings|5347,5350|false|false|false|||RUE
Event|Event|Findings|5357,5367|false|false|false|||IMPRESSION
Finding|Intellectual Product|Findings|5357,5367|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|Findings|5357,5367|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Intellectual Product|Findings|5374,5379|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Attribute|Clinical Attribute|Findings|5380,5384|false|false|false|C4318566|Deep Resection Margin|deep
Anatomy|Body Part, Organ, or Organ Component|Findings|5380,5389|false|false|false|C0226514|Structure of deep vein|deep vein
Disorder|Disease or Syndrome|Findings|5380,5400|false|false|false|C0149871;C0340708|Deep Vein Thrombosis;Deep vein thrombosis of lower limb|deep vein thrombosis
Anatomy|Body Part, Organ, or Organ Component|Findings|5385,5389|false|false|false|C0042449|Veins|vein
Finding|Pathologic Function|Findings|5385,5400|false|false|false|C0042487|Venous Thrombosis|vein thrombosis
Event|Event|Findings|5390,5400|false|false|false|||thrombosis
Finding|Pathologic Function|Findings|5390,5400|false|false|false|C0040053|Thrombosis|thrombosis
Event|Event|Findings|5401,5406|false|false|false|||noted
Finding|Functional Concept|Findings|5423,5428|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|Findings|5429,5442|false|false|false|C0226812|Structure of brachial vein|brachial vein
Anatomy|Body Part, Organ, or Organ Component|Findings|5438,5442|false|false|false|C0042449|Veins|vein
Finding|Idea or Concept|Findings|5455,5460|false|false|false|C1552828|Table Frame - above|above
Event|Event|Findings|5468,5471|false|false|false|||CXR
Procedure|Diagnostic Procedure|Findings|5468,5471|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|Findings|5474,5484|false|false|false|||IMPRESSION
Finding|Intellectual Product|Findings|5474,5484|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|Findings|5474,5484|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Functional Concept|Findings|5503,5507|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Finding|Gene or Genome|Findings|5503,5507|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Event|Event|Findings|5508,5511|false|false|false|||tip
Finding|Gene or Genome|Findings|5508,5511|false|false|false|C1705504;C1823282;C1825626;C1825978|ITFG1 gene;KAT5 wt Allele;METTL8 gene;TIPRL gene|tip
Procedure|Therapeutic or Preventive Procedure|Findings|5508,5511|false|false|false|C0673828|TIP regimen|tip
Anatomy|Body Part, Organ, or Organ Component|Findings|5530,5536|false|false|false|C0225594;C4521147|Keel structure;Structure of carina|carina
Anatomy|Body Location or Region|Findings|5540,5551|false|false|false|C3282907|Nasogastric|Nasogastric
Finding|Functional Concept|Findings|5540,5551|false|false|false|C0694637|Nasogastric Route of Administration|Nasogastric
Procedure|Therapeutic or Preventive Procedure|Findings|5540,5556|false|false|false|C0812428|Nasogastric tube procedures|Nasogastric tube
Event|Event|Findings|5552,5556|false|false|false|||tube
Finding|Functional Concept|Findings|5552,5556|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Finding|Gene or Genome|Findings|5552,5556|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Event|Event|Findings|5557,5560|false|false|false|||tip
Finding|Gene or Genome|Findings|5557,5560|false|false|false|C1705504;C1823282;C1825626;C1825978|ITFG1 gene;KAT5 wt Allele;METTL8 gene;TIPRL gene|tip
Procedure|Therapeutic or Preventive Procedure|Findings|5557,5560|false|false|false|C0673828|TIP regimen|tip
Finding|Conceptual Entity|Findings|5599,5603|false|false|false|C2697523|Graph Edge|edge
Drug|Biomedical or Dental Material|Findings|5612,5616|false|false|false|C1561572;C1704608|Film Dosage Form;film - layer|film
Drug|Substance|Findings|5612,5616|false|false|false|C1561572;C1704608|Film Dosage Form;film - layer|film
Event|Event|Findings|5612,5616|false|false|false|||film
Finding|Intellectual Product|Findings|5612,5616|false|false|false|C4019020||film
Finding|Functional Concept|Findings|5621,5625|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Drug|Pharmacologic Substance|Findings|5626,5633|false|false|false|C0719205|Central brand of multivitamin with minerals|central
Drug|Vitamin|Findings|5626,5633|false|false|false|C0719205|Central brand of multivitamin with minerals|central
Procedure|Laboratory Procedure|Findings|5626,5633|false|false|false|C1879652|Central Minus|central
Drug|Biologically Active Substance|Findings|5634,5638|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Findings|5634,5638|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Substance|Findings|5634,5638|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Event|Event|Findings|5634,5638|false|false|false|||line
Finding|Intellectual Product|Findings|5634,5638|false|false|false|C1546701|line source specimen code|line
Event|Event|Findings|5642,5649|false|false|false|||present
Finding|Finding|Findings|5642,5649|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|Findings|5642,5649|false|false|false|C0150312;C0449450|Present;Presentation|present
Event|Event|Findings|5657,5660|false|false|false|||tip
Finding|Gene or Genome|Findings|5657,5660|false|false|false|C1705504;C1823282;C1825626;C1825978|ITFG1 gene;KAT5 wt Allele;METTL8 gene;TIPRL gene|tip
Procedure|Therapeutic or Preventive Procedure|Findings|5657,5660|false|false|false|C0673828|TIP regimen|tip
Event|Event|Findings|5676,5679|false|false|false|||SVC
Finding|Finding|Findings|5676,5679|false|false|false|C0231957|Slow vital capacity|SVC
Event|Event|Findings|5684,5693|false|false|false|||pacemaker
Finding|Intellectual Product|Findings|5684,5693|false|false|false|C1546728||pacemaker
Event|Event|Findings|5697,5702|false|false|false|||noted
Event|Event|Findings|5710,5715|false|false|false|||right
Finding|Functional Concept|Findings|5710,5715|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Drug|Element, Ion, or Isotope|Findings|5723,5727|false|false|false|C0023175;C1442948|Plumbum metallicum, homeopathic preparation;lead|lead
Drug|Hazardous or Poisonous Substance|Findings|5723,5727|false|false|false|C0023175;C1442948|Plumbum metallicum, homeopathic preparation;lead|lead
Drug|Inorganic Chemical|Findings|5723,5727|false|false|false|C0023175;C1442948|Plumbum metallicum, homeopathic preparation;lead|lead
Drug|Pharmacologic Substance|Findings|5723,5727|false|false|false|C0023175;C1442948|Plumbum metallicum, homeopathic preparation;lead|lead
Event|Event|Findings|5723,5727|false|false|false|||lead
Finding|Functional Concept|Findings|5723,5727|false|false|false|C1522538|Leading|lead
Procedure|Diagnostic Procedure|Findings|5723,5727|false|false|false|C0524167;C5575683|Lead measurement;Long Ensemble Angular-Coherence Doppler Ultrasound|lead
Procedure|Laboratory Procedure|Findings|5723,5727|false|false|false|C0524167;C5575683|Lead measurement;Long Ensemble Angular-Coherence Doppler Ultrasound|lead
Event|Event|Findings|5729,5737|false|false|false|||projects
Finding|Functional Concept|Findings|5747,5752|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|Findings|5747,5762|false|false|false|C0225883|Right ventricular structure|right ventricle
Anatomy|Body Part, Organ, or Organ Component|Findings|5753,5762|false|false|false|C0007799;C0018827;C2355627|Cerebral Ventricles;Heart Ventricle;Ventricle|ventricle
Anatomy|Body Space or Junction|Findings|5753,5762|false|false|false|C0007799;C0018827;C2355627|Cerebral Ventricles;Heart Ventricle;Ventricle|ventricle
Finding|Finding|Findings|5774,5782|false|false|false|C0332148|Probable diagnosis|probable
Event|Event|Findings|5783,5791|false|false|false|||scarring
Finding|Pathologic Function|Findings|5783,5791|false|true|false|C0008767;C2004491|Cicatrix;Cicatrization|scarring
Anatomy|Body Location or Region|Findings|5801,5805|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Findings|5801,5805|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Findings|5801,5805|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Findings|5801,5805|false|false|false|C0740941|Lung Problem|lung
Event|Event|Findings|5806,5812|false|false|false|||apices
Finding|Finding|Findings|5828,5831|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Findings|5828,5831|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Event|Event|Findings|5832,5837|false|false|false|||areas
Disorder|Disease or Syndrome|Findings|5841,5854|false|false|false|C0521530|Lung consolidation|consolidation
Event|Event|Findings|5841,5854|false|false|false|||consolidation
Event|Event|Findings|5878,5892|false|false|false|||redistribution
Finding|Functional Concept|Findings|5878,5892|false|false|false|C0332620|Redistribution|redistribution
Event|Event|Findings|5897,5909|false|false|false|||cardiomegaly
Finding|Finding|Findings|5897,5909|false|false|false|C0018800|Cardiomegaly|cardiomegaly
Event|Event|Findings|5910,5920|false|false|false|||suggesting
Anatomy|Body Part, Organ, or Organ Component|Findings|5922,5931|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Findings|5922,5931|false|false|false|C2707265||pulmonary
Finding|Finding|Findings|5922,5931|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|Findings|5922,5951|false|false|false|C4477098|Pulmonary venous hypertension|pulmonary venous hypertension
Anatomy|Body Part, Organ, or Organ Component|Findings|5932,5938|false|false|false|C0042449|Veins|venous
Disorder|Disease or Syndrome|Findings|5932,5951|false|false|false|C0340766|Venous hypertension|venous hypertension
Disorder|Disease or Syndrome|Findings|5939,5951|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|Findings|5939,5951|false|false|false|||hypertension
Disorder|Disease or Syndrome|Findings|5965,5977|true|false|false|C0032326|Pneumothorax|pneumothorax
Event|Event|Findings|5965,5977|false|false|false|||pneumothorax
Finding|Finding|Hospital Course|6012,6018|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Hospital Course|6012,6018|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|Hospital Course|6019,6023|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|6019,6023|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|6019,6023|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|6019,6023|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|Hospital Course|6025,6029|false|false|false|C0004238|Atrial Fibrillation|AFib
Event|Event|Hospital Course|6025,6029|false|false|false|||AFib
Lab|Laboratory or Test Result|Hospital Course|6025,6029|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|AFib
Disorder|Disease or Syndrome|Hospital Course|6031,6034|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6031,6034|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|6031,6034|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Hospital Course|6031,6034|false|false|false|||CAD
Finding|Gene or Genome|Hospital Course|6031,6034|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|6031,6034|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|6031,6034|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6031,6034|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|Hospital Course|6036,6039|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|Hospital Course|6036,6039|false|false|false|||HTN
Event|Event|Hospital Course|6041,6044|false|false|false|||HLD
Event|Event|Hospital Course|6053,6069|false|false|false|||hospitalizations
Procedure|Health Care Activity|Hospital Course|6053,6069|false|false|false|C0019993|Hospitalization|hospitalizations
Disorder|Disease or Syndrome|Hospital Course|6085,6089|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|6085,6089|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|6085,6089|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|6085,6089|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|Hospital Course|6090,6103|false|false|false|||exacerbations
Event|Event|Hospital Course|6139,6148|false|false|false|||presented
Event|Event|Hospital Course|6154,6161|false|false|false|||dyspnea
Finding|Finding|Hospital Course|6154,6161|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|Hospital Course|6154,6161|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Event|Event|Hospital Course|6176,6184|false|false|false|||wheezing
Finding|Sign or Symptom|Hospital Course|6176,6184|false|false|false|C0043144|Wheezing|wheezing
Disorder|Neoplastic Process|Hospital Course|6185,6194|false|false|false|C0027627|Neoplasm Metastasis|secondary
Event|Event|Hospital Course|6185,6194|false|false|false|||secondary
Finding|Functional Concept|Hospital Course|6185,6194|false|false|false|C1522484|metastatic qualifier|secondary
Event|Event|Hospital Course|6199,6205|false|false|false|||severe
Finding|Finding|Hospital Course|6199,6205|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Hospital Course|6199,6205|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|Hospital Course|6206,6210|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|6206,6210|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|6206,6210|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|6206,6210|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|Hospital Course|6222,6229|false|false|false|||treated
Disorder|Disease or Syndrome|Hospital Course|6238,6242|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|6238,6242|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|6238,6242|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|6238,6242|false|false|false|C1412502|ARCN1 gene|COPD
Drug|Pharmacologic Substance|Hospital Course|6248,6258|false|false|false|C2064916|nebulizers (medication)|nebulizers
Event|Event|Hospital Course|6248,6258|false|false|false|||nebulizers
Drug|Organic Chemical|Hospital Course|6263,6271|false|false|false|C0038317|Steroids|steroids
Drug|Pharmacologic Substance|Hospital Course|6263,6271|false|false|false|C0038317|Steroids|steroids
Event|Event|Hospital Course|6263,6271|false|false|false|||steroids
Event|Event|Hospital Course|6278,6287|false|false|false|||continued
Event|Event|Hospital Course|6310,6319|false|false|false|||suffering
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6322,6325|false|false|false|C3496006|area PEa of Pandya|PEA
Disorder|Disease or Syndrome|Hospital Course|6322,6325|false|false|false|C0340861|Electromechanical dissociation|PEA
Drug|Biologically Active Substance|Hospital Course|6322,6325|false|false|false|C0030738;C0069964;C0070939;C1572795;C2702415;C3257529|PEA Preparation;Pisum sativum (pea) extract;palmidrol;pea allergenic extract;phosphoethanolamine|PEA
Drug|Food|Hospital Course|6322,6325|false|false|false|C0030738;C0069964;C0070939;C1572795;C2702415;C3257529|PEA Preparation;Pisum sativum (pea) extract;palmidrol;pea allergenic extract;phosphoethanolamine|PEA
Drug|Immunologic Factor|Hospital Course|6322,6325|false|false|false|C0030738;C0069964;C0070939;C1572795;C2702415;C3257529|PEA Preparation;Pisum sativum (pea) extract;palmidrol;pea allergenic extract;phosphoethanolamine|PEA
Drug|Organic Chemical|Hospital Course|6322,6325|false|false|false|C0030738;C0069964;C0070939;C1572795;C2702415;C3257529|PEA Preparation;Pisum sativum (pea) extract;palmidrol;pea allergenic extract;phosphoethanolamine|PEA
Drug|Pharmacologic Substance|Hospital Course|6322,6325|false|false|false|C0030738;C0069964;C0070939;C1572795;C2702415;C3257529|PEA Preparation;Pisum sativum (pea) extract;palmidrol;pea allergenic extract;phosphoethanolamine|PEA
Event|Event|Hospital Course|6322,6325|false|false|false|||PEA
Disorder|Disease or Syndrome|Hospital Course|6326,6332|false|false|false|C0018790|Cardiac Arrest|arrest
Event|Event|Hospital Course|6326,6332|false|false|false|||arrest
Event|Governmental or Regulatory Activity|Hospital Course|6326,6332|false|false|false|C0392351|Law enforcement arrest|arrest
Finding|Finding|Hospital Course|6326,6332|false|false|false|C2919124|Encounter due to problems related to other legal circumstances - arrest|arrest
Event|Event|Hospital Course|6333,6340|false|false|false|||thought
Finding|Idea or Concept|Hospital Course|6333,6340|false|false|false|C0039869;C4319827|Thought|thought
Finding|Mental Process|Hospital Course|6333,6340|false|false|false|C0039869;C4319827|Thought|thought
Event|Event|Hospital Course|6349,6358|false|false|false|||hypoxemia
Finding|Finding|Hospital Course|6349,6358|false|false|false|C0700292;C5548348|Blood oxygen concentration below reference range (finding);Hypoxemia|hypoxemia
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6369,6392|false|false|false|C0021932|Intubation, Intratracheal|endotracheal intubation
Event|Event|Hospital Course|6382,6392|false|false|false|||intubation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6382,6392|false|false|false|C0021925|Intubation (procedure)|intubation
Event|Event|Hospital Course|6398,6408|false|false|false|||mechanical
Finding|Functional Concept|Hospital Course|6398,6408|false|false|false|C0443254|mechanical method|mechanical
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6398,6408|false|false|false|C0699886|Mechanical Treatments|mechanical
Finding|Finding|Hospital Course|6398,6420|false|false|false|C4760388|Mechanical ventilation finding|mechanical ventilation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6398,6420|false|false|false|C0199470|Mechanical ventilation|mechanical ventilation
Event|Event|Hospital Course|6409,6420|false|false|false|||ventilation
Finding|Physiologic Function|Hospital Course|6409,6420|false|false|false|C0035203;C2945579|Respiration;Ventilation, function (observable entity)|ventilation
Phenomenon|Phenomenon or Process|Hospital Course|6409,6420|false|false|false|C0042491|Environmental air flow|ventilation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6409,6420|false|false|false|C0554804|Assisted breathing|ventilation
Finding|Idea or Concept|Hospital Course|6424,6433|false|false|false|C1548539;C3245481|EntityNameUseR2 - temporary;Job Status - Temporary|temporary
Finding|Intellectual Product|Hospital Course|6424,6433|false|false|false|C1548539;C3245481|EntityNameUseR2 - temporary;Job Status - Temporary|temporary
Event|Event|Hospital Course|6434,6443|false|false|false|||pacemaker
Finding|Intellectual Product|Hospital Course|6434,6443|false|false|false|C1546728||pacemaker
Event|Event|Hospital Course|6448,6454|false|false|false|||placed
Event|Event|Hospital Course|6460,6467|false|false|false|||periods
Finding|Organism Function|Hospital Course|6460,6467|false|false|false|C0025344|Menstruation|periods
Event|Event|Hospital Course|6471,6482|false|false|false|||bradycardia
Finding|Finding|Hospital Course|6471,6482|false|false|false|C0428977;C3812171|Bradycardia;Bradycardia by ECG Finding|bradycardia
Event|Event|Hospital Course|6502,6513|false|false|false|||contributed
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6521,6524|false|false|false|C3496006|area PEa of Pandya|PEA
Disorder|Disease or Syndrome|Hospital Course|6521,6524|false|false|false|C0340861|Electromechanical dissociation|PEA
Drug|Biologically Active Substance|Hospital Course|6521,6524|false|false|false|C0030738;C0069964;C0070939;C1572795;C2702415;C3257529|PEA Preparation;Pisum sativum (pea) extract;palmidrol;pea allergenic extract;phosphoethanolamine|PEA
Drug|Food|Hospital Course|6521,6524|false|false|false|C0030738;C0069964;C0070939;C1572795;C2702415;C3257529|PEA Preparation;Pisum sativum (pea) extract;palmidrol;pea allergenic extract;phosphoethanolamine|PEA
Drug|Immunologic Factor|Hospital Course|6521,6524|false|false|false|C0030738;C0069964;C0070939;C1572795;C2702415;C3257529|PEA Preparation;Pisum sativum (pea) extract;palmidrol;pea allergenic extract;phosphoethanolamine|PEA
Drug|Organic Chemical|Hospital Course|6521,6524|false|false|false|C0030738;C0069964;C0070939;C1572795;C2702415;C3257529|PEA Preparation;Pisum sativum (pea) extract;palmidrol;pea allergenic extract;phosphoethanolamine|PEA
Drug|Pharmacologic Substance|Hospital Course|6521,6524|false|false|false|C0030738;C0069964;C0070939;C1572795;C2702415;C3257529|PEA Preparation;Pisum sativum (pea) extract;palmidrol;pea allergenic extract;phosphoethanolamine|PEA
Event|Event|Hospital Course|6521,6524|false|false|false|||PEA
Disorder|Disease or Syndrome|Hospital Course|6526,6532|false|false|false|C0018790|Cardiac Arrest|arrest
Event|Event|Hospital Course|6526,6532|false|false|false|||arrest
Event|Governmental or Regulatory Activity|Hospital Course|6526,6532|false|false|false|C0392351|Law enforcement arrest|arrest
Finding|Finding|Hospital Course|6526,6532|false|false|false|C2919124|Encounter due to problems related to other legal circumstances - arrest|arrest
Event|Event|Hospital Course|6549,6562|false|false|false|||manifestation
Finding|Finding|Hospital Course|6566,6572|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Hospital Course|6566,6572|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Event|Event|Hospital Course|6573,6582|false|false|false|||hypoxemia
Finding|Finding|Hospital Course|6573,6582|false|false|false|C0700292;C5548348|Blood oxygen concentration below reference range (finding);Hypoxemia|hypoxemia
Event|Event|Hospital Course|6583,6589|false|false|false|||severe
Finding|Finding|Hospital Course|6583,6589|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Hospital Course|6583,6589|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Event|Event|Hospital Course|6591,6602|false|false|false|||hypercarbia
Finding|Finding|Hospital Course|6591,6602|false|false|false|C0020440|Hypercapnia|hypercarbia
Event|Event|Hospital Course|6603,6612|false|false|false|||preceding
Disorder|Disease or Syndrome|Hospital Course|6617,6623|false|false|false|C0018790|Cardiac Arrest|arrest
Event|Event|Hospital Course|6617,6623|false|false|false|||arrest
Event|Governmental or Regulatory Activity|Hospital Course|6617,6623|false|false|false|C0392351|Law enforcement arrest|arrest
Finding|Finding|Hospital Course|6617,6623|false|false|false|C2919124|Encounter due to problems related to other legal circumstances - arrest|arrest
Finding|Functional Concept|Hospital Course|6637,6646|false|false|false|C1516691|Cognitive|cognitive
Event|Activity|Hospital Course|6647,6655|false|false|false|C0237820||recovery
Event|Event|Hospital Course|6647,6655|false|false|false|||recovery
Finding|Organism Function|Hospital Course|6647,6655|false|false|false|C2004454|Recovery - healing process|recovery
Event|Event|Hospital Course|6665,6671|false|false|false|||unable
Finding|Finding|Hospital Course|6665,6671|false|false|false|C1299582|Unable|unable
Event|Event|Hospital Course|6691,6697|false|false|false|||weaned
Event|Event|Hospital Course|6728,6736|false|false|false|||capacity
Event|Event|Hospital Course|6745,6749|false|false|false|||able
Finding|Finding|Hospital Course|6745,6749|false|false|false|C1299581|Able (qualifier value)|able
Event|Event|Hospital Course|6753,6757|false|false|false|||make
Event|Event|Hospital Course|6761,6771|false|false|false|||understand
Event|Event|Hospital Course|6790,6794|false|false|false|||wish
Event|Event|Hospital Course|6796,6805|false|false|false|||continued
Event|Event|Hospital Course|6806,6816|false|false|false|||intubation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6806,6816|false|false|false|C0021925|Intubation (procedure)|intubation
Finding|Functional Concept|Hospital Course|6819,6829|false|false|false|C0443254|mechanical method|mechanical
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6819,6829|false|false|false|C0699886|Mechanical Treatments|mechanical
Finding|Finding|Hospital Course|6819,6841|false|false|false|C4760388|Mechanical ventilation finding|mechanical ventilation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6819,6841|false|false|false|C0199470|Mechanical ventilation|mechanical ventilation
Event|Event|Hospital Course|6830,6841|false|false|false|||ventilation
Finding|Physiologic Function|Hospital Course|6830,6841|false|false|false|C0035203;C2945579|Respiration;Ventilation, function (observable entity)|ventilation
Phenomenon|Phenomenon or Process|Hospital Course|6830,6841|false|false|false|C0042491|Environmental air flow|ventilation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6830,6841|false|false|false|C0554804|Assisted breathing|ventilation
Event|Event|Hospital Course|6844,6857|false|false|false|||re-intubation
Finding|Functional Concept|Hospital Course|6862,6872|false|false|false|C0443254|mechanical method|mechanical
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6862,6872|false|false|false|C0699886|Mechanical Treatments|mechanical
Finding|Finding|Hospital Course|6862,6884|false|false|false|C4760388|Mechanical ventilation finding|mechanical ventilation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6862,6884|false|false|false|C0199470|Mechanical ventilation|mechanical ventilation
Event|Event|Hospital Course|6873,6884|false|false|false|||ventilation
Finding|Physiologic Function|Hospital Course|6873,6884|false|false|false|C0035203;C2945579|Respiration;Ventilation, function (observable entity)|ventilation
Phenomenon|Phenomenon or Process|Hospital Course|6873,6884|false|false|false|C0042491|Environmental air flow|ventilation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6873,6884|false|false|false|C0554804|Assisted breathing|ventilation
Finding|Intellectual Product|Hospital Course|6885,6889|false|false|false|C1720092|Once - dosing instruction fragment|once
Event|Event|Hospital Course|6890,6899|false|false|false|||extubated
Disorder|Cell or Molecular Dysfunction|Hospital Course|6906,6914|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Event|Event|Hospital Course|6906,6914|false|false|false|||positive
Finding|Classification|Hospital Course|6906,6914|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|Hospital Course|6906,6914|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|Hospital Course|6928,6936|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|Hospital Course|6928,6936|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|Hospital Course|6928,6936|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|Hospital Course|6928,6936|false|false|false|C0033095||pressure
Event|Event|Hospital Course|6937,6948|false|false|false|||ventilation
Finding|Physiologic Function|Hospital Course|6937,6948|false|false|false|C0035203;C2945579|Respiration;Ventilation, function (observable entity)|ventilation
Phenomenon|Phenomenon or Process|Hospital Course|6937,6948|false|false|false|C0042491|Environmental air flow|ventilation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6937,6948|false|false|false|C0554804|Assisted breathing|ventilation
Event|Event|Hospital Course|6967,6978|false|false|false|||discussions
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6967,6978|false|false|false|C0557061|Discussion (procedure)|discussions
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6992,7002|false|false|false|C3812393|ErbB Receptors|her family
Drug|Enzyme|Hospital Course|6992,7002|false|false|false|C3812393|ErbB Receptors|her family
Finding|Receptor|Hospital Course|6992,7002|false|false|false|C3812393|ErbB Receptors|her family
Event|Event|Hospital Course|6996,7002|false|false|false|||family
Finding|Classification|Hospital Course|6996,7002|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Hospital Course|6996,7002|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Hospital Course|6996,7002|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Hospital Course|6996,7002|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Event|Event|Hospital Course|7012,7024|false|false|false|||transitioned
Attribute|Clinical Attribute|Hospital Course|7029,7032|false|false|false|C4285234||DNR
Drug|Antibiotic|Hospital Course|7029,7032|false|false|false|C0011015|daunorubicin|DNR
Drug|Organic Chemical|Hospital Course|7029,7032|false|false|false|C0011015|daunorubicin|DNR
Event|Event|Hospital Course|7029,7032|false|false|false|||DNR
Finding|Finding|Hospital Course|7029,7032|false|false|false|C0079252;C0582114|Do not resuscitate status;Do-Not-Resuscitate Orders|DNR
Finding|Intellectual Product|Hospital Course|7029,7032|false|false|false|C0079252;C0582114|Do not resuscitate status;Do-Not-Resuscitate Orders|DNR
Drug|Organic Chemical|Hospital Course|7041,7048|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Drug|Pharmacologic Substance|Hospital Course|7041,7048|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Event|Event|Hospital Course|7041,7048|false|false|false|||comfort
Finding|Mental Process|Hospital Course|7041,7048|false|false|false|C1331418|Comfort|comfort
Finding|Finding|Hospital Course|7049,7057|false|false|false|C1961028|Oriented to place|oriented
Event|Activity|Hospital Course|7058,7062|false|false|false|C1947933|care activity|care
Event|Event|Hospital Course|7058,7062|false|false|false|||care
Finding|Finding|Hospital Course|7058,7062|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Hospital Course|7058,7062|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Event|Event|Hospital Course|7072,7081|false|false|false|||extubated
Finding|Finding|Hospital Course|7100,7104|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Hospital Course|7100,7104|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Hospital Course|7100,7104|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7110,7120|false|false|false|C3812393|ErbB Receptors|her family
Drug|Enzyme|Hospital Course|7110,7120|false|false|false|C3812393|ErbB Receptors|her family
Finding|Receptor|Hospital Course|7110,7120|false|false|false|C3812393|ErbB Receptors|her family
Event|Event|Hospital Course|7114,7120|false|false|false|||family
Finding|Classification|Hospital Course|7114,7120|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Hospital Course|7114,7120|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Hospital Course|7114,7120|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Hospital Course|7114,7120|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Event|Event|Hospital Course|7128,7135|false|false|false|||passing
Attribute|Clinical Attribute|Hospital Course|7141,7152|false|false|false|C0231832|Respiratory rate|respiratory
Event|Event|Hospital Course|7141,7152|false|false|false|||respiratory
Finding|Body Substance|Hospital Course|7141,7152|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|Hospital Course|7141,7152|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|Hospital Course|7141,7152|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Event|Event|Hospital Course|7154,7161|false|false|false|||failure
Finding|Functional Concept|Hospital Course|7154,7161|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|Hospital Course|7154,7161|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|Hospital Course|7154,7161|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|Hospital Course|7193,7200|false|false|false|||Autopsy
Finding|Intellectual Product|Hospital Course|7193,7200|false|false|false|C1546546||Autopsy
Procedure|Diagnostic Procedure|Hospital Course|7193,7200|false|false|false|C0004398;C1548821|Autopsy;Autopsy - Consent type|Autopsy
Procedure|Health Care Activity|Hospital Course|7193,7200|false|false|false|C0004398;C1548821|Autopsy;Autopsy - Consent type|Autopsy
Event|Event|Hospital Course|7205,7213|false|false|false|||declined
Finding|Classification|Hospital Course|7218,7224|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Hospital Course|7218,7224|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Hospital Course|7218,7224|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Hospital Course|7218,7224|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Event|Event|Hospital Course|7248,7253|false|false|false|||found
Drug|Organic Chemical|Hospital Course|7264,7267|false|false|false|C0939812|Ruta graveolens preparation|RUE
Drug|Pharmacologic Substance|Hospital Course|7264,7267|false|false|false|C0939812|Ruta graveolens preparation|RUE
Anatomy|Body Location or Region|Hospital Course|7268,7271|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Hospital Course|7268,7271|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Hospital Course|7268,7271|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|Hospital Course|7268,7271|false|false|false|||DVT
Event|Event|Hospital Course|7281,7288|false|false|false|||treated
Drug|Biologically Active Substance|Hospital Course|7295,7302|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|Hospital Course|7295,7302|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|Hospital Course|7295,7302|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Disorder|Neoplastic Process|Hospital Course|7303,7306|false|false|false|C1135868|Gestational Trophoblastic Neoplasms|gtt
Drug|Biomedical or Dental Material|Hospital Course|7303,7306|false|false|false|C0991568|Drops - Drug Form|gtt
Event|Event|Hospital Course|7303,7306|false|false|false|||gtt
Procedure|Laboratory Procedure|Hospital Course|7303,7306|false|false|false|C0017741|Glucose tolerance test|gtt
Event|Event|Hospital Course|7323,7327|false|false|false|||used
Event|Event|Hospital Course|7332,7347|false|false|false|||anticoagulation
Finding|Finding|Hospital Course|7332,7347|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|Hospital Course|7332,7347|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7332,7347|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7357,7363|false|false|false|C0018792|Heart Atrium|atrial
Attribute|Clinical Attribute|Hospital Course|7357,7376|false|false|false|C2926591||atrial fibrillation
Disorder|Disease or Syndrome|Hospital Course|7357,7376|false|false|false|C0004238|Atrial Fibrillation|atrial fibrillation
Lab|Laboratory or Test Result|Hospital Course|7357,7376|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|atrial fibrillation
Disorder|Disease or Syndrome|Hospital Course|7364,7376|false|false|false|C0232197|Fibrillation|fibrillation
Event|Event|Hospital Course|7364,7376|false|false|false|||fibrillation
Event|Event|Hospital Course|7398,7410|false|false|false|||transitioned
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7415,7425|false|false|false|C0048470|argatroban|argatroban
Drug|Pharmacologic Substance|Hospital Course|7415,7425|false|false|false|C0048470|argatroban|argatroban
Event|Event|Hospital Course|7415,7425|false|false|false|||argatroban
Event|Event|Hospital Course|7430,7437|false|false|false|||concern
Finding|Idea or Concept|Hospital Course|7430,7437|false|false|false|C2699424|Concern|concern
Disorder|Disease or Syndrome|Hospital Course|7441,7444|false|false|false|C0272285|Heparin-induced thrombocytopenia|HIT
Event|Event|Hospital Course|7441,7444|false|false|false|||HIT
Finding|Functional Concept|Hospital Course|7441,7444|false|false|false|C1708373|Hit - database search return|HIT
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7450,7453|false|false|false|C0032183;C3887656|Platelet Factor 4;Platelet Factor 4, human|PF4
Drug|Immunologic Factor|Hospital Course|7450,7453|false|false|false|C0032183;C3887656|Platelet Factor 4;Platelet Factor 4, human|PF4
Finding|Gene or Genome|Hospital Course|7450,7453|false|false|false|C1335206|PF4 gene|PF4
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7454,7464|false|false|false|C0003241;C3495458|Antibodies;antibodies (medication)|antibodies
Drug|Immunologic Factor|Hospital Course|7454,7464|false|false|false|C0003241;C3495458|Antibodies;antibodies (medication)|antibodies
Drug|Pharmacologic Substance|Hospital Course|7454,7464|false|false|false|C0003241;C3495458|Antibodies;antibodies (medication)|antibodies
Event|Event|Hospital Course|7454,7464|false|false|false|||antibodies
Event|Event|Hospital Course|7465,7473|false|false|false|||returned
Finding|Finding|Hospital Course|7478,7486|false|false|false|C0442811;C5202917|IPSS-R Risk Category Very Low;Very low (qualifier value)|very low
Finding|Finding|Hospital Course|7483,7486|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Hospital Course|7483,7486|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Attribute|Clinical Attribute|Hospital Course|7503,7512|false|false|false|C0945731||diagnosis
Event|Event|Hospital Course|7503,7512|false|false|false|||diagnosis
Finding|Classification|Hospital Course|7503,7512|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|Hospital Course|7503,7512|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|Hospital Course|7503,7512|false|false|false|C0011900|Diagnosis|diagnosis
Event|Event|Hospital Course|7513,7521|false|false|false|||unlikely
Finding|Finding|Hospital Course|7513,7521|false|false|false|C0750558|Unlikely|unlikely
Event|Event|Hospital Course|7538,7545|false|false|false|||treated
Finding|Intellectual Product|Hospital Course|7553,7558|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Disease or Syndrome|Hospital Course|7553,7568|false|false|false|C0149512|Acute sinusitis|acute sinusitis
Disorder|Disease or Syndrome|Hospital Course|7559,7568|false|false|false|C0037199|Sinusitis|sinusitis
Event|Event|Hospital Course|7559,7568|false|false|false|||sinusitis
Drug|Antibiotic|Hospital Course|7574,7583|false|false|false|C0591132|Augmentin|Augmentin
Drug|Organic Chemical|Hospital Course|7574,7583|false|false|false|C0591132|Augmentin|Augmentin
Event|Event|Hospital Course|7574,7583|false|false|false|||Augmentin
Finding|Idea or Concept|Hospital Course|7596,7604|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|Hospital Course|7605,7609|false|false|false|||stay
Attribute|Clinical Attribute|Hospital Course|7614,7625|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|7614,7625|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|7614,7625|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|7614,7625|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|7614,7638|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|7629,7638|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|7629,7638|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|Hospital Course|7657,7667|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Hospital Course|7657,7667|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|Hospital Course|7657,7672|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|Hospital Course|7668,7672|false|false|false|||list
Finding|Intellectual Product|Hospital Course|7668,7672|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|Hospital Course|7676,7684|false|false|false|||accurate
Drug|Organic Chemical|Hospital Course|7689,7697|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Hospital Course|7689,7697|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Hospital Course|7689,7697|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|Hospital Course|7689,7697|false|false|false|||complete
Finding|Functional Concept|Hospital Course|7689,7697|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|7689,7697|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|Hospital Course|7702,7715|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|7702,7715|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Hospital Course|7702,7715|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|7702,7715|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|Hospital Course|7730,7733|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|7734,7738|false|false|false|C2598155||Pain
Event|Event|Hospital Course|7734,7738|false|false|false|||Pain
Finding|Functional Concept|Hospital Course|7734,7738|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Hospital Course|7734,7738|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Drug|Organic Chemical|Hospital Course|7743,7753|false|false|false|C3464797|Calcitrate|Calcitrate
Drug|Pharmacologic Substance|Hospital Course|7743,7753|false|false|false|C3464797|Calcitrate|Calcitrate
Drug|Organic Chemical|Hospital Course|7754,7761|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|7754,7761|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|7754,7761|false|false|false|C0042890|Vitamins|Vitamin
Event|Event|Hospital Course|7754,7761|false|false|false|||Vitamin
Drug|Hormone|Hospital Course|7754,7763|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|Hospital Course|7754,7763|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|Hospital Course|7754,7763|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|Hospital Course|7754,7763|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|Hospital Course|7754,7763|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|Hospital Course|7762,7763|false|false|false|||D
Drug|Biologically Active Substance|Hospital Course|7765,7772|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Element, Ion, or Isotope|Hospital Course|7765,7772|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Inorganic Chemical|Hospital Course|7765,7772|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Pharmacologic Substance|Hospital Course|7765,7772|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Vitamin|Hospital Course|7765,7772|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Event|Event|Hospital Course|7765,7772|false|false|false|||calcium
Finding|Physiologic Function|Hospital Course|7765,7772|false|false|false|C4553026|Calcium metabolic function|calcium
Procedure|Laboratory Procedure|Hospital Course|7765,7772|false|false|false|C0201925|Calcium measurement|calcium
Drug|Organic Chemical|Hospital Course|7765,7780|false|false|false|C0108101|calcium citrate|calcium citrate
Drug|Pharmacologic Substance|Hospital Course|7765,7780|false|false|false|C0108101|calcium citrate|calcium citrate
Drug|Organic Chemical|Hospital Course|7773,7780|false|false|false|C0008857;C0376259|Citrates;citrate|citrate
Drug|Pharmacologic Substance|Hospital Course|7773,7780|false|false|false|C0008857;C0376259|Citrates;citrate|citrate
Event|Event|Hospital Course|7773,7780|false|false|false|||citrate
Procedure|Laboratory Procedure|Hospital Course|7773,7780|false|false|false|C0201956|Citrate measurement|citrate
Drug|Organic Chemical|Hospital Course|7781,7788|false|false|false|C0042890|Vitamins|vitamin
Drug|Pharmacologic Substance|Hospital Course|7781,7788|false|false|false|C0042890|Vitamins|vitamin
Drug|Vitamin|Hospital Course|7781,7788|false|false|false|C0042890|Vitamins|vitamin
Event|Event|Hospital Course|7781,7788|false|false|false|||vitamin
Drug|Organic Chemical|Hospital Course|7781,7791|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Pharmacologic Substance|Hospital Course|7781,7791|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Vitamin|Hospital Course|7781,7791|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Anatomy|Body Space or Junction|Hospital Course|7814,7818|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|7814,7818|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|7814,7818|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|7814,7818|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|Hospital Course|7819,7824|false|false|false|||DAILY
Drug|Organic Chemical|Hospital Course|7829,7839|false|false|false|C0213771|tiotropium|Tiotropium
Drug|Pharmacologic Substance|Hospital Course|7829,7839|false|false|false|C0213771|tiotropium|Tiotropium
Event|Event|Hospital Course|7829,7839|false|false|false|||Tiotropium
Drug|Organic Chemical|Hospital Course|7829,7847|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Pharmacologic Substance|Hospital Course|7829,7847|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Inorganic Chemical|Hospital Course|7840,7847|false|false|false|C0006222|Bromides|Bromide
Event|Event|Hospital Course|7840,7847|false|false|false|||Bromide
Procedure|Laboratory Procedure|Hospital Course|7840,7847|false|false|false|C0202341|Bromides measurement|Bromide
Disorder|Congenital Abnormality|Hospital Course|7850,7853|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|CAP
Drug|Biomedical or Dental Material|Hospital Course|7850,7853|false|false|false|C0006935|capsule (pharmacologic)|CAP
Event|Event|Hospital Course|7850,7853|false|false|false|||CAP
Finding|Gene or Genome|Hospital Course|7850,7853|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|CAP
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7850,7853|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|CAP
Drug|Organic Chemical|Hospital Course|7867,7879|false|false|false|C0039771|theophylline|Theophylline
Drug|Pharmacologic Substance|Hospital Course|7867,7879|false|false|false|C0039771|theophylline|Theophylline
Event|Event|Hospital Course|7867,7879|false|false|false|||Theophylline
Procedure|Laboratory Procedure|Hospital Course|7867,7879|false|false|false|C0039773|Assay of theophylline|Theophylline
Drug|Organic Chemical|Hospital Course|7867,7882|false|false|false|C0939729|Theophylline SR|Theophylline SR
Drug|Pharmacologic Substance|Hospital Course|7867,7882|false|false|false|C0939729|Theophylline SR|Theophylline SR
Disorder|Mental or Behavioral Dysfunction|Hospital Course|7893,7896|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7893,7896|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|7893,7896|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|7893,7896|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|7893,7896|false|false|false|C1332410|BID gene|BID
Drug|Antibiotic|Hospital Course|7911,7923|false|false|false|C0041041|trimethoprim|Trimethoprim
Drug|Organic Chemical|Hospital Course|7911,7923|false|false|false|C0041041|trimethoprim|Trimethoprim
Drug|Biomedical or Dental Material|Hospital Course|7929,7932|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|Hospital Course|7929,7932|false|false|false|||TAB
Event|Event|Hospital Course|7942,7953|false|false|false|||prophylaxis
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7942,7953|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Finding|Idea or Concept|Hospital Course|7964,7968|false|false|false|C0233324;C1705313|Term (lexical);Term Birth|term
Finding|Organism Function|Hospital Course|7964,7968|false|false|false|C0233324;C1705313|Term (lexical);Term Birth|term
Drug|Organic Chemical|Hospital Course|7969,7976|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Drug|Pharmacologic Substance|Hospital Course|7969,7976|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Finding|Individual Behavior|Hospital Course|7969,7980|false|false|false|C0281991|Use of steroids|steroid use
Event|Event|Hospital Course|7977,7980|false|false|false|||use
Finding|Functional Concept|Hospital Course|7977,7980|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|Hospital Course|7977,7980|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Drug|Organic Chemical|Hospital Course|7985,7995|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Pharmacologic Substance|Hospital Course|7985,7995|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Hormone|Hospital Course|8016,8026|false|false|false|C0032952|prednisone|PredniSONE
Drug|Organic Chemical|Hospital Course|8016,8026|false|false|false|C0032952|prednisone|PredniSONE
Drug|Pharmacologic Substance|Hospital Course|8016,8026|false|false|false|C0032952|prednisone|PredniSONE
Drug|Organic Chemical|Hospital Course|8046,8055|false|false|false|C0024002|lorazepam|Lorazepam
Drug|Pharmacologic Substance|Hospital Course|8046,8055|false|false|false|C0024002|lorazepam|Lorazepam
Finding|Gene or Genome|Hospital Course|8070,8073|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Pharmacologic Substance|Hospital Course|8074,8082|false|false|false|C1950154|Insomnia homeopathic medication|Insomnia
Event|Event|Hospital Course|8074,8082|false|false|false|||Insomnia
Finding|Sign or Symptom|Hospital Course|8074,8082|false|false|false|C0917801|Sleeplessness|Insomnia
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8084,8091|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|Hospital Course|8084,8091|false|false|false|||anxiety
Finding|Sign or Symptom|Hospital Course|8084,8091|false|false|false|C0860603|Anxiety symptoms|anxiety
Disorder|Disease or Syndrome|Hospital Course|8093,8100|false|false|false|C1135208|Vertigo as late effect of cerebrovascular disease|vertigo
Event|Event|Hospital Course|8093,8100|false|false|false|||vertigo
Finding|Sign or Symptom|Hospital Course|8093,8100|false|false|false|C0042571|Vertigo|vertigo
Drug|Organic Chemical|Hospital Course|8105,8116|false|false|false|C0090306|latanoprost|Latanoprost
Drug|Pharmacologic Substance|Hospital Course|8105,8116|false|false|false|C0090306|latanoprost|Latanoprost
Finding|Functional Concept|Hospital Course|8124,8129|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|Hospital Course|8139,8143|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|Hospital Course|8139,8143|false|false|false|C1705648|Dropping|DROP
Event|Event|Hospital Course|8139,8143|false|false|false|||DROP
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8144,8153|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8149,8153|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|Hospital Course|8149,8153|false|false|false|C5848506||EYES
Drug|Organic Chemical|Hospital Course|8163,8173|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|Hospital Course|8163,8173|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|Hospital Course|8163,8185|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|Hospital Course|8163,8185|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Event|Event|Hospital Course|8174,8185|false|false|false|||Mononitrate
Finding|Finding|Hospital Course|8187,8195|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|8187,8195|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Hospital Course|8196,8203|false|false|false|||Release
Finding|Functional Concept|Hospital Course|8196,8203|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|8196,8203|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8196,8203|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Hospital Course|8226,8237|false|false|false|C0027235|ipratropium|Ipratropium
Drug|Pharmacologic Substance|Hospital Course|8226,8237|false|false|false|C0027235|ipratropium|Ipratropium
Event|Event|Hospital Course|8226,8237|false|false|false|||Ipratropium
Drug|Organic Chemical|Hospital Course|8226,8245|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Pharmacologic Substance|Hospital Course|8226,8245|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Inorganic Chemical|Hospital Course|8238,8245|false|false|false|C0006222|Bromides|Bromide
Event|Event|Hospital Course|8238,8245|false|false|false|||Bromide
Procedure|Laboratory Procedure|Hospital Course|8238,8245|false|false|false|C0202341|Bromides measurement|Bromide
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8246,8249|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|Hospital Course|8246,8249|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|Hospital Course|8246,8249|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Event|Event|Hospital Course|8246,8249|false|false|false|||Neb
Finding|Cell Function|Hospital Course|8246,8249|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|Hospital Course|8246,8249|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8252,8255|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|Hospital Course|8252,8255|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|Hospital Course|8252,8255|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|Hospital Course|8252,8255|false|false|false|||NEB
Finding|Cell Function|Hospital Course|8252,8255|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|8252,8255|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Event|Event|Hospital Course|8263,8271|false|false|false|||Wheezing
Finding|Sign or Symptom|Hospital Course|8263,8271|false|false|false|C0043144|Wheezing|Wheezing
Drug|Organic Chemical|Hospital Course|8277,8296|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Pharmacologic Substance|Hospital Course|8277,8296|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Organic Chemical|Hospital Course|8317,8328|false|false|false|C0018305|guaifenesin|Guaifenesin
Drug|Pharmacologic Substance|Hospital Course|8317,8328|false|false|false|C0018305|guaifenesin|Guaifenesin
Finding|Gene or Genome|Hospital Course|8343,8346|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|Hospital Course|8347,8352|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|Hospital Course|8347,8352|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|Hospital Course|8347,8352|false|false|false|||cough
Finding|Sign or Symptom|Hospital Course|8347,8352|false|false|false|C0010200|Coughing|cough
Drug|Organic Chemical|Hospital Course|8358,8369|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|8358,8369|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|8358,8380|false|false|false|C0939232|fluticasone / salmeterol|Fluticasone-Salmeterol
Drug|Organic Chemical|Hospital Course|8358,8387|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Pharmacologic Substance|Hospital Course|8358,8387|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Organic Chemical|Hospital Course|8370,8380|false|false|false|C0073992|salmeterol|Salmeterol
Drug|Pharmacologic Substance|Hospital Course|8370,8380|false|false|false|C0073992|salmeterol|Salmeterol
Event|Event|Hospital Course|8381,8387|false|false|false|||Diskus
Drug|Biomedical or Dental Material|Hospital Course|8400,8403|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Organic Chemical|Hospital Course|8400,8403|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Pharmacologic Substance|Hospital Course|8400,8403|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Event|Event|Hospital Course|8400,8403|false|false|false|||INH
Finding|Functional Concept|Hospital Course|8400,8403|false|false|false|C0205535|Inhalation Route of Administration|INH
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8407,8410|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8407,8410|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8407,8410|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|8407,8410|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|8407,8410|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|8416,8427|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|8416,8427|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|Hospital Course|8416,8427|false|false|false|||Fluticasone
Drug|Organic Chemical|Hospital Course|8416,8438|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|Hospital Course|8416,8438|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|Hospital Course|8428,8438|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8439,8444|false|false|false|C0028429||NASAL
Drug|Biomedical or Dental Material|Hospital Course|8439,8444|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Organic Chemical|Hospital Course|8439,8444|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Pharmacologic Substance|Hospital Course|8439,8444|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Finding|Finding|Hospital Course|8439,8444|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Finding|Functional Concept|Hospital Course|8439,8444|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Event|Event|Hospital Course|8447,8451|false|false|false|||SPRY
Event|Event|Hospital Course|8455,8460|false|false|false|||DAILY
Finding|Gene or Genome|Hospital Course|8461,8464|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|8465,8474|false|false|false|C1717415||allergies
Event|Event|Hospital Course|8465,8474|false|false|false|||allergies
Finding|Pathologic Function|Hospital Course|8465,8474|false|false|false|C0020517|Hypersensitivity|allergies
Drug|Element, Ion, or Isotope|Hospital Course|8480,8487|false|false|false|C2346592|Ferrous|Ferrous
Drug|Inorganic Chemical|Hospital Course|8480,8495|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Pharmacologic Substance|Hospital Course|8480,8495|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Element, Ion, or Isotope|Hospital Course|8488,8495|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Inorganic Chemical|Hospital Course|8488,8495|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Pharmacologic Substance|Hospital Course|8488,8495|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Organic Chemical|Hospital Course|8517,8528|false|false|false|C0165590|dorzolamide|Dorzolamide
Drug|Pharmacologic Substance|Hospital Course|8517,8528|false|false|false|C0165590|dorzolamide|Dorzolamide
Event|Event|Hospital Course|8532,8537|false|false|false|||Ophth
Finding|Functional Concept|Hospital Course|8532,8537|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|Hospital Course|8547,8551|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|Hospital Course|8547,8551|false|false|false|C1705648|Dropping|DROP
Event|Event|Hospital Course|8547,8551|false|false|false|||DROP
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8552,8561|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8557,8561|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|Hospital Course|8557,8561|false|false|false|C5848506||EYES
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8562,8565|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8562,8565|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8562,8565|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|8562,8565|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|8562,8565|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|8571,8580|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|Hospital Course|8571,8580|false|false|false|C0001927|albuterol|albuterol
Event|Event|Hospital Course|8571,8580|false|false|false|||albuterol
Drug|Organic Chemical|Hospital Course|8571,8588|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|Hospital Course|8571,8588|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|Hospital Course|8581,8588|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|Hospital Course|8581,8588|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|Hospital Course|8581,8588|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Event|Event|Hospital Course|8581,8588|false|false|false|||sulfate
Finding|Functional Concept|Hospital Course|8606,8616|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Organism Function|Hospital Course|8606,8616|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Event|Event|Hospital Course|8617,8620|false|false|false|||Q4H
Drug|Organic Chemical|Hospital Course|8626,8634|false|false|false|C1831808|apixaban|Apixaban
Drug|Pharmacologic Substance|Hospital Course|8626,8634|false|false|false|C1831808|apixaban|Apixaban
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8643,8646|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8643,8646|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8643,8646|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|8643,8646|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|8643,8646|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|8652,8659|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Hospital Course|8652,8659|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|Hospital Course|8680,8692|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|8680,8692|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|Hospital Course|8711,8720|false|false|false|C0012373|diltiazem|Diltiazem
Drug|Pharmacologic Substance|Hospital Course|8711,8720|false|false|false|C0012373|diltiazem|Diltiazem
Finding|Finding|Hospital Course|8721,8729|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|8721,8729|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Hospital Course|8730,8737|false|false|false|||Release
Finding|Functional Concept|Hospital Course|8730,8737|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|8730,8737|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8730,8737|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8748,8751|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8748,8751|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8748,8751|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|8748,8751|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|8748,8751|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|8757,8765|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|8757,8765|false|false|false|C1692318|docusate|Docusate
Drug|Organic Chemical|Hospital Course|8757,8772|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|Hospital Course|8757,8772|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|Hospital Course|8766,8772|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|8766,8772|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|8766,8772|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|8766,8772|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|8766,8772|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|8766,8772|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8783,8786|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8783,8786|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8783,8786|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|8783,8786|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|8783,8786|false|false|false|C1332410|BID gene|BID
Drug|Biologically Active Substance|Hospital Course|8792,8798|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|8792,8798|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|8792,8798|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|8792,8798|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|8792,8798|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|8792,8798|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Inorganic Chemical|Hospital Course|8792,8807|false|false|false|C0037494|sodium chloride|Sodium Chloride
Drug|Clinical Drug|Hospital Course|8792,8813|false|false|false|C3213708|Sodium Chloride Nasal Product|Sodium Chloride Nasal
Drug|Element, Ion, or Isotope|Hospital Course|8799,8807|false|false|false|C0008203;C0596019|Chlorides;chloride ion|Chloride
Event|Event|Hospital Course|8799,8807|false|false|false|||Chloride
Finding|Physiologic Function|Hospital Course|8799,8807|false|false|false|C4553021|Chloride metabolic function|Chloride
Procedure|Laboratory Procedure|Hospital Course|8799,8807|false|false|false|C0201952|Chloride measurement|Chloride
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8808,8813|false|false|false|C0028429||Nasal
Drug|Biomedical or Dental Material|Hospital Course|8808,8813|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Organic Chemical|Hospital Course|8808,8813|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Pharmacologic Substance|Hospital Course|8808,8813|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Finding|Finding|Hospital Course|8808,8813|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Functional Concept|Hospital Course|8808,8813|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Event|Event|Hospital Course|8818,8822|false|false|false|||SPRY
Finding|Gene or Genome|Hospital Course|8830,8833|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8834,8839|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|Hospital Course|8834,8839|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|Hospital Course|8834,8839|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|Hospital Course|8834,8839|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|Hospital Course|8834,8839|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|Hospital Course|8834,8839|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Sign or Symptom|Hospital Course|8834,8850|false|false|false|C0858259|Nasal discomfort|nasal discomfort
Event|Event|Hospital Course|8840,8850|false|false|false|||discomfort
Finding|Sign or Symptom|Hospital Course|8840,8850|false|false|false|C2364135|Discomfort|discomfort
Drug|Organic Chemical|Hospital Course|8856,8864|false|false|false|C0026549|morphine|Morphine
Drug|Pharmacologic Substance|Hospital Course|8856,8864|false|false|false|C0026549|morphine|Morphine
Drug|Organic Chemical|Hospital Course|8856,8872|false|false|false|C0066814|morphine sulfate|Morphine Sulfate
Drug|Pharmacologic Substance|Hospital Course|8856,8872|false|false|false|C0066814|morphine sulfate|Morphine Sulfate
Drug|Element, Ion, or Isotope|Hospital Course|8865,8872|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Inorganic Chemical|Hospital Course|8865,8872|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Pharmacologic Substance|Hospital Course|8865,8872|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Event|Event|Hospital Course|8865,8872|false|false|false|||Sulfate
Anatomy|Body Space or Junction|Hospital Course|8874,8878|false|false|false|C0226896|Oral cavity|Oral
Drug|Biomedical or Dental Material|Hospital Course|8874,8878|false|false|false|C1272919|Oral Dosage Form|Oral
Finding|Finding|Hospital Course|8874,8878|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Finding|Functional Concept|Hospital Course|8874,8878|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Drug|Biomedical or Dental Material|Hospital Course|8874,8887|false|false|false|C0991536|Oral Solution|Oral Solution
Drug|Biomedical or Dental Material|Hospital Course|8879,8887|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|Solution
Drug|Substance|Hospital Course|8879,8887|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|Solution
Event|Event|Hospital Course|8879,8887|false|false|false|||Solution
Finding|Conceptual Entity|Hospital Course|8879,8887|false|false|false|C2699488|Resolution|Solution
Finding|Gene or Genome|Hospital Course|8909,8912|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|8914,8923|false|false|false|||shortness
Attribute|Clinical Attribute|Hospital Course|8914,8933|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|Hospital Course|8914,8933|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|Hospital Course|8927,8933|false|false|false|C0225386|Breath|breath
Drug|Organic Chemical|Hospital Course|8939,8949|false|false|false|C0054201|budesonide|Budesonide
Drug|Pharmacologic Substance|Hospital Course|8939,8949|false|false|false|C0054201|budesonide|Budesonide
Drug|Clinical Drug|Hospital Course|8939,8955|false|false|false|C0360546;C3832695|Budesonide Nasal (Brand Name);Budesonide Nasal Product|Budesonide Nasal
Drug|Pharmacologic Substance|Hospital Course|8939,8955|false|false|false|C0360546;C3832695|Budesonide Nasal (Brand Name);Budesonide Nasal Product|Budesonide Nasal
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8950,8955|false|false|false|C0028429||Nasal
Drug|Biomedical or Dental Material|Hospital Course|8950,8955|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Organic Chemical|Hospital Course|8950,8955|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Pharmacologic Substance|Hospital Course|8950,8955|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Finding|Finding|Hospital Course|8950,8955|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Functional Concept|Hospital Course|8950,8955|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Event|Event|Hospital Course|8956,8963|false|false|false|||Inhaler
Finding|Functional Concept|Hospital Course|8956,8963|false|false|false|C4319647|Inhaler (unit of presentation)|Inhaler
Event|Event|Hospital Course|8988,8997|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|8988,8997|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|8988,8997|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|8988,8997|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|8988,8997|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|8988,9009|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|8998,9009|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|8998,9009|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|8998,9009|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|8998,9009|false|false|false|C4284232|Medications|Medications
Event|Event|Hospital Course|9019,9028|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|9019,9028|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|9019,9028|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|9019,9028|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|9019,9028|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|9019,9040|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|9019,9040|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|9029,9040|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|9029,9040|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|9029,9040|false|false|false|C0184758|Patient disposition|Disposition
Finding|Idea or Concept|Hospital Course|9042,9049|false|false|false|C0011065;C0231800;C1548436;C1549070;C1704631|Certificate Status - Expired;Cessation of life;Expiration;Expiration, Respiratory;Referral status - Expired|Expired
Finding|Organism Function|Hospital Course|9042,9049|false|false|false|C0011065;C0231800;C1548436;C1549070;C1704631|Certificate Status - Expired;Cessation of life;Expiration;Expiration, Respiratory;Referral status - Expired|Expired
Event|Event|Hospital Course|9052,9061|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|9052,9061|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|9052,9061|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|9052,9061|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|9052,9061|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|9052,9071|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|9062,9071|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|9062,9071|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|9062,9071|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|9062,9071|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|9062,9071|false|false|false|C0011900|Diagnosis|Diagnosis
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|9096,9099|false|false|false|C3496006|area PEa of Pandya|PEA
Disorder|Disease or Syndrome|Principle Diagnosis|9096,9099|false|false|false|C0340861|Electromechanical dissociation|PEA
Drug|Biologically Active Substance|Principle Diagnosis|9096,9099|false|false|false|C0030738;C0069964;C0070939;C1572795;C2702415;C3257529|PEA Preparation;Pisum sativum (pea) extract;palmidrol;pea allergenic extract;phosphoethanolamine|PEA
Drug|Food|Principle Diagnosis|9096,9099|false|false|false|C0030738;C0069964;C0070939;C1572795;C2702415;C3257529|PEA Preparation;Pisum sativum (pea) extract;palmidrol;pea allergenic extract;phosphoethanolamine|PEA
Drug|Immunologic Factor|Principle Diagnosis|9096,9099|false|false|false|C0030738;C0069964;C0070939;C1572795;C2702415;C3257529|PEA Preparation;Pisum sativum (pea) extract;palmidrol;pea allergenic extract;phosphoethanolamine|PEA
Drug|Organic Chemical|Principle Diagnosis|9096,9099|false|false|false|C0030738;C0069964;C0070939;C1572795;C2702415;C3257529|PEA Preparation;Pisum sativum (pea) extract;palmidrol;pea allergenic extract;phosphoethanolamine|PEA
Drug|Pharmacologic Substance|Principle Diagnosis|9096,9099|false|false|false|C0030738;C0069964;C0070939;C1572795;C2702415;C3257529|PEA Preparation;Pisum sativum (pea) extract;palmidrol;pea allergenic extract;phosphoethanolamine|PEA
Disorder|Disease or Syndrome|Principle Diagnosis|9100,9106|false|false|false|C0018790|Cardiac Arrest|Arrest
Event|Event|Principle Diagnosis|9100,9106|false|false|false|||Arrest
Event|Governmental or Regulatory Activity|Principle Diagnosis|9100,9106|false|false|false|C0392351|Law enforcement arrest|Arrest
Finding|Finding|Principle Diagnosis|9100,9106|false|false|false|C2919124|Encounter due to problems related to other legal circumstances - arrest|Arrest
Attribute|Clinical Attribute|Principle Diagnosis|9108,9119|false|false|false|C0231832|Respiratory rate|Respiratory
Finding|Body Substance|Principle Diagnosis|9108,9119|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|Respiratory
Finding|Functional Concept|Principle Diagnosis|9108,9119|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|Respiratory
Finding|Intellectual Product|Principle Diagnosis|9108,9119|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|Respiratory
Disorder|Disease or Syndrome|Principle Diagnosis|9108,9127|false|false|false|C1145670|Respiratory Failure|Respiratory Failure
Event|Event|Principle Diagnosis|9120,9127|false|false|false|||Failure
Finding|Functional Concept|Principle Diagnosis|9120,9127|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|Failure
Finding|Idea or Concept|Principle Diagnosis|9120,9127|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|Failure
Finding|Individual Behavior|Principle Diagnosis|9120,9127|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|Failure
Disorder|Disease or Syndrome|Principle Diagnosis|9128,9132|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Principle Diagnosis|9128,9132|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Principle Diagnosis|9128,9132|false|false|false|||COPD
Finding|Gene or Genome|Principle Diagnosis|9128,9132|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|Principle Diagnosis|9133,9142|false|false|false|C0037199|Sinusitis|Sinusitis
Event|Event|Principle Diagnosis|9133,9142|false|false|false|||Sinusitis
Drug|Organic Chemical|Principle Diagnosis|9143,9146|false|false|false|C0939812|Ruta graveolens preparation|RUE
Drug|Pharmacologic Substance|Principle Diagnosis|9143,9146|false|false|false|C0939812|Ruta graveolens preparation|RUE
Anatomy|Body Location or Region|Principle Diagnosis|9147,9150|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Principle Diagnosis|9147,9150|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Principle Diagnosis|9147,9150|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|Principle Diagnosis|9147,9150|false|false|false|||DVT
Disorder|Neoplastic Process|Principle Diagnosis|9152,9161|false|false|false|C0027627|Neoplasm Metastasis|SECONDARY
Finding|Functional Concept|Principle Diagnosis|9152,9161|false|false|false|C1522484|metastatic qualifier|SECONDARY
Event|Event|Principle Diagnosis|9162,9171|false|false|false|||DIAGNOSES
Procedure|Diagnostic Procedure|Principle Diagnosis|9162,9171|false|false|false|C0011900|Diagnosis|DIAGNOSES
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|9173,9179|false|false|false|C0018792|Heart Atrium|Atrial
Attribute|Clinical Attribute|Principle Diagnosis|9173,9192|false|false|false|C2926591||Atrial fibrillation
Disorder|Disease or Syndrome|Principle Diagnosis|9173,9192|false|false|false|C0004238|Atrial Fibrillation|Atrial fibrillation
Lab|Laboratory or Test Result|Principle Diagnosis|9173,9192|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Atrial fibrillation
Disorder|Disease or Syndrome|Principle Diagnosis|9180,9192|false|false|false|C0232197|Fibrillation|fibrillation
Event|Event|Principle Diagnosis|9180,9192|false|false|false|||fibrillation
Disorder|Disease or Syndrome|Principle Diagnosis|9193,9205|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|Principle Diagnosis|9193,9205|false|false|false|||Hypertension
Disorder|Disease or Syndrome|Principle Diagnosis|9206,9209|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Principle Diagnosis|9206,9209|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Principle Diagnosis|9206,9209|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Principle Diagnosis|9206,9209|false|false|false|||CAD
Finding|Gene or Genome|Principle Diagnosis|9206,9209|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Principle Diagnosis|9206,9209|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Principle Diagnosis|9206,9209|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Principle Diagnosis|9206,9209|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|Discharge Condition|9233,9241|false|false|false|||Deceased
Event|Event|Discharge Instructions|9270,9271|false|false|false|||N
Procedure|Health Care Activity|Discharge Instructions|9276,9284|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|9285,9297|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|9285,9297|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|9285,9297|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

