 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|48,57|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|48,57|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|48,62|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|82,91|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|82,91|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|82,91|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|82,91|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|82,91|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|82,96|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|114,119|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|114,119|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|114,119|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|138,141|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|138,141|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|138,141|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|138,141|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|138,141|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|149,156|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|149,156|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|158,166|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|169,178|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|169,178|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|169,178|false|false|false|C0020517|Hypersensitivity|Allergies
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|181,186|false|false|false|C0749139|sulfa|Sulfa
Event|Event|SIMPLE_SEGMENT|181,186|false|false|false|||Sulfa
Drug|Antibiotic|SIMPLE_SEGMENT|188,199|false|false|false|C0038760;C0599503;C3536763|Sulfonamide Anti-Infective Agents;Sulfonamide [EPC];Sulfonamides|Sulfonamide
Drug|Organic Chemical|SIMPLE_SEGMENT|188,199|false|false|false|C0038760;C0599503;C3536763|Sulfonamide Anti-Infective Agents;Sulfonamide [EPC];Sulfonamides|Sulfonamide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|188,199|false|false|false|C0038760;C0599503;C3536763|Sulfonamide Anti-Infective Agents;Sulfonamide [EPC];Sulfonamides|Sulfonamide
Drug|Antibiotic|SIMPLE_SEGMENT|200,211|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|Antibiotics
Event|Event|SIMPLE_SEGMENT|200,211|false|false|false|||Antibiotics
Drug|Organic Chemical|SIMPLE_SEGMENT|215,222|false|false|false|C0009214|codeine|Codeine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|215,222|false|false|false|C0009214|codeine|Codeine
Drug|Organic Chemical|SIMPLE_SEGMENT|225,232|false|false|false|C0591139|Bactrim|Bactrim
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|225,232|false|false|false|C0591139|Bactrim|Bactrim
Event|Event|SIMPLE_SEGMENT|235,244|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|235,244|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|253,268|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|259,268|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|259,268|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|259,268|false|false|false|C5441521|Complaint (finding)|Complaint
Event|Event|SIMPLE_SEGMENT|271,279|false|false|false|||Weakness
Finding|Sign or Symptom|SIMPLE_SEGMENT|271,279|false|false|false|C0004093;C3714552|Asthenia;Weakness|Weakness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|281,287|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|281,287|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|281,287|false|false|false|C0027497|Nausea|nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|281,296|false|false|false|C0027498|Nausea and vomiting|nausea/vomiting
Event|Event|SIMPLE_SEGMENT|288,296|false|false|false|||vomiting
Finding|Sign or Symptom|SIMPLE_SEGMENT|288,296|false|false|false|C0042963|Vomiting|vomiting
Finding|Classification|SIMPLE_SEGMENT|302,307|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|308,316|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|308,316|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|320,338|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|329,338|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|329,338|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|329,338|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|329,338|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|329,338|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|SIMPLE_SEGMENT|348,355|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|348,355|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|348,355|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|348,355|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|348,358|false|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|348,374|false|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|348,374|false|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|359,366|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|359,366|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|359,374|false|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|367,374|false|false|false|C0221423|Illness (finding)|Illness
Event|Event|SIMPLE_SEGMENT|393,394|false|false|false|||f
Event|Event|SIMPLE_SEGMENT|413,422|false|false|false|||diagnosed
Finding|Functional Concept|SIMPLE_SEGMENT|423,433|false|false|false|C0036525;C1522484|Metastatic to;metastatic qualifier|metastatic
Disorder|Neoplastic Process|SIMPLE_SEGMENT|423,440|false|false|false|C0027627;C0346957;C2939419|Disseminated Malignant Neoplasm;Metastatic malignant neoplasm;Neoplasm Metastasis|metastatic cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|434,440|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|SIMPLE_SEGMENT|434,440|false|false|false|||cancer
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|445,452|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Immunologic Factor|SIMPLE_SEGMENT|445,452|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|445,452|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Event|Event|SIMPLE_SEGMENT|445,452|false|false|false|||unknown
Finding|Finding|SIMPLE_SEGMENT|445,452|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Functional Concept|SIMPLE_SEGMENT|445,452|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Idea or Concept|SIMPLE_SEGMENT|445,452|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Intellectual Product|SIMPLE_SEGMENT|445,452|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Event|Event|SIMPLE_SEGMENT|459,469|false|false|false|||presenting
Finding|Idea or Concept|SIMPLE_SEGMENT|459,469|false|false|false|C0449450|Presentation|presenting
Attribute|Clinical Attribute|SIMPLE_SEGMENT|475,481|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|475,481|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|475,481|false|false|false|C0027497|Nausea|nausea
Event|Event|SIMPLE_SEGMENT|483,491|false|false|false|||vomiting
Finding|Sign or Symptom|SIMPLE_SEGMENT|483,491|false|false|false|C0042963|Vomiting|vomiting
Event|Event|SIMPLE_SEGMENT|497,502|false|false|false|||fever
Finding|Finding|SIMPLE_SEGMENT|497,502|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|497,502|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Body Substance|SIMPLE_SEGMENT|518,525|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|518,525|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|518,525|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Functional Concept|SIMPLE_SEGMENT|518,529|false|false|false|C0332310|Has patient|Patient has
Event|Event|SIMPLE_SEGMENT|535,543|false|false|false|||vomiting
Finding|Sign or Symptom|SIMPLE_SEGMENT|535,543|false|false|false|C0042963|Vomiting|vomiting
Event|Event|SIMPLE_SEGMENT|593,602|false|false|false|||diagnosed
Finding|Functional Concept|SIMPLE_SEGMENT|608,618|false|false|false|C0036525;C1522484|Metastatic to;metastatic qualifier|metastatic
Disorder|Neoplastic Process|SIMPLE_SEGMENT|608,625|false|false|false|C0027627;C0346957;C2939419|Disseminated Malignant Neoplasm;Metastatic malignant neoplasm;Neoplasm Metastasis|metastatic cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|619,625|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|SIMPLE_SEGMENT|619,625|false|false|false|||cancer
Event|Event|SIMPLE_SEGMENT|637,644|false|false|false|||reports
Attribute|Clinical Attribute|SIMPLE_SEGMENT|645,649|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|645,649|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|645,649|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|645,649|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Location or Region|SIMPLE_SEGMENT|659,672|false|false|false|C0230165;C2937240|Upper abdomen (surface region);Upper abdomen structure|upper abdomen
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|659,672|false|false|false|C0230165;C2937240|Upper abdomen (surface region);Upper abdomen structure|upper abdomen
Anatomy|Body Location or Region|SIMPLE_SEGMENT|665,672|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|665,672|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Finding|Finding|SIMPLE_SEGMENT|665,672|false|false|false|C0941288|Abdomen problem|abdomen
Anatomy|Body Location or Region|SIMPLE_SEGMENT|665,676|false|false|false|C0000726|Abdomen|abdomen and
Finding|Finding|SIMPLE_SEGMENT|681,690|false|false|false|C3641766|Very Poor|very poor
Finding|Intellectual Product|SIMPLE_SEGMENT|686,690|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Event|Event|SIMPLE_SEGMENT|694,700|false|false|false|||intake
Finding|Functional Concept|SIMPLE_SEGMENT|694,700|false|false|false|C1512806|Intake|intake
Procedure|Health Care Activity|SIMPLE_SEGMENT|694,700|false|false|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|intake
Event|Event|SIMPLE_SEGMENT|716,723|false|false|false|||feeling
Event|Event|SIMPLE_SEGMENT|738,742|false|false|false|||weak
Finding|Intellectual Product|SIMPLE_SEGMENT|738,742|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|weak
Finding|Sign or Symptom|SIMPLE_SEGMENT|738,742|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|weak
Finding|Finding|SIMPLE_SEGMENT|753,757|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|753,757|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|753,757|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|SIMPLE_SEGMENT|758,764|false|false|false|||period
Finding|Organism Function|SIMPLE_SEGMENT|758,764|false|false|false|C0025344|Menstruation|period
Procedure|Research Activity|SIMPLE_SEGMENT|758,764|false|false|false|C2347804|Clinical Trial Period|period
Event|Event|SIMPLE_SEGMENT|771,779|false|false|false|||vomiting
Finding|Sign or Symptom|SIMPLE_SEGMENT|771,779|false|false|false|C0042963|Vomiting|vomiting
Anatomy|Body Location or Region|SIMPLE_SEGMENT|784,793|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|SIMPLE_SEGMENT|784,798|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|794,798|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|794,798|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|794,798|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|794,798|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|807,816|false|false|false|||increased
Event|Event|SIMPLE_SEGMENT|852,857|false|false|false|||feels
Event|Event|SIMPLE_SEGMENT|863,871|false|false|false|||fatigued
Finding|Sign or Symptom|SIMPLE_SEGMENT|863,871|false|false|false|C0015672|Fatigue|fatigued
Event|Event|SIMPLE_SEGMENT|883,890|false|false|false|||chronic
Finding|Intellectual Product|SIMPLE_SEGMENT|883,890|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|883,890|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Drug|Organic Chemical|SIMPLE_SEGMENT|907,912|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|907,912|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|SIMPLE_SEGMENT|907,912|false|false|false|||cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|907,912|false|false|false|C0010200|Coughing|cough
Finding|Finding|SIMPLE_SEGMENT|916,920|false|false|false|C5575035|Well (answer to question)|well
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|925,928|false|false|false|C0041912|Upper Respiratory Infections|URI
Event|Event|SIMPLE_SEGMENT|925,928|false|false|false|||URI
Finding|Gene or Genome|SIMPLE_SEGMENT|925,928|false|false|false|C1421895;C1548524;C3272713|URI1 gene;URI1 wt Allele;Uniform Resource Identifier|URI
Finding|Intellectual Product|SIMPLE_SEGMENT|925,928|false|false|false|C1421895;C1548524;C3272713|URI1 gene;URI1 wt Allele;Uniform Resource Identifier|URI
Event|Event|SIMPLE_SEGMENT|929,937|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|929,937|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|929,937|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|942,949|false|false|false|C0042027|Urinary tract|urinary
Event|Event|SIMPLE_SEGMENT|951,961|false|false|false|||complaints
Finding|Finding|SIMPLE_SEGMENT|951,961|false|false|false|C5441521|Complaint (finding)|complaints
Event|Event|SIMPLE_SEGMENT|976,987|false|false|false|||constipated
Finding|Sign or Symptom|SIMPLE_SEGMENT|976,987|false|false|false|C0009806|Constipation|constipated
Event|Event|SIMPLE_SEGMENT|995,1003|false|false|false|||improves
Event|Event|SIMPLE_SEGMENT|1014,1019|false|false|false|||stops
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1024,1036|false|false|false|C0003297|Antiemetics|anti-emetics
Event|Event|SIMPLE_SEGMENT|1024,1036|false|false|false|||anti-emetics
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1043,1048|false|false|false|C0021853|Intestines|bowel
Finding|Organism Function|SIMPLE_SEGMENT|1043,1057|false|false|false|C0011135|Defecation|bowel movement
Event|Event|SIMPLE_SEGMENT|1049,1057|false|false|false|||movement
Finding|Organism Function|SIMPLE_SEGMENT|1049,1057|false|false|false|C0026649|Movement|movement
Event|Event|SIMPLE_SEGMENT|1062,1071|false|false|false|||yesterday
Event|Event|SIMPLE_SEGMENT|1081,1088|false|false|false|||passing
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1089,1092|false|false|false|C0017110;C1550641;C1704673|Gas - SpecimenType;Gas Dosage Form;Gases|gas
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|1089,1092|false|false|false|C0017110;C1550641;C1704673|Gas - SpecimenType;Gas Dosage Form;Gases|gas
Drug|Substance|SIMPLE_SEGMENT|1089,1092|false|false|false|C0017110;C1550641;C1704673|Gas - SpecimenType;Gas Dosage Form;Gases|gas
Event|Event|SIMPLE_SEGMENT|1089,1092|false|false|false|||gas
Finding|Gene or Genome|SIMPLE_SEGMENT|1089,1092|false|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|gas
Finding|Intellectual Product|SIMPLE_SEGMENT|1089,1092|false|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|gas
Finding|Molecular Function|SIMPLE_SEGMENT|1089,1092|false|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|gas
Finding|Sign or Symptom|SIMPLE_SEGMENT|1089,1092|false|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|gas
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1102,1107|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|1102,1107|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1102,1117|false|false|false|C0023216|Lower Extremity|lower extremity
Finding|Pathologic Function|SIMPLE_SEGMENT|1102,1123|false|false|false|C0239340|Edema of lower extremity|lower extremity edema
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1108,1117|false|false|false|C0015385|Limb structure|extremity
Finding|Pathologic Function|SIMPLE_SEGMENT|1108,1123|false|false|false|C0085649|Peripheral edema|extremity edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1118,1123|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|1118,1123|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|1118,1123|false|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|1141,1148|false|false|false|||present
Finding|Finding|SIMPLE_SEGMENT|1141,1148|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|SIMPLE_SEGMENT|1141,1148|false|false|false|C0150312;C0449450|Present;Presentation|present
Event|Event|SIMPLE_SEGMENT|1196,1204|false|false|false|||supposed
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1224,1229|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1224,1229|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1224,1229|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|SIMPLE_SEGMENT|1224,1229|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1224,1229|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|SIMPLE_SEGMENT|1224,1229|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Finding|Finding|SIMPLE_SEGMENT|1224,1229|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|SIMPLE_SEGMENT|1224,1229|false|false|false|C0872387|Procedures on liver|liver
Event|Event|SIMPLE_SEGMENT|1230,1234|false|false|false|||mets
Finding|Gene or Genome|SIMPLE_SEGMENT|1230,1234|false|false|false|C0812270;C1705694|ETV3 gene;ETV3 wt Allele|mets
Event|Event|SIMPLE_SEGMENT|1235,1243|false|false|false|||biopsied
Event|Event|SIMPLE_SEGMENT|1284,1290|false|false|false|||taking
Drug|Organic Chemical|SIMPLE_SEGMENT|1291,1300|false|false|false|C0020740|ibuprofen|ibuprofen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1291,1300|false|false|false|C0020740|ibuprofen|ibuprofen
Event|Event|SIMPLE_SEGMENT|1291,1300|false|false|false|||ibuprofen
Event|Event|SIMPLE_SEGMENT|1309,1315|false|false|false|||biopsy
Finding|Finding|SIMPLE_SEGMENT|1309,1315|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Finding|Intellectual Product|SIMPLE_SEGMENT|1309,1315|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1309,1315|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Procedure|Health Care Activity|SIMPLE_SEGMENT|1309,1315|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Event|Event|SIMPLE_SEGMENT|1326,1335|false|false|false|||postponed
Finding|Idea or Concept|SIMPLE_SEGMENT|1352,1359|false|false|false|C1555582|Initial (abbreviation)|initial
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1396,1400|false|false|false|C0587081|Laboratory test finding|Labs
Event|Event|SIMPLE_SEGMENT|1407,1418|false|false|false|||significant
Finding|Idea or Concept|SIMPLE_SEGMENT|1407,1418|false|false|false|C0750502|Significant|significant
Anatomy|Cell|SIMPLE_SEGMENT|1423,1426|false|false|false|C0023516|Leukocytes|WBC
Event|Event|SIMPLE_SEGMENT|1423,1426|false|false|false|||WBC
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|1445,1450|false|false|false|C0032400;C0071360|5'-Inosinic acid, 2'-deoxy-2'-fluoro-, homopolymer;Poly A|polys
Event|Event|SIMPLE_SEGMENT|1445,1450|false|false|false|||polys
Event|Event|SIMPLE_SEGMENT|1452,1454|false|false|false|||UA
Event|Event|SIMPLE_SEGMENT|1459,1470|false|false|false|||significant
Finding|Idea or Concept|SIMPLE_SEGMENT|1459,1470|false|false|false|C0750502|Significant|significant
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|1476,1483|false|false|false|C0497010|Toxic effect of ketones|ketones
Drug|Organic Chemical|SIMPLE_SEGMENT|1476,1483|false|false|false|C0022634|Ketones|ketones
Event|Event|SIMPLE_SEGMENT|1476,1483|false|false|false|||ketones
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1476,1483|false|false|false|C0202110;C0555179|Ketone bodies measurement, quantitative;Urine ketone test|ketones
Finding|Body Substance|SIMPLE_SEGMENT|1485,1492|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1485,1492|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1485,1492|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Organic Chemical|SIMPLE_SEGMENT|1502,1508|false|false|false|C0206046|Zofran|zofran
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1502,1508|false|false|false|C0206046|Zofran|zofran
Event|Event|SIMPLE_SEGMENT|1502,1508|false|false|false|||zofran
Event|Event|SIMPLE_SEGMENT|1510,1512|false|false|false|||NS
Event|Event|SIMPLE_SEGMENT|1524,1527|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1524,1527|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|SIMPLE_SEGMENT|1534,1540|false|false|false|||showed
Finding|Finding|SIMPLE_SEGMENT|1541,1544|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|1541,1544|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Functional Concept|SIMPLE_SEGMENT|1545,1549|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Event|Event|SIMPLE_SEGMENT|1556,1563|false|false|false|||opacity
Finding|Finding|SIMPLE_SEGMENT|1556,1563|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacity
Finding|Pathologic Function|SIMPLE_SEGMENT|1556,1563|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacity
Event|Event|SIMPLE_SEGMENT|1573,1580|false|false|false|||reflect
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|1581,1584|false|false|false|C0600500|Peptide Nucleic Acids|PNA
Event|Event|SIMPLE_SEGMENT|1581,1584|false|false|false|||PNA
Event|Event|SIMPLE_SEGMENT|1585,1597|false|false|false|||superimposed
Finding|Functional Concept|SIMPLE_SEGMENT|1602,1612|false|false|false|C0036525;C1522484|Metastatic to;metastatic qualifier|metastatic
Event|Event|SIMPLE_SEGMENT|1613,1619|false|false|false|||diseae
Event|Activity|SIMPLE_SEGMENT|1638,1644|false|false|false|C1947932|Smear - instruction imperative|spread
Event|Event|SIMPLE_SEGMENT|1638,1644|false|false|false|||spread
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1648,1654|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|SIMPLE_SEGMENT|1648,1654|false|false|false|||cancer
Event|Event|SIMPLE_SEGMENT|1670,1674|false|false|false|||vanc
Drug|Antibiotic|SIMPLE_SEGMENT|1679,1687|false|false|false|C0055003|cefepime|cefepime
Drug|Organic Chemical|SIMPLE_SEGMENT|1679,1687|false|false|false|C0055003|cefepime|cefepime
Event|Event|SIMPLE_SEGMENT|1679,1687|false|false|false|||cefepime
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1692,1701|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|SIMPLE_SEGMENT|1692,1701|false|false|false|||pneumonia
Event|Event|SIMPLE_SEGMENT|1703,1709|false|false|false|||Vitals
Event|Event|SIMPLE_SEGMENT|1713,1721|false|false|false|||transfer
Finding|Functional Concept|SIMPLE_SEGMENT|1713,1721|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|SIMPLE_SEGMENT|1713,1721|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|SIMPLE_SEGMENT|1713,1721|false|false|false|C4706767|Transfer (immobility management)|transfer
Event|Event|SIMPLE_SEGMENT|1769,1778|false|false|false|||continues
Event|Event|SIMPLE_SEGMENT|1782,1786|false|false|false|||feel
Finding|Intellectual Product|SIMPLE_SEGMENT|1782,1791|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|feel weak
Finding|Sign or Symptom|SIMPLE_SEGMENT|1782,1791|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|feel weak
Event|Event|SIMPLE_SEGMENT|1787,1791|false|false|false|||weak
Finding|Intellectual Product|SIMPLE_SEGMENT|1787,1791|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|weak
Finding|Sign or Symptom|SIMPLE_SEGMENT|1787,1791|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|weak
Event|Event|SIMPLE_SEGMENT|1796,1804|false|false|false|||nauseous
Finding|Sign or Symptom|SIMPLE_SEGMENT|1796,1804|false|false|false|C0027497|Nausea|nauseous
Event|Event|SIMPLE_SEGMENT|1814,1820|false|false|false|||trying
Event|Event|SIMPLE_SEGMENT|1824,1828|false|false|false|||take
Event|Event|SIMPLE_SEGMENT|1833,1838|false|false|false|||pants
Finding|Gene or Genome|SIMPLE_SEGMENT|1833,1838|false|false|false|C2240332|C22orf39 gene|pants
Event|Event|SIMPLE_SEGMENT|1848,1853|false|false|false|||feels
Event|Event|SIMPLE_SEGMENT|1858,1862|false|false|false|||weak
Finding|Intellectual Product|SIMPLE_SEGMENT|1858,1862|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|weak
Finding|Sign or Symptom|SIMPLE_SEGMENT|1858,1862|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|weak
Event|Event|SIMPLE_SEGMENT|1867,1872|false|false|false|||tired
Finding|Finding|SIMPLE_SEGMENT|1867,1872|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Finding|Intellectual Product|SIMPLE_SEGMENT|1867,1872|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Finding|Sign or Symptom|SIMPLE_SEGMENT|1867,1872|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Event|Event|SIMPLE_SEGMENT|1886,1892|false|false|false|||REVIEW
Finding|Idea or Concept|SIMPLE_SEGMENT|1886,1892|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|REVIEW
Finding|Intellectual Product|SIMPLE_SEGMENT|1886,1892|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|REVIEW
Finding|Functional Concept|SIMPLE_SEGMENT|1886,1895|false|false|false|C0699752|Review of|REVIEW OF
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1886,1903|false|false|false|C0488564;C0488565||REVIEW OF SYSTEMS
Procedure|Health Care Activity|SIMPLE_SEGMENT|1886,1903|false|false|false|C0489633|Review of systems (procedure)|REVIEW OF SYSTEMS
Event|Event|SIMPLE_SEGMENT|1896,1903|false|false|false|||SYSTEMS
Finding|Functional Concept|SIMPLE_SEGMENT|1896,1903|false|false|false|C0449913|System|SYSTEMS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1915,1918|false|false|false|C0268529|Proline dehydrogenase deficiency|HPI
Event|Event|SIMPLE_SEGMENT|1915,1918|false|false|false|||HPI
Finding|Finding|SIMPLE_SEGMENT|1915,1918|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Finding|Molecular Function|SIMPLE_SEGMENT|1915,1918|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Finding|Sign or Symptom|SIMPLE_SEGMENT|1925,1937|false|false|false|C0028081|Night sweats|night sweats
Event|Event|SIMPLE_SEGMENT|1931,1937|false|false|false|||sweats
Finding|Body Substance|SIMPLE_SEGMENT|1931,1937|false|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Finding|Finding|SIMPLE_SEGMENT|1931,1937|false|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Event|Event|SIMPLE_SEGMENT|1939,1947|false|false|false|||headache
Finding|Sign or Symptom|SIMPLE_SEGMENT|1939,1947|false|false|false|C0018681|Headache|headache
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1949,1955|false|false|false|C2707266||vision
Finding|Organism Function|SIMPLE_SEGMENT|1949,1955|false|false|false|C0042789|Vision|vision
Event|Event|SIMPLE_SEGMENT|1956,1963|false|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|1956,1963|false|false|false|C0392747|Changing|changes
Event|Event|SIMPLE_SEGMENT|1965,1975|false|false|false|||rhinorrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1965,1975|false|false|false|C1260880|Rhinorrhea|rhinorrhea
Event|Event|SIMPLE_SEGMENT|1978,1988|false|false|false|||congestion
Finding|Pathologic Function|SIMPLE_SEGMENT|1978,1988|false|false|false|C0700148|Congestion|congestion
Finding|Sign or Symptom|SIMPLE_SEGMENT|1990,1994|false|false|false|C0234233;C1442877|Sore skin;Sore to touch|sore
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1990,2001|false|false|false|C0031350|Pharyngitis|sore throat
Drug|Organic Chemical|SIMPLE_SEGMENT|1990,2001|false|false|false|C0723402;C3244654|Sore Throat brand of Phenol;Sore Throat brand of benzocaine & menthol|sore throat
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1990,2001|false|false|false|C0723402;C3244654|Sore Throat brand of Phenol;Sore Throat brand of benzocaine & menthol|sore throat
Finding|Sign or Symptom|SIMPLE_SEGMENT|1990,2001|false|false|false|C0242429|Sore Throat|sore throat
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1995,2001|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1995,2001|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1995,2001|false|false|false|C1950455|Throat Homeopathic Medication|throat
Event|Event|SIMPLE_SEGMENT|1995,2001|false|false|false|||throat
Finding|Body Substance|SIMPLE_SEGMENT|1995,2001|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Finding|Intellectual Product|SIMPLE_SEGMENT|1995,2001|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2003,2008|false|false|false|C0018932|Hematochezia|BRBPR
Event|Event|SIMPLE_SEGMENT|2003,2008|false|false|false|||BRBPR
Event|Event|SIMPLE_SEGMENT|2010,2016|false|false|false|||melena
Finding|Pathologic Function|SIMPLE_SEGMENT|2010,2016|false|false|false|C0025222|Melena|melena
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2018,2030|false|false|false|C0018932|Hematochezia|hematochezia
Event|Event|SIMPLE_SEGMENT|2018,2030|false|false|false|||hematochezia
Finding|Sign or Symptom|SIMPLE_SEGMENT|2018,2030|false|false|false|C1321898|Blood in stool|hematochezia
Event|Event|SIMPLE_SEGMENT|2032,2039|false|false|false|||dysuria
Finding|Sign or Symptom|SIMPLE_SEGMENT|2032,2039|false|false|false|C0013428|Dysuria|dysuria
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2042,2051|false|false|false|C0018965|Hematuria|hematuria
Event|Event|SIMPLE_SEGMENT|2042,2051|false|false|false|||hematuria
Finding|Finding|SIMPLE_SEGMENT|2060,2080|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|2065,2072|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|2065,2072|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|2065,2072|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|2065,2072|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2065,2072|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|2065,2080|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2073,2080|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2073,2080|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2073,2080|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Event|Event|SIMPLE_SEGMENT|2082,2085|false|false|false|||PMH
Finding|Finding|SIMPLE_SEGMENT|2082,2085|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|PMH
Finding|Finding|SIMPLE_SEGMENT|2090,2094|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|SIMPLE_SEGMENT|2090,2094|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|SIMPLE_SEGMENT|2090,2094|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Finding|SIMPLE_SEGMENT|2090,2100|false|false|false|C0205082;C4554016|Enneking High Surgical Grade;Severe (severity modifier)|high grade
Finding|Intellectual Product|SIMPLE_SEGMENT|2090,2100|false|false|false|C0205082;C4554016|Enneking High Surgical Grade;Severe (severity modifier)|high grade
Finding|Classification|SIMPLE_SEGMENT|2095,2100|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Finding|Finding|SIMPLE_SEGMENT|2095,2100|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Event|Event|SIMPLE_SEGMENT|2101,2104|false|false|false|||SBO
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2113,2135|false|false|false|C0085704|Exploratory laparotomy|exploratory laparotomy
Event|Event|SIMPLE_SEGMENT|2125,2135|false|false|false|||laparotomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2125,2135|false|false|false|C0023038|Laparotomy|laparotomy
Event|Event|SIMPLE_SEGMENT|2137,2142|false|false|false|||lysis
Finding|Cell Function|SIMPLE_SEGMENT|2137,2142|false|false|false|C0024348;C1536403|Lysis;pathologic cytolysis|lysis
Finding|Pathologic Function|SIMPLE_SEGMENT|2137,2142|false|false|false|C0024348;C1536403|Lysis;pathologic cytolysis|lysis
Event|Event|SIMPLE_SEGMENT|2147,2156|false|false|false|||adhesions
Finding|Pathologic Function|SIMPLE_SEGMENT|2147,2156|false|false|false|C0001511|Tissue Adhesions|adhesions
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2162,2173|false|false|false|C0021852;C4319010|Abdomen>Small bowel;Intestines, Small|small bowel
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2162,2173|false|false|false|C0021852;C4319010|Abdomen>Small bowel;Intestines, Small|small bowel
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2162,2183|false|false|false|C0192601|Small intestine excision|small bowel resection
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2168,2173|false|false|false|C0021853|Intestines|bowel
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2168,2183|false|false|false|C0741614|Bowel resection|bowel resection
Event|Event|SIMPLE_SEGMENT|2174,2183|false|false|false|||resection
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2174,2183|false|false|false|C0015252;C0728940|Excision;removal technique|resection
Event|Event|SIMPLE_SEGMENT|2189,2206|false|false|false|||enteroenterostomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2189,2206|false|false|false|C0192711;C0192741|Anastomosis of intestine;Anastomosis of small intestine to small intestine|enteroenterostomy
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2210,2219|false|false|false|C0007095|Carcinoid Tumor|carcinoid
Event|Event|SIMPLE_SEGMENT|2210,2219|false|false|false|||carcinoid
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2222,2236|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|hyperlipidemia
Event|Event|SIMPLE_SEGMENT|2222,2236|false|false|false|||hyperlipidemia
Finding|Finding|SIMPLE_SEGMENT|2222,2236|false|false|false|C0428465|Serum lipids high (finding)|hyperlipidemia
Drug|Organic Chemical|SIMPLE_SEGMENT|2239,2246|false|false|false|C0042890|Vitamins|vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2239,2246|false|false|false|C0042890|Vitamins|vitamin
Drug|Vitamin|SIMPLE_SEGMENT|2239,2246|false|false|false|C0042890|Vitamins|vitamin
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|2239,2250|false|false|false|C0042845;C0086024;C2936883|Vitamin B12 [EPC];cobalamins;vitamin B12|vitamin B12
Drug|Organic Chemical|SIMPLE_SEGMENT|2239,2250|false|false|false|C0042845;C0086024;C2936883|Vitamin B12 [EPC];cobalamins;vitamin B12|vitamin B12
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2239,2250|false|false|false|C0042845;C0086024;C2936883|Vitamin B12 [EPC];cobalamins;vitamin B12|vitamin B12
Drug|Vitamin|SIMPLE_SEGMENT|2239,2250|false|false|false|C0042845;C0086024;C2936883|Vitamin B12 [EPC];cobalamins;vitamin B12|vitamin B12
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2239,2250|false|false|false|C0202252|VITAMIN B12 MEASUREMENT|vitamin B12
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2239,2261|false|false|false|C0042847|Vitamin B 12 Deficiency|vitamin B12 deficiency
Finding|Finding|SIMPLE_SEGMENT|2239,2261|false|false|false|C5886863|Decreased circulating vitamin B12 concentration|vitamin B12 deficiency
Event|Event|SIMPLE_SEGMENT|2247,2250|false|false|false|||B12
Finding|Gene or Genome|SIMPLE_SEGMENT|2247,2250|false|false|false|C1417635;C1420797;C3538796|NDUFB3 gene;TNFAIP1 gene;TNFAIP1 wt Allele|B12
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2251,2261|false|false|false|C0162429|Malnutrition|deficiency
Event|Event|SIMPLE_SEGMENT|2251,2261|false|false|false|||deficiency
Finding|Functional Concept|SIMPLE_SEGMENT|2251,2261|false|false|false|C0011155|Deficiency|deficiency
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2264,2272|false|false|false|C0027530|Neck|cervical
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2273,2276|false|false|false|C0029408|Degenerative polyarthritis|DJD
Event|Event|SIMPLE_SEGMENT|2273,2276|false|false|false|||DJD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2279,2293|false|false|false|C0029408|Degenerative polyarthritis|osteoarthritis
Event|Event|SIMPLE_SEGMENT|2279,2293|false|false|false|||osteoarthritis
Event|Event|SIMPLE_SEGMENT|2296,2299|false|false|false|||PSH
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2308,2312|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2308,2312|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2308,2312|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|2308,2312|false|false|false|C0740941|Lung Problem|lung
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2308,2322|false|false|false|C0396565|Lung excision|lung resection
Event|Event|SIMPLE_SEGMENT|2313,2322|false|false|false|||resection
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2313,2322|false|false|false|C0015252;C0728940|Excision;removal technique|resection
Event|Event|SIMPLE_SEGMENT|2341,2353|false|false|false|||hysterectomy
Finding|Finding|SIMPLE_SEGMENT|2341,2353|false|false|false|C1548863|Consent Type - Hysterectomy|hysterectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2341,2353|false|false|false|C0020699|Hysterectomy|hysterectomy
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2365,2370|false|false|false|C4048756|Right arm|R arm
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2367,2370|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|2367,2370|false|false|false|C3495676|Anorectal Malformations|arm
Finding|Gene or Genome|SIMPLE_SEGMENT|2367,2370|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2367,2370|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|SIMPLE_SEGMENT|2367,2370|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2367,2370|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Event|Event|SIMPLE_SEGMENT|2371,2378|false|false|false|||surgery
Finding|Finding|SIMPLE_SEGMENT|2371,2378|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|2371,2378|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|2371,2378|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2371,2378|false|false|false|C0543467|Operative Surgical Procedures|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|2382,2388|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|2382,2396|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|2389,2396|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2389,2396|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2389,2396|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2389,2396|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|2402,2408|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2402,2408|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|2402,2408|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|2402,2408|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|2402,2416|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|2409,2416|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2409,2416|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2409,2416|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2409,2416|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Idea or Concept|SIMPLE_SEGMENT|2418,2424|false|false|false|C1546508|Relationship - Mother|Mother
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2431,2437|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|SIMPLE_SEGMENT|2431,2437|false|false|false|||cancer
Event|Event|SIMPLE_SEGMENT|2475,2480|false|false|false|||touch
Finding|Mental Process|SIMPLE_SEGMENT|2475,2480|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|2475,2480|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2475,2480|false|false|false|C0152054|Therapeutic Touch|touch
Event|Event|SIMPLE_SEGMENT|2486,2494|false|false|false|||siblings
Finding|Conceptual Entity|SIMPLE_SEGMENT|2497,2503|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|SIMPLE_SEGMENT|2497,2503|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Event|Event|SIMPLE_SEGMENT|2525,2533|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|2525,2533|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|2525,2533|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2525,2533|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|2525,2538|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2525,2538|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|2534,2538|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|2534,2538|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2534,2538|false|false|false|C0582103|Medical Examination|Exam
Event|Event|SIMPLE_SEGMENT|2540,2549|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|2540,2549|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Finding|Finding|SIMPLE_SEGMENT|2550,2558|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|2550,2558|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2550,2558|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|2550,2563|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2550,2563|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|2559,2563|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|2559,2563|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2559,2563|false|false|false|C0582103|Medical Examination|Exam
Event|Event|SIMPLE_SEGMENT|2605,2612|false|false|false|||GENERAL
Finding|Classification|SIMPLE_SEGMENT|2605,2612|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|2605,2612|false|false|false|C3812897|General medical service|GENERAL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2614,2619|false|false|false|C0028754|Obesity|Obese
Event|Event|SIMPLE_SEGMENT|2635,2646|false|false|false|||comfortable
Finding|Finding|SIMPLE_SEGMENT|2635,2646|false|false|false|C5546696|Feeling comfortable|comfortable
Finding|Finding|SIMPLE_SEGMENT|2648,2668|false|false|false|C2051415|patient appears in no acute distress (physical finding)|in no acute distress
Finding|Intellectual Product|SIMPLE_SEGMENT|2654,2659|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|SIMPLE_SEGMENT|2660,2668|false|false|false|||distress
Finding|Finding|SIMPLE_SEGMENT|2660,2668|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|SIMPLE_SEGMENT|2660,2668|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2672,2677|false|false|false|C1512338|HEENT|HEENT
Event|Event|SIMPLE_SEGMENT|2679,2685|false|false|false|||PERRLA
Finding|Finding|SIMPLE_SEGMENT|2679,2685|false|false|false|C2143306|PERRLA|PERRLA
Event|Event|SIMPLE_SEGMENT|2687,2691|false|false|false|||EOMI
Event|Event|SIMPLE_SEGMENT|2701,2710|false|false|false|||anicteric
Finding|Finding|SIMPLE_SEGMENT|2701,2710|false|false|false|C0205180|Anicteric|anicteric
Event|Event|SIMPLE_SEGMENT|2725,2730|false|false|false|||mucus
Finding|Body Substance|SIMPLE_SEGMENT|2725,2730|false|false|false|C0026727;C1546714;C2753459|Mucus (substance);mucus layer|mucus
Finding|Intellectual Product|SIMPLE_SEGMENT|2725,2730|false|false|false|C0026727;C1546714;C2753459|Mucus (substance);mucus layer|mucus
Anatomy|Tissue|SIMPLE_SEGMENT|2732,2741|false|false|false|C0025255|Membrane Tissue|membranes
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2744,2748|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|SIMPLE_SEGMENT|2744,2748|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|SIMPLE_SEGMENT|2744,2748|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|SIMPLE_SEGMENT|2750,2756|false|false|false|||supple
Finding|Functional Concept|SIMPLE_SEGMENT|2750,2756|false|false|false|C0332254|Supple|supple
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2758,2763|false|false|false|C0028754|Obesity|obese
Event|Event|SIMPLE_SEGMENT|2758,2763|false|false|false|||obese
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2766,2771|false|false|false|C0024109|Lung|LUNGS
Finding|Pathologic Function|SIMPLE_SEGMENT|2773,2780|false|false|false|C5441917|Distant Metastasis|Distant
Finding|Body Substance|SIMPLE_SEGMENT|2781,2787|false|false|false|C0225386|Breath|breath
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2781,2794|false|false|false|C0035234;C3484186|Respiratory Sounds|breath sounds
Event|Event|SIMPLE_SEGMENT|2788,2794|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2788,2794|false|false|false|C0037709||sounds
Event|Event|SIMPLE_SEGMENT|2796,2805|false|false|false|||decreased
Finding|Functional Concept|SIMPLE_SEGMENT|2813,2818|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Event|Event|SIMPLE_SEGMENT|2825,2833|false|false|false|||crackles
Finding|Finding|SIMPLE_SEGMENT|2825,2833|false|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2840,2845|false|false|false|C0018787;C4037974|Chest>Heart;Heart|HEART
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2840,2845|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|HEART
Event|Event|SIMPLE_SEGMENT|2840,2845|false|false|false|||HEART
Finding|Sign or Symptom|SIMPLE_SEGMENT|2840,2845|false|false|false|C0795691|HEART PROBLEM|HEART
Event|Event|SIMPLE_SEGMENT|2847,2850|false|false|false|||RRR
Event|Event|SIMPLE_SEGMENT|2855,2858|false|false|false|||MRG
Finding|Gene or Genome|SIMPLE_SEGMENT|2855,2858|true|false|false|C1422304|MAS1L gene|MRG
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2871,2878|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2871,2878|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|SIMPLE_SEGMENT|2871,2878|false|false|false|||ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|2871,2878|false|false|false|C0941288|Abdomen problem|ABDOMEN
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2882,2887|false|false|false|C0021853|Intestines|bowel
Finding|Finding|SIMPLE_SEGMENT|2882,2894|false|false|false|C0232693|Bowel sounds|bowel sounds
Event|Event|SIMPLE_SEGMENT|2888,2894|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2888,2894|false|false|false|C0037709||sounds
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2896,2900|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|SIMPLE_SEGMENT|2896,2900|false|false|false|||soft
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2902,2912|false|false|false|C0521440|Epigastric|epigastric
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2917,2920|false|false|false|C0230177|Structure of right upper quadrant of abdomen|RUQ
Event|Event|SIMPLE_SEGMENT|2921,2931|false|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|2921,2931|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|2921,2931|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Event|SIMPLE_SEGMENT|2936,2945|false|false|false|||palpation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2936,2945|false|false|false|C0030247|Palpation|palpation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2956,2964|false|false|false|C1293134|Enlargement procedure|enlarged
Finding|Finding|SIMPLE_SEGMENT|2956,2970|false|false|false|C0019209|Hepatomegaly|enlarged liver
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2965,2970|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2965,2970|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2965,2970|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|SIMPLE_SEGMENT|2965,2970|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2965,2970|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|SIMPLE_SEGMENT|2965,2970|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|SIMPLE_SEGMENT|2965,2970|false|false|false|||liver
Finding|Finding|SIMPLE_SEGMENT|2965,2970|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|SIMPLE_SEGMENT|2965,2970|false|false|false|C0872387|Procedures on liver|liver
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2977,2982|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2977,2982|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2977,2982|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|SIMPLE_SEGMENT|2977,2982|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2977,2982|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|SIMPLE_SEGMENT|2977,2982|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|SIMPLE_SEGMENT|2977,2982|false|false|false|||liver
Finding|Finding|SIMPLE_SEGMENT|2977,2982|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|SIMPLE_SEGMENT|2977,2982|false|false|false|C0872387|Procedures on liver|liver
Finding|Finding|SIMPLE_SEGMENT|2977,2987|false|false|false|C0426689|Liver edge|liver edge
Finding|Finding|SIMPLE_SEGMENT|2977,2996|false|false|false|C0426690|Liver edge palpable|liver edge palpable
Finding|Conceptual Entity|SIMPLE_SEGMENT|2983,2987|false|false|false|C2697523|Graph Edge|edge
Event|Event|SIMPLE_SEGMENT|2988,2996|false|false|false|||palpable
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3009,3012|false|false|false|C0035561|Bone structure of rib|rib
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3009,3017|false|false|false|C0222762|Rib Cage|rib cage
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3013,3017|false|false|false|C4555210|CAGE Antibody|cage
Drug|Immunologic Factor|SIMPLE_SEGMENT|3013,3017|false|false|false|C4555210|CAGE Antibody|cage
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3013,3017|false|false|false|C4555210|CAGE Antibody|cage
Event|Event|SIMPLE_SEGMENT|3013,3017|false|false|false|||cage
Finding|Gene or Genome|SIMPLE_SEGMENT|3013,3017|false|false|false|C1426669|DDX53 gene|cage
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3013,3017|false|false|false|C5552712|CAP Analysis of Gene Expression|cage
Event|Event|SIMPLE_SEGMENT|3022,3029|false|false|false|||rebound
Event|Event|SIMPLE_SEGMENT|3030,3038|false|false|false|||guarding
Finding|Finding|SIMPLE_SEGMENT|3030,3038|true|false|false|C0427198|Protective muscle spasm|guarding
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3042,3053|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3058,3063|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|3058,3063|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3058,3073|false|false|false|C0023216|Lower Extremity|lower extremity
Finding|Pathologic Function|SIMPLE_SEGMENT|3058,3079|false|false|false|C0239340|Edema of lower extremity|lower extremity edema
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3064,3073|false|false|false|C0015385|Limb structure|extremity
Finding|Pathologic Function|SIMPLE_SEGMENT|3064,3079|false|false|false|C0085649|Peripheral edema|extremity edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3074,3079|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|3074,3079|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|3074,3079|false|false|false|C0013604|Edema|edema
Drug|Food|SIMPLE_SEGMENT|3084,3090|false|false|false|C5890763||pulses
Event|Event|SIMPLE_SEGMENT|3084,3090|false|false|false|||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|3084,3090|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|3084,3090|false|false|false|C0034107|Pulse taking|pulses
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3084,3097|false|false|false|C0232142||pulses radial
Event|Event|SIMPLE_SEGMENT|3091,3097|false|false|false|||radial
Finding|Conceptual Entity|SIMPLE_SEGMENT|3091,3097|false|false|false|C0442038;C0920847|Circumpennate;Radial|radial
Event|Event|SIMPLE_SEGMENT|3114,3119|false|false|false|||awake
Finding|Finding|SIMPLE_SEGMENT|3114,3119|false|false|false|C0234422|Awake (finding)|awake
Event|Event|SIMPLE_SEGMENT|3121,3122|false|false|false|||A
Anatomy|Body System|SIMPLE_SEGMENT|3128,3131|false|false|false|C3714787|Central Nervous System|CNs
Finding|Finding|SIMPLE_SEGMENT|3147,3153|false|false|false|C1554187|Gender Status - Intact|intact
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3155,3161|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|SIMPLE_SEGMENT|3155,3161|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3155,3170|false|false|false|C4050373||muscle strength
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3155,3170|false|false|false|C0517349|Muscle Strength|muscle strength
Event|Event|SIMPLE_SEGMENT|3162,3170|false|false|false|||strength
Finding|Idea or Concept|SIMPLE_SEGMENT|3162,3170|false|false|false|C0808080|Strength (attribute)|strength
Event|Event|SIMPLE_SEGMENT|3190,3199|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|3190,3199|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|3190,3199|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|3190,3199|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|3190,3199|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|3200,3208|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|3200,3208|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|3200,3208|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|3200,3213|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3200,3213|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|3209,3213|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|3209,3213|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3209,3213|false|false|false|C0582103|Medical Examination|Exam
Event|Event|SIMPLE_SEGMENT|3260,3267|false|false|false|||General
Finding|Classification|SIMPLE_SEGMENT|3260,3267|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|SIMPLE_SEGMENT|3260,3267|false|false|false|C3812897|General medical service|General
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3269,3274|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|3269,3274|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3269,3274|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|3269,3274|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|3269,3274|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|3269,3274|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|3269,3274|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|3276,3284|false|false|false|||oriented
Finding|Intellectual Product|SIMPLE_SEGMENT|3289,3294|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|SIMPLE_SEGMENT|3295,3303|false|false|false|||distress
Finding|Finding|SIMPLE_SEGMENT|3295,3303|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|SIMPLE_SEGMENT|3295,3303|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3305,3310|false|false|false|C0028754|Obesity|obese
Event|Event|SIMPLE_SEGMENT|3311,3320|false|false|false|||appearing
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3330,3335|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3337,3343|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3337,3343|false|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|SIMPLE_SEGMENT|3337,3343|false|false|false|||Sclera
Procedure|Health Care Activity|SIMPLE_SEGMENT|3337,3343|false|false|false|C2228481|examination of sclera|Sclera
Event|Event|SIMPLE_SEGMENT|3344,3353|false|false|false|||anicteric
Finding|Finding|SIMPLE_SEGMENT|3344,3353|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3355,3358|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3355,3358|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3360,3370|false|false|false|C0521367|Oropharyngeal|oropharynx
Event|Event|SIMPLE_SEGMENT|3371,3376|false|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|3371,3376|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3379,3383|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|SIMPLE_SEGMENT|3379,3383|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|SIMPLE_SEGMENT|3379,3383|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|SIMPLE_SEGMENT|3385,3391|false|false|false|||supple
Finding|Functional Concept|SIMPLE_SEGMENT|3385,3391|false|false|false|C0332254|Supple|supple
Event|Event|SIMPLE_SEGMENT|3393,3396|false|false|false|||JVP
Finding|Finding|SIMPLE_SEGMENT|3393,3396|false|false|false|C0428897|Jugular venous pressure|JVP
Event|Event|SIMPLE_SEGMENT|3401,3409|false|false|false|||elevated
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3414,3417|true|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3414,3417|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|SIMPLE_SEGMENT|3414,3417|false|false|false|||LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|3414,3417|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3420,3425|false|false|false|C0024109|Lung|Lungs
Event|Event|SIMPLE_SEGMENT|3427,3432|false|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|3427,3432|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|3436,3448|false|false|false|||auscultation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3436,3448|false|false|false|C0004339|Auscultation|auscultation
Event|Event|SIMPLE_SEGMENT|3476,3482|false|false|false|||breath
Finding|Body Substance|SIMPLE_SEGMENT|3476,3482|false|false|false|C0225386|Breath|breath
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3484,3489|false|false|false|C0037709||sound
Finding|Functional Concept|SIMPLE_SEGMENT|3493,3497|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3498,3507|false|false|false|C0751438|Posterior pituitary disease|posterior
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3516,3520|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3516,3520|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3516,3520|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|3516,3520|false|false|false|C0740941|Lung Problem|lung
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3516,3526|false|false|false|C0225759|Lung field|lung field
Event|Event|SIMPLE_SEGMENT|3521,3526|false|false|false|||field
Finding|Conceptual Entity|SIMPLE_SEGMENT|3521,3526|false|false|false|C1521738;C2346620;C2349184|Field;Force Field;Knowledge Field|field
Procedure|Health Care Activity|SIMPLE_SEGMENT|3521,3526|false|false|false|C1553496|field - patient encounter|field
Event|Event|SIMPLE_SEGMENT|3531,3538|false|false|false|||wheezes
Finding|Sign or Symptom|SIMPLE_SEGMENT|3531,3538|true|false|false|C0043144|Wheezing|wheezes
Event|Event|SIMPLE_SEGMENT|3540,3545|false|false|false|||rales
Finding|Finding|SIMPLE_SEGMENT|3540,3545|true|false|false|C0034642;C0240859|Basilar Rales;Rales|rales
Event|Activity|SIMPLE_SEGMENT|3569,3573|false|false|false|C0871208|Rating (action)|rate
Event|Event|SIMPLE_SEGMENT|3569,3573|false|false|false|||rate
Finding|Idea or Concept|SIMPLE_SEGMENT|3569,3573|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|SIMPLE_SEGMENT|3578,3584|false|false|false|||rhythm
Finding|Finding|SIMPLE_SEGMENT|3578,3584|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|SIMPLE_SEGMENT|3578,3584|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Event|Event|SIMPLE_SEGMENT|3605,3612|false|false|false|||murmurs
Finding|Finding|SIMPLE_SEGMENT|3605,3612|true|false|false|C0018808|Heart murmur|murmurs
Event|Event|SIMPLE_SEGMENT|3614,3618|false|false|false|||rubs
Finding|Finding|SIMPLE_SEGMENT|3614,3618|true|false|false|C0232267|Pericardial friction rub|rubs
Event|Event|SIMPLE_SEGMENT|3621,3628|false|false|false|||gallops
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3631,3638|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3631,3638|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Finding|Finding|SIMPLE_SEGMENT|3631,3638|false|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3640,3644|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|SIMPLE_SEGMENT|3640,3644|false|false|false|||soft
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3646,3651|false|false|false|C0028754|Obesity|obese
Event|Event|SIMPLE_SEGMENT|3646,3651|false|false|false|||obese
Event|Event|SIMPLE_SEGMENT|3663,3669|false|false|false|||tender
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3686,3691|false|false|false|C0021853|Intestines|bowel
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3693,3699|false|false|false|C0037709||sounds
Event|Event|SIMPLE_SEGMENT|3700,3707|false|false|false|||present
Finding|Finding|SIMPLE_SEGMENT|3700,3707|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|SIMPLE_SEGMENT|3700,3707|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Sign or Symptom|SIMPLE_SEGMENT|3712,3730|true|false|false|C0234246|Rebound tenderness|rebound tenderness
Event|Event|SIMPLE_SEGMENT|3720,3730|false|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|3720,3730|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|3720,3730|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Event|SIMPLE_SEGMENT|3734,3742|false|false|false|||guarding
Finding|Finding|SIMPLE_SEGMENT|3734,3742|true|false|false|C0427198|Protective muscle spasm|guarding
Event|Event|SIMPLE_SEGMENT|3744,3746|false|false|false|||no
Event|Event|SIMPLE_SEGMENT|3748,3760|false|false|false|||organomegaly
Finding|Finding|SIMPLE_SEGMENT|3748,3760|false|false|false|C4054315|Organomegaly|organomegaly
Event|Event|SIMPLE_SEGMENT|3770,3775|false|false|false|||foley
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|3778,3781|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|SIMPLE_SEGMENT|3778,3781|false|false|false|||Ext
Finding|Gene or Genome|SIMPLE_SEGMENT|3778,3781|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|SIMPLE_SEGMENT|3783,3787|false|false|false|||warm
Finding|Finding|SIMPLE_SEGMENT|3783,3787|false|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3783,3787|false|false|false|C0687712|warming process|warm
Finding|Finding|SIMPLE_SEGMENT|3789,3793|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|3794,3802|false|false|false|||perfused
Drug|Food|SIMPLE_SEGMENT|3807,3813|false|false|false|C5890763||pulses
Event|Event|SIMPLE_SEGMENT|3807,3813|false|false|false|||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|3807,3813|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|3807,3813|false|false|false|C0034107|Pulse taking|pulses
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|3818,3826|true|false|false|C0149651|Clubbing|clubbing
Event|Event|SIMPLE_SEGMENT|3818,3826|false|false|false|||clubbing
Event|Event|SIMPLE_SEGMENT|3828,3836|false|false|false|||cyanosis
Finding|Sign or Symptom|SIMPLE_SEGMENT|3828,3836|true|false|false|C0010520|Cyanosis|cyanosis
Finding|Functional Concept|SIMPLE_SEGMENT|3842,3849|false|false|false|C0205323|Pitting|pitting
Finding|Finding|SIMPLE_SEGMENT|3842,3855|false|false|false|C0333243|Pitting edema|pitting edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3850,3855|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|3850,3855|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|3850,3855|false|false|false|C0013604|Edema|edema
Finding|Classification|SIMPLE_SEGMENT|3865,3869|false|false|false|C3899749|CNS 2|CNs2
Event|Event|SIMPLE_SEGMENT|3873,3879|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|3873,3879|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Functional Concept|SIMPLE_SEGMENT|3881,3886|false|false|false|C1513492|motor movement|motor
Finding|Finding|SIMPLE_SEGMENT|3881,3895|false|false|false|C5551447|Motor function (finding)|motor function
Phenomenon|Biologic Function|SIMPLE_SEGMENT|3881,3895|false|false|false|C0234130|Motor function (observable entity)|motor function
Event|Event|SIMPLE_SEGMENT|3887,3895|false|false|false|||function
Finding|Finding|SIMPLE_SEGMENT|3887,3895|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|3887,3895|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|3887,3895|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|SIMPLE_SEGMENT|3887,3895|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Event|Event|SIMPLE_SEGMENT|3904,3910|false|false|false|||normal
Event|Event|SIMPLE_SEGMENT|3913,3917|false|false|false|||Labs
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3913,3917|false|false|false|C0587081|Laboratory test finding|Labs
Event|Event|SIMPLE_SEGMENT|3919,3927|false|false|false|||Reviewed
Event|Event|SIMPLE_SEGMENT|3936,3939|false|false|false|||see
Procedure|Health Care Activity|SIMPLE_SEGMENT|3971,3976|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMIT
Event|Event|SIMPLE_SEGMENT|3977,3981|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3977,3981|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3996,4001|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3996,4001|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3996,4001|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|4002,4005|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|4013,4016|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4013,4016|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4013,4016|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4023,4026|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4023,4026|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|4023,4026|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4023,4026|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4032,4035|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4032,4035|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|4043,4046|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|4043,4046|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4043,4046|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4043,4046|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4043,4046|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|4050,4053|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4050,4053|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|4050,4053|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|4050,4053|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|4050,4053|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4050,4053|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4060,4064|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4081,4084|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4101,4106|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4101,4106|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4101,4106|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4119,4125|false|false|false|C0024202|Lymph|Lymphs
Drug|Antibiotic|SIMPLE_SEGMENT|4132,4137|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4132,4137|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|SIMPLE_SEGMENT|4132,4137|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4143,4146|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Finding|Gene or Genome|SIMPLE_SEGMENT|4143,4146|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4172,4177|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4172,4177|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4172,4177|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4178,4181|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4198,4203|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4198,4203|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4198,4203|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|4198,4211|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4198,4211|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4198,4211|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4204,4211|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|4204,4211|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4204,4211|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|4204,4211|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4204,4211|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4204,4211|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4253,4257|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4253,4257|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4253,4257|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4282,4287|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4282,4287|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4282,4287|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4288,4291|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4288,4291|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|4288,4291|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|4288,4291|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|4288,4291|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|4288,4291|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|4288,4291|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4288,4291|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4295,4298|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4295,4298|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4295,4298|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4295,4298|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|4295,4298|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|4295,4298|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|4295,4298|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4303,4310|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|SIMPLE_SEGMENT|4303,4310|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4340,4345|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4340,4345|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4340,4345|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4340,4353|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4346,4353|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4346,4353|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4346,4353|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4346,4353|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|4346,4353|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|4346,4353|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|4346,4353|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4346,4353|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4388,4393|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4388,4393|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4388,4393|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4388,4401|false|false|false|C0853248|Blood albumin|BLOOD Albumin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4394,4401|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4394,4401|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4394,4401|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Event|Event|SIMPLE_SEGMENT|4394,4401|false|false|false|||Albumin
Finding|Gene or Genome|SIMPLE_SEGMENT|4394,4401|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Finding|Physiologic Function|SIMPLE_SEGMENT|4394,4401|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4394,4401|false|false|false|C0201838|Albumin measurement|Albumin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4419,4424|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4419,4424|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4419,4424|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4419,4432|false|false|false|C3824990|lactate in blood (lab test)|BLOOD Lactate
Drug|Organic Chemical|SIMPLE_SEGMENT|4425,4432|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4425,4432|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Event|Event|SIMPLE_SEGMENT|4425,4432|false|false|false|||Lactate
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4425,4432|false|false|false|C0202115|Lactic acid measurement|Lactate
Finding|Body Substance|SIMPLE_SEGMENT|4438,4447|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|4438,4447|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|4438,4447|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|4438,4447|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|SIMPLE_SEGMENT|4449,4453|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4449,4453|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4468,4473|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4468,4473|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4468,4473|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|4474,4477|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|4484,4487|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4484,4487|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4484,4487|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4494,4497|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4494,4497|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|4494,4497|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4494,4497|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4503,4506|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4503,4506|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|4514,4517|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|4514,4517|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4514,4517|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4514,4517|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4514,4517|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|4521,4524|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4521,4524|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|4521,4524|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|4521,4524|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|4521,4524|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4521,4524|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4531,4535|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4552,4555|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4572,4577|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4572,4577|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4572,4577|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|4572,4585|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4572,4585|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4572,4585|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4578,4585|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|4578,4585|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4578,4585|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|4578,4585|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4578,4585|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4578,4585|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4628,4632|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4628,4632|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4628,4632|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4657,4662|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4657,4662|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4657,4662|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4663,4666|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4663,4666|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|4663,4666|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|4663,4666|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|4663,4666|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|4663,4666|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|4663,4666|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4663,4666|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4670,4673|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4670,4673|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4670,4673|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4670,4673|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|4670,4673|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|4670,4673|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|4670,4673|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4681,4684|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Drug|Enzyme|SIMPLE_SEGMENT|4681,4684|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Event|Event|SIMPLE_SEGMENT|4681,4684|false|false|false|||LDH
Finding|Finding|SIMPLE_SEGMENT|4681,4684|false|false|false|C0851148|Lifetime Drinking History|LDH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4681,4684|false|false|false|C0202113|Lactate dehydrogenase measurement|LDH
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4691,4698|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|SIMPLE_SEGMENT|4691,4698|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4729,4734|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4729,4734|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4729,4734|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4729,4742|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4735,4742|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4735,4742|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4735,4742|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4735,4742|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|4735,4742|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|4735,4742|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|4735,4742|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4735,4742|false|false|false|C0201925|Calcium measurement|Calcium
Event|Event|SIMPLE_SEGMENT|4764,4771|false|false|false|||IMAGING
Finding|Finding|SIMPLE_SEGMENT|4764,4771|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4764,4771|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Finding|Idea or Concept|SIMPLE_SEGMENT|4777,4782|false|false|false|C1546485|Diagnosis Type - Final|Final
Finding|Intellectual Product|SIMPLE_SEGMENT|4777,4789|false|false|false|C0460114|Final report|Final Report
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4783,4789|false|false|false|C4255046||Report
Event|Event|SIMPLE_SEGMENT|4783,4789|false|false|false|||Report
Finding|Intellectual Product|SIMPLE_SEGMENT|4783,4789|false|false|false|C0684224|Report (document)|Report
Procedure|Health Care Activity|SIMPLE_SEGMENT|4783,4789|false|false|false|C0700287|Reporting|Report
Event|Event|SIMPLE_SEGMENT|4791,4798|false|false|false|||HISTORY
Finding|Conceptual Entity|SIMPLE_SEGMENT|4791,4798|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|HISTORY
Finding|Finding|SIMPLE_SEGMENT|4791,4798|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|HISTORY
Finding|Functional Concept|SIMPLE_SEGMENT|4791,4798|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|HISTORY
Finding|Finding|SIMPLE_SEGMENT|4801,4804|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Finding|Idea or Concept|SIMPLE_SEGMENT|4801,4804|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Finding|Finding|SIMPLE_SEGMENT|4801,4814|false|false|false|C2585997|New diagnosis (finding)|New diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4801,4814|false|false|false|C1882082|New Diagnosis Procedure|New diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4805,4814|false|false|false|C0945731||diagnosis
Event|Event|SIMPLE_SEGMENT|4805,4814|false|false|false|||diagnosis
Finding|Classification|SIMPLE_SEGMENT|4805,4814|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|4805,4814|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4805,4814|false|false|false|C0011900|Diagnosis|diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|4818,4828|false|false|false|C0036525;C1522484|Metastatic to;metastatic qualifier|metastatic
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4818,4835|false|true|false|C0027627;C0346957;C2939419|Disseminated Malignant Neoplasm;Metastatic malignant neoplasm;Neoplasm Metastasis|metastatic cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4829,4835|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|SIMPLE_SEGMENT|4829,4835|false|false|false|||cancer
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4841,4848|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Immunologic Factor|SIMPLE_SEGMENT|4841,4848|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4841,4848|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Event|Event|SIMPLE_SEGMENT|4841,4848|false|false|false|||unknown
Finding|Finding|SIMPLE_SEGMENT|4841,4848|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Functional Concept|SIMPLE_SEGMENT|4841,4848|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Idea or Concept|SIMPLE_SEGMENT|4841,4848|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Intellectual Product|SIMPLE_SEGMENT|4841,4848|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Event|Event|SIMPLE_SEGMENT|4860,4866|false|false|false|||Assess
Event|Event|SIMPLE_SEGMENT|4871,4877|false|false|false|||extent
Event|Event|SIMPLE_SEGMENT|4881,4888|false|false|false|||lesions
Finding|Finding|SIMPLE_SEGMENT|4881,4888|false|false|false|C0221198|Lesion|lesions
Event|Activity|SIMPLE_SEGMENT|4893,4903|false|false|false|C1707455|Comparison|COMPARISON
Event|Event|SIMPLE_SEGMENT|4893,4903|false|false|false|||COMPARISON
Event|Event|SIMPLE_SEGMENT|4906,4908|false|false|false|||CT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4906,4916|false|false|false|C1644645||CT abdomen
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4906,4916|false|false|false|C0412620|CT of abdomen|CT abdomen
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4906,4927|false|false|false|C1715387||CT abdomen and pelvis
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4909,4916|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4909,4916|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Event|Event|SIMPLE_SEGMENT|4909,4916|false|false|false|||abdomen
Finding|Finding|SIMPLE_SEGMENT|4909,4916|false|false|false|C0941288|Abdomen problem|abdomen
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4909,4920|false|false|false|C0000726|Abdomen|abdomen and
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4909,4927|false|false|false|C1508499|Abdominopelvic structure|abdomen and pelvis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4921,4927|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4921,4927|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4921,4927|false|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Finding|Finding|SIMPLE_SEGMENT|4921,4927|false|false|false|C0812455|Pelvis problem|pelvis
Event|Event|SIMPLE_SEGMENT|4928,4933|false|false|false|||dated
Finding|Functional Concept|SIMPLE_SEGMENT|4941,4950|false|false|false|C0449851|Techniques|TECHNIQUE
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4953,4969|false|false|false|C3179130|Multidetector Computed Tomography|Multidetector CT
Event|Event|SIMPLE_SEGMENT|4967,4969|false|false|false|||CT
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4977,4982|false|false|false|C0460005|Trunk structure|torso
Event|Event|SIMPLE_SEGMENT|5003,5014|false|false|false|||intravenous
Finding|Functional Concept|SIMPLE_SEGMENT|5003,5014|false|false|false|C1522726|Intravenous Route of Administration|intravenous
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5019,5023|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5019,5023|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|5019,5023|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|5019,5023|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|5024,5032|false|false|false|C0009924|Contrast Media|contrast
Event|Event|SIMPLE_SEGMENT|5024,5032|false|false|false|||contrast
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5047,5055|false|false|false|C0935598|Sagittal plane|sagittal
Event|Event|SIMPLE_SEGMENT|5057,5069|false|false|false|||reformations
Event|Event|SIMPLE_SEGMENT|5075,5083|false|false|false|||provided
Event|Event|SIMPLE_SEGMENT|5086,5092|false|false|false|||Images
Event|Event|SIMPLE_SEGMENT|5111,5119|false|false|false|||degraded
Finding|Body Substance|SIMPLE_SEGMENT|5132,5139|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|5132,5139|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|5132,5139|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|5142,5146|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5142,5146|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Finding|Intellectual Product|SIMPLE_SEGMENT|5142,5146|false|false|false|C1551342|Document Body|body
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5142,5154|false|false|false|C1318474|Assessment of body build|body habitus
Event|Event|SIMPLE_SEGMENT|5147,5154|false|false|false|||habitus
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5159,5167|false|false|false|C2926606||FINDINGS
Event|Event|SIMPLE_SEGMENT|5159,5167|false|false|false|||FINDINGS
Finding|Functional Concept|SIMPLE_SEGMENT|5159,5167|false|false|false|C2607943|findings aspects|FINDINGS
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5170,5175|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|CHEST
Finding|Finding|SIMPLE_SEGMENT|5170,5175|false|false|false|C0741025|Chest problem|CHEST
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5201,5210|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5201,5210|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|5201,5210|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Finding|SIMPLE_SEGMENT|5201,5218|false|false|false|C0748164|Multiple Pulmonary Nodules|pulmonary nodules
Event|Event|SIMPLE_SEGMENT|5211,5218|false|false|false|||nodules
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5241,5245|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|SIMPLE_SEGMENT|5241,5245|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Event|Event|SIMPLE_SEGMENT|5247,5259|false|false|false|||predilection
Finding|Functional Concept|SIMPLE_SEGMENT|5281,5285|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5281,5296|false|false|false|C1261076|Structure of left upper lobe of lung|left upper lobe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5286,5296|false|false|false|C0225756|Structure of upper lobe of lung|upper lobe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5292,5296|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|SIMPLE_SEGMENT|5292,5296|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Finding|Functional Concept|SIMPLE_SEGMENT|5347,5355|false|false|false|C0004793;C0162326;C0162327;C1519249;C1547787;C3853789|Base Sequence;DNA Sequence;RNA Sequence;Sequence;Sequence - ParameterizedDataType;Sequence - TransmissionRelationshipTypeCode|sequence
Finding|Intellectual Product|SIMPLE_SEGMENT|5347,5355|false|false|false|C0004793;C0162326;C0162327;C1519249;C1547787;C3853789|Base Sequence;DNA Sequence;RNA Sequence;Sequence;Sequence - ParameterizedDataType;Sequence - TransmissionRelationshipTypeCode|sequence
Finding|Nucleotide Sequence|SIMPLE_SEGMENT|5347,5355|false|false|false|C0004793;C0162326;C0162327;C1519249;C1547787;C3853789|Base Sequence;DNA Sequence;RNA Sequence;Sequence;Sequence - ParameterizedDataType;Sequence - TransmissionRelationshipTypeCode|sequence
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5358,5363|false|false|false|C1846009|Intrauterine growth restriction, metaphyseal dysplasia, adrenal hypoplasia congenita, and genital anomaly syndrome|image
Event|Event|SIMPLE_SEGMENT|5358,5363|false|false|false|||image
Finding|Intellectual Product|SIMPLE_SEGMENT|5358,5363|false|false|false|C1696103;C1704254;C1704922;C3542466|Image;Image (foundation metadata concept);Medical Image;image - dosage form|image
Event|Event|SIMPLE_SEGMENT|5369,5382|false|false|false|||Calcification
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5369,5382|false|false|false|C0006660;C0006663;C1533591|Calcification;Calcinosis;Physiologic calcification|Calcification
Finding|Pathologic Function|SIMPLE_SEGMENT|5369,5382|false|false|false|C0006660;C0006663;C1533591|Calcification;Calcinosis;Physiologic calcification|Calcification
Event|Event|SIMPLE_SEGMENT|5387,5392|false|false|false|||noted
Finding|Functional Concept|SIMPLE_SEGMENT|5405,5410|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5405,5425|false|false|false|C0225782|Structure of right pleural cavity|right pleural cavity
Anatomy|Tissue|SIMPLE_SEGMENT|5411,5418|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5411,5418|false|false|false|C0032226|Pleural Diseases|pleural
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5411,5425|false|false|false|C0178802|Pleural cavity|pleural cavity
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5419,5425|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|5419,5425|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5419,5425|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Finding|Functional Concept|SIMPLE_SEGMENT|5427,5435|false|false|false|C0004793;C0162326;C0162327;C1519249;C1547787;C3853789|Base Sequence;DNA Sequence;RNA Sequence;Sequence;Sequence - ParameterizedDataType;Sequence - TransmissionRelationshipTypeCode|sequence
Finding|Intellectual Product|SIMPLE_SEGMENT|5427,5435|false|false|false|C0004793;C0162326;C0162327;C1519249;C1547787;C3853789|Base Sequence;DNA Sequence;RNA Sequence;Sequence;Sequence - ParameterizedDataType;Sequence - TransmissionRelationshipTypeCode|sequence
Finding|Nucleotide Sequence|SIMPLE_SEGMENT|5427,5435|false|false|false|C0004793;C0162326;C0162327;C1519249;C1547787;C3853789|Base Sequence;DNA Sequence;RNA Sequence;Sequence;Sequence - ParameterizedDataType;Sequence - TransmissionRelationshipTypeCode|sequence
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5438,5443|false|false|false|C1846009|Intrauterine growth restriction, metaphyseal dysplasia, adrenal hypoplasia congenita, and genital anomaly syndrome|image
Event|Event|SIMPLE_SEGMENT|5438,5443|false|false|false|||image
Finding|Intellectual Product|SIMPLE_SEGMENT|5438,5443|false|false|false|C1696103;C1704254;C1704922;C3542466|Image;Image (foundation metadata concept);Medical Image;image - dosage form|image
Finding|Finding|SIMPLE_SEGMENT|5459,5465|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|5459,5465|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Drug|Organic Chemical|SIMPLE_SEGMENT|5466,5473|false|true|false|C0163712|Relate - vinyl resin|related
Event|Event|SIMPLE_SEGMENT|5466,5473|false|false|false|||related
Finding|Finding|SIMPLE_SEGMENT|5466,5473|false|true|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|SIMPLE_SEGMENT|5466,5473|false|true|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Body Substance|SIMPLE_SEGMENT|5481,5488|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|5481,5488|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|5481,5488|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|5491,5498|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|5491,5498|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|5491,5498|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|5491,5498|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|5491,5501|false|false|false|C0262926|Medical History|history of
Event|Event|SIMPLE_SEGMENT|5502,5510|false|false|false|||previous
Finding|Functional Concept|SIMPLE_SEGMENT|5512,5517|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5512,5522|false|false|false|C0225706|Right lung|right lung
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5518,5522|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5518,5522|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5518,5522|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|5518,5522|false|false|false|C0740941|Lung Problem|lung
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5518,5530|false|false|false|C0038903|Pulmonary Surgical Procedures|lung surgery
Event|Event|SIMPLE_SEGMENT|5523,5530|false|false|false|||surgery
Finding|Finding|SIMPLE_SEGMENT|5523,5530|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|5523,5530|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|5523,5530|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5523,5530|false|false|false|C0543467|Operative Surgical Procedures|surgery
Anatomy|Tissue|SIMPLE_SEGMENT|5536,5543|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5536,5543|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Body Substance|SIMPLE_SEGMENT|5536,5552|true|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Finding|SIMPLE_SEGMENT|5536,5552|true|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|5536,5552|true|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Event|Event|SIMPLE_SEGMENT|5544,5552|false|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|5544,5552|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|5544,5552|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|5544,5552|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5558,5570|true|false|false|C0032326|Pneumothorax|pneumothorax
Event|Event|SIMPLE_SEGMENT|5558,5570|false|false|false|||pneumothorax
Finding|Idea or Concept|SIMPLE_SEGMENT|5577,5588|false|false|false|C0750502|Significant|significant
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5589,5600|false|false|false|C0025066|Mediastinum|mediastinal
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5602,5610|false|false|false|C0004454|Axilla|axillary
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5614,5630|true|false|false|C0456973|Hilar lymphadenopathy|hilar adenopathy
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5620,5630|false|false|false|C0497156|Lymphadenopathy|adenopathy
Event|Event|SIMPLE_SEGMENT|5620,5630|false|false|false|||adenopathy
Finding|Sign or Symptom|SIMPLE_SEGMENT|5620,5630|false|false|false|C4282165|Swollen Lymph Node|adenopathy
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5634,5641|false|false|false|C0018787|Heart|Cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|5634,5641|false|false|false|C1314974|Cardiac attachment|Cardiac
Event|Event|SIMPLE_SEGMENT|5651,5657|false|false|false|||normal
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5663,5674|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5663,5674|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5663,5683|true|false|false|C0031039|Pericardial effusion|pericardial effusion
Finding|Body Substance|SIMPLE_SEGMENT|5663,5683|true|false|false|C1253937|Pericardial effusion body substance|pericardial effusion
Event|Event|SIMPLE_SEGMENT|5675,5683|false|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|5675,5683|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|5675,5683|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|5675,5683|true|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5687,5694|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5687,5694|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|SIMPLE_SEGMENT|5687,5694|false|false|false|||ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|5687,5694|false|false|false|C0941288|Abdomen problem|ABDOMEN
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5702,5707|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5702,5707|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5702,5707|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|SIMPLE_SEGMENT|5702,5707|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5702,5707|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|SIMPLE_SEGMENT|5702,5707|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|SIMPLE_SEGMENT|5702,5707|false|false|false|||liver
Finding|Finding|SIMPLE_SEGMENT|5702,5707|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|SIMPLE_SEGMENT|5702,5707|false|false|false|C0872387|Procedures on liver|liver
Event|Event|SIMPLE_SEGMENT|5711,5719|false|false|false|||enlarged
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5711,5719|false|false|false|C1293134|Enlargement procedure|enlarged
Event|Event|SIMPLE_SEGMENT|5750,5757|false|false|false|||density
Event|Event|SIMPLE_SEGMENT|5759,5766|false|false|false|||lesions
Finding|Finding|SIMPLE_SEGMENT|5759,5766|false|false|false|C0221198|Lesion|lesions
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5783,5788|false|false|false|C0796494|lobe|lobes
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5796,5801|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5796,5801|true|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5796,5801|true|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|SIMPLE_SEGMENT|5796,5801|true|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5796,5801|true|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|SIMPLE_SEGMENT|5796,5801|true|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|SIMPLE_SEGMENT|5796,5801|false|false|false|||liver
Finding|Finding|SIMPLE_SEGMENT|5796,5801|true|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|SIMPLE_SEGMENT|5796,5801|true|false|false|C0872387|Procedures on liver|liver
Event|Event|SIMPLE_SEGMENT|5812,5821|false|false|false|||replacing
Finding|Intellectual Product|SIMPLE_SEGMENT|5827,5831|false|false|false|C0814230|veterans alcoholism screening test (VAST)|vast
Event|Event|SIMPLE_SEGMENT|5832,5840|false|false|false|||majority
Finding|Social Behavior|SIMPLE_SEGMENT|5832,5840|false|false|false|C0680220|majority|majority
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5848,5855|false|false|false|C0205054|Hepatic|hepatic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5848,5866|false|false|false|C0736268|Liver parenchyma|hepatic parenchyma
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5856,5866|false|false|false|C0933845|Parenchyma|parenchyma
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5873,5879|false|false|false|C0205054|Hepatic|portal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5873,5884|false|false|false|C0032718;C1305775;C4266644|Abdomen>Portal vein;Portal vein structure|portal vein
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5880,5884|false|false|false|C0042449|Veins|vein
Event|Event|SIMPLE_SEGMENT|5889,5895|false|false|false|||patent
Finding|Intellectual Product|SIMPLE_SEGMENT|5889,5895|false|false|false|C0030650|Legal patent|patent
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5923,5927|false|false|false|C0687028;C1550227|Duct (organ) structure;canal [body parts]|duct
Event|Event|SIMPLE_SEGMENT|5928,5938|false|false|false|||dilatation
Finding|Finding|SIMPLE_SEGMENT|5928,5938|true|false|false|C0012359;C0700124|Dilated;Pathological Dilatation|dilatation
Finding|Pathologic Function|SIMPLE_SEGMENT|5928,5938|true|false|false|C0012359;C0700124|Dilated;Pathological Dilatation|dilatation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5928,5938|true|false|false|C1322279|Dilate procedure|dilatation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5946,5957|false|false|false|C0016976;C1524055;C4071903|Abdomen>Gallbladder;Gallbladder;Gallbladder (MMHCC)|gallbladder
Anatomy|Tissue|SIMPLE_SEGMENT|5946,5957|false|false|false|C0016976;C1524055;C4071903|Abdomen>Gallbladder;Gallbladder;Gallbladder (MMHCC)|gallbladder
Event|Event|SIMPLE_SEGMENT|5946,5957|false|false|false|||gallbladder
Procedure|Health Care Activity|SIMPLE_SEGMENT|5946,5957|false|false|false|C2032932|examination of gallbladder|gallbladder
Event|Event|SIMPLE_SEGMENT|5961,5973|false|false|false|||unremarkable
Event|Event|SIMPLE_SEGMENT|5993,5999|false|false|false|||amount
Finding|Intellectual Product|SIMPLE_SEGMENT|5993,5999|false|false|false|C1561574|Amount class - Amount|amount
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6003,6010|false|false|false|C0003962|Ascites|ascites
Event|Event|SIMPLE_SEGMENT|6003,6010|false|false|false|||ascites
Finding|Pathologic Function|SIMPLE_SEGMENT|6003,6010|false|false|false|C5441966|Peritoneal Effusion|ascites
Event|Event|SIMPLE_SEGMENT|6012,6020|false|false|false|||adjacent
Finding|Functional Concept|SIMPLE_SEGMENT|6028,6033|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6028,6051|false|false|false|C0227481|Right lobe of liver|right lobe of the liver
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6034,6038|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|SIMPLE_SEGMENT|6034,6038|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6046,6051|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6046,6051|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6046,6051|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|SIMPLE_SEGMENT|6046,6051|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6046,6051|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|SIMPLE_SEGMENT|6046,6051|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|SIMPLE_SEGMENT|6046,6051|false|false|false|||liver
Finding|Finding|SIMPLE_SEGMENT|6046,6051|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|SIMPLE_SEGMENT|6046,6051|false|false|false|C0872387|Procedures on liver|liver
Finding|Functional Concept|SIMPLE_SEGMENT|6063,6068|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6063,6075|false|false|false|C0227613|Right kidney|right kidney
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6069,6075|false|false|false|C0022646;C0227665|Both kidneys;Kidney|kidney
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6069,6075|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|kidney
Event|Event|SIMPLE_SEGMENT|6069,6075|false|false|false|||kidney
Finding|Sign or Symptom|SIMPLE_SEGMENT|6069,6075|false|false|false|C0812426|Kidney problem|kidney
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6069,6075|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6069,6075|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Event|Event|SIMPLE_SEGMENT|6086,6096|false|false|false|||compressed
Event|Event|SIMPLE_SEGMENT|6120,6128|false|false|false|||enlarged
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6120,6128|false|false|false|C1293134|Enlargement procedure|enlarged
Finding|Finding|SIMPLE_SEGMENT|6120,6134|false|false|false|C0019209|Hepatomegaly|enlarged liver
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6129,6134|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6129,6134|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6129,6134|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|SIMPLE_SEGMENT|6129,6134|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6129,6134|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|SIMPLE_SEGMENT|6129,6134|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|SIMPLE_SEGMENT|6129,6134|false|false|false|||liver
Finding|Finding|SIMPLE_SEGMENT|6129,6134|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|SIMPLE_SEGMENT|6129,6134|false|false|false|C0872387|Procedures on liver|liver
Event|Event|SIMPLE_SEGMENT|6173,6179|false|false|false|||lesion
Finding|Finding|SIMPLE_SEGMENT|6173,6179|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|SIMPLE_SEGMENT|6173,6179|false|false|false|C0221198;C1546698|Lesion|lesion
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6194,6198|false|false|false|C0935623|anatomical pole|pole
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6194,6198|false|false|false|C3811771|DNA Polymerase Epsilon Catalytic Subunit A, Human|pole
Drug|Enzyme|SIMPLE_SEGMENT|6194,6198|false|false|false|C3811771|DNA Polymerase Epsilon Catalytic Subunit A, Human|pole
Finding|Gene or Genome|SIMPLE_SEGMENT|6194,6198|false|false|false|C1418729|POLE gene|pole
Finding|Functional Concept|SIMPLE_SEGMENT|6206,6211|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6206,6218|false|false|false|C0227613|Right kidney|right kidney
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6212,6218|false|false|false|C0022646;C0227665|Both kidneys;Kidney|kidney
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6212,6218|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|kidney
Event|Event|SIMPLE_SEGMENT|6212,6218|false|false|false|||kidney
Finding|Sign or Symptom|SIMPLE_SEGMENT|6212,6218|false|false|false|C0812426|Kidney problem|kidney
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6212,6218|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6212,6218|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Finding|Finding|SIMPLE_SEGMENT|6220,6226|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|6220,6226|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|SIMPLE_SEGMENT|6227,6239|false|false|false|||representing
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|6257,6261|false|false|false|C0010709|Cyst|cyst
Event|Event|SIMPLE_SEGMENT|6257,6261|false|false|false|||cyst
Finding|Body Substance|SIMPLE_SEGMENT|6257,6261|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Finding|Intellectual Product|SIMPLE_SEGMENT|6257,6261|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Finding|Functional Concept|SIMPLE_SEGMENT|6263,6271|false|false|false|C0004793;C0162326;C0162327;C1519249;C1547787;C3853789|Base Sequence;DNA Sequence;RNA Sequence;Sequence;Sequence - ParameterizedDataType;Sequence - TransmissionRelationshipTypeCode|sequence
Finding|Intellectual Product|SIMPLE_SEGMENT|6263,6271|false|false|false|C0004793;C0162326;C0162327;C1519249;C1547787;C3853789|Base Sequence;DNA Sequence;RNA Sequence;Sequence;Sequence - ParameterizedDataType;Sequence - TransmissionRelationshipTypeCode|sequence
Finding|Nucleotide Sequence|SIMPLE_SEGMENT|6263,6271|false|false|false|C0004793;C0162326;C0162327;C1519249;C1547787;C3853789|Base Sequence;DNA Sequence;RNA Sequence;Sequence;Sequence - ParameterizedDataType;Sequence - TransmissionRelationshipTypeCode|sequence
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6274,6279|false|false|false|C1846009|Intrauterine growth restriction, metaphyseal dysplasia, adrenal hypoplasia congenita, and genital anomaly syndrome|image
Event|Event|SIMPLE_SEGMENT|6274,6279|false|false|false|||image
Finding|Intellectual Product|SIMPLE_SEGMENT|6274,6279|false|false|false|C1696103;C1704254;C1704922;C3542466|Image;Image (foundation metadata concept);Medical Image;image - dosage form|image
Finding|Functional Concept|SIMPLE_SEGMENT|6290,6295|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6290,6302|false|false|false|C0227613|Right kidney|right kidney
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6296,6302|false|false|false|C0022646;C0227665|Both kidneys;Kidney|kidney
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6296,6302|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|kidney
Event|Event|SIMPLE_SEGMENT|6296,6302|false|false|false|||kidney
Finding|Sign or Symptom|SIMPLE_SEGMENT|6296,6302|false|false|false|C0812426|Kidney problem|kidney
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6296,6302|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6296,6302|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Event|Event|SIMPLE_SEGMENT|6317,6329|false|false|false|||unremarkable
Finding|Functional Concept|SIMPLE_SEGMENT|6336,6340|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6336,6347|false|false|false|C0227614|Left kidney|left kidney
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6341,6347|false|false|false|C0022646;C0227665|Both kidneys;Kidney|kidney
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6341,6347|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|kidney
Event|Event|SIMPLE_SEGMENT|6341,6347|false|false|false|||kidney
Finding|Sign or Symptom|SIMPLE_SEGMENT|6341,6347|false|false|false|C0812426|Kidney problem|kidney
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6341,6347|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6341,6347|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Event|Event|SIMPLE_SEGMENT|6358,6364|false|false|false|||normal
Event|Event|SIMPLE_SEGMENT|6366,6372|false|false|false|||limits
Finding|Functional Concept|SIMPLE_SEGMENT|6366,6372|false|false|false|C0439801|Limited (extensiveness)|limits
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6379,6387|false|false|false|C0001625|Adrenal Glands|adrenals
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6392,6398|false|false|false|C0037993;C4037984|Abdomen>Spleen;Spleen|spleen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6392,6398|false|false|false|C0153470|Malignant neoplasm of spleen|spleen
Event|Event|SIMPLE_SEGMENT|6392,6398|false|false|false|||spleen
Finding|Finding|SIMPLE_SEGMENT|6392,6398|false|false|false|C0812414|Spleen problem|spleen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6392,6398|false|false|false|C0869677|Procedures on Spleen|spleen
Event|Event|SIMPLE_SEGMENT|6403,6415|false|false|false|||unremarkable
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6422,6430|false|false|false|C0030274;C4037927|Abdomen>Pancreas;Pancreas|pancreas
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6422,6430|false|false|false|C0030286;C0347284|Benign tumor of pancreas;Pancreatic Diseases|pancreas
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6422,6430|false|false|false|C0030286;C0347284|Benign tumor of pancreas;Pancreatic Diseases|pancreas
Drug|Organic Chemical|SIMPLE_SEGMENT|6422,6430|false|false|false|C0771711|pancreas extract|pancreas
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6422,6430|false|false|false|C0771711|pancreas extract|pancreas
Event|Event|SIMPLE_SEGMENT|6422,6430|false|false|false|||pancreas
Finding|Finding|SIMPLE_SEGMENT|6422,6430|false|false|false|C0813176|Pancreas problem|pancreas
Procedure|Health Care Activity|SIMPLE_SEGMENT|6422,6430|false|false|false|C0869826|Procedures on Pancreas|pancreas
Finding|Finding|SIMPLE_SEGMENT|6435,6455|false|false|false|C0442816||within normal limits
Event|Event|SIMPLE_SEGMENT|6449,6455|false|false|false|||limits
Finding|Functional Concept|SIMPLE_SEGMENT|6449,6455|false|false|false|C0439801|Limited (extensiveness)|limits
Finding|Gene or Genome|SIMPLE_SEGMENT|6472,6477|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6472,6483|false|false|false|C0021851|Large Intestine|large bowel
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6478,6483|false|false|false|C0021853|Intestines|bowel
Event|Event|SIMPLE_SEGMENT|6489,6501|false|false|false|||unremarkable
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6507,6522|false|false|false|C0035359|Retroperitoneal Space|retroperitoneal
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6526,6536|false|false|false|C0025474|Mesentery|mesenteric
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6537,6547|true|false|false|C0497156|Lymphadenopathy|adenopathy
Event|Event|SIMPLE_SEGMENT|6537,6547|false|false|false|||adenopathy
Finding|Sign or Symptom|SIMPLE_SEGMENT|6537,6547|true|false|false|C4282165|Swollen Lymph Node|adenopathy
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6554,6560|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|PELVIS
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6554,6560|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|PELVIS
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6554,6560|false|false|false|C0153663|Malignant neoplasm of pelvis|PELVIS
Event|Event|SIMPLE_SEGMENT|6554,6560|false|false|false|||PELVIS
Finding|Finding|SIMPLE_SEGMENT|6554,6560|false|false|false|C0812455|Pelvis problem|PELVIS
Event|Event|SIMPLE_SEGMENT|6568,6574|false|false|false|||images
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6582,6588|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6582,6588|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6582,6588|false|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Finding|Finding|SIMPLE_SEGMENT|6582,6588|false|false|false|C0812455|Pelvis problem|pelvis
Event|Event|SIMPLE_SEGMENT|6607,6615|false|false|false|||degraded
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6616,6625|false|false|false|C0027627|Neoplasm Metastasis|secondary
Event|Event|SIMPLE_SEGMENT|6616,6625|false|false|false|||secondary
Finding|Functional Concept|SIMPLE_SEGMENT|6616,6625|false|false|false|C1522484|metastatic qualifier|secondary
Finding|Body Substance|SIMPLE_SEGMENT|6634,6641|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6634,6641|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6634,6641|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|6644,6648|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6644,6648|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Finding|Intellectual Product|SIMPLE_SEGMENT|6644,6648|false|false|false|C1551342|Document Body|body
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6644,6656|false|false|false|C1318474|Assessment of body build|body habitus
Event|Event|SIMPLE_SEGMENT|6649,6656|false|false|false|||habitus
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6662,6668|false|false|false|C0030797|Pelvis|pelvic
Event|Event|SIMPLE_SEGMENT|6669,6675|false|false|false|||masses
Event|Event|SIMPLE_SEGMENT|6680,6690|false|false|false|||identified
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6698,6705|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6698,6705|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Event|Event|SIMPLE_SEGMENT|6698,6705|false|false|false|||bladder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6698,6705|false|false|false|C0872388|Procedures on bladder|bladder
Event|Event|SIMPLE_SEGMENT|6709,6721|false|false|false|||unremarkable
Finding|Body Substance|SIMPLE_SEGMENT|6728,6735|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6728,6735|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6728,6735|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6739,6745|false|false|false|C5889824||status
Event|Event|SIMPLE_SEGMENT|6739,6745|false|false|false|||status
Finding|Idea or Concept|SIMPLE_SEGMENT|6739,6745|false|false|false|C1546481|What subject filter - Status|status
Finding|Gene or Genome|SIMPLE_SEGMENT|6746,6750|false|false|false|C3469826;C3470073|DESI1 gene;SLC35G1 gene|post
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6752,6778|false|false|false|C1270947;C1270948|Partial hysterectomy;Supracervical hysterectomy|supracervical hysterectomy
Event|Event|SIMPLE_SEGMENT|6766,6778|false|false|false|||hysterectomy
Finding|Finding|SIMPLE_SEGMENT|6766,6778|false|false|false|C1548863|Consent Type - Hysterectomy|hysterectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6766,6778|false|false|false|C0020699|Hysterectomy|hysterectomy
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6784,6790|false|false|false|C0030797|Pelvis|pelvic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6791,6801|true|false|false|C0497156|Lymphadenopathy|adenopathy
Event|Event|SIMPLE_SEGMENT|6791,6801|false|false|false|||adenopathy
Finding|Sign or Symptom|SIMPLE_SEGMENT|6791,6801|true|false|false|C4282165|Swollen Lymph Node|adenopathy
Event|Event|SIMPLE_SEGMENT|6806,6810|false|false|false|||free
Finding|Functional Concept|SIMPLE_SEGMENT|6806,6810|true|false|false|C0332296|Free of (attribute)|free
Finding|Pathologic Function|SIMPLE_SEGMENT|6806,6816|true|false|false|C0013687|effusion|free fluid
Drug|Substance|SIMPLE_SEGMENT|6811,6816|true|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|6811,6816|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|6811,6816|true|false|false|C1546638|Fluid Specimen Code|fluid
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6829,6835|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6829,6835|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6829,6835|false|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Finding|Finding|SIMPLE_SEGMENT|6829,6835|false|false|false|C0812455|Pelvis problem|pelvis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6842,6849|false|false|false|C0262950;C4520924|Bone Tissue, Human;Skeletal bone|OSSEOUS
Anatomy|Tissue|SIMPLE_SEGMENT|6842,6849|false|false|false|C0262950;C4520924|Bone Tissue, Human;Skeletal bone|OSSEOUS
Event|Event|SIMPLE_SEGMENT|6850,6860|false|false|false|||STRUCTURES
Finding|Finding|SIMPLE_SEGMENT|6874,6885|false|false|false|C0332516|Symmetrical|symmetrical
Event|Event|SIMPLE_SEGMENT|6886,6895|false|false|false|||sclerosis
Finding|Pathologic Function|SIMPLE_SEGMENT|6886,6895|false|false|false|C0036429|Sclerosis|sclerosis
Event|Event|SIMPLE_SEGMENT|6899,6909|false|false|false|||identified
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6917,6922|false|false|false|C0020889|Bone structure of ilium|iliac
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6937,6947|false|false|false|C0555898|sacroiliac|sacroiliac
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6937,6954|false|false|false|C0036036|Sacroiliac joint structure|sacroiliac joints
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6948,6954|false|false|false|C0022417;C0392905|Articular system;Joints|joints
Anatomy|Body System|SIMPLE_SEGMENT|6948,6954|false|false|false|C0022417;C0392905|Articular system;Joints|joints
Event|Event|SIMPLE_SEGMENT|6956,6966|false|false|false|||consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|6956,6966|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|6956,6971|false|false|false|C0332290|Consistent with|consistent with
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6972,6980|false|false|false|C0029400|Osteitis|osteitis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6972,6991|false|false|false|C0152263|Osteitis condensans|osteitis condensans
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6972,6996|false|false|false|C0343261|Osteitis condensans ilii|osteitis condensans ilii
Event|Event|SIMPLE_SEGMENT|6992,6996|false|false|false|||ilii
Finding|Finding|SIMPLE_SEGMENT|7009,7015|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|7009,7015|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Functional Concept|SIMPLE_SEGMENT|7016,7028|false|false|false|C0011164;C1880269|Abnormal degeneration;biologic degeneration|degenerative
Finding|Pathologic Function|SIMPLE_SEGMENT|7016,7028|false|false|false|C0011164;C1880269|Abnormal degeneration;biologic degeneration|degenerative
Finding|Pathologic Function|SIMPLE_SEGMENT|7016,7035|false|false|false|C0011164|Abnormal degeneration|degenerative change
Event|Event|SIMPLE_SEGMENT|7029,7035|false|false|false|||change
Finding|Functional Concept|SIMPLE_SEGMENT|7029,7035|false|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7029,7035|false|false|false|C4319952|Change - procedure|change
Finding|Functional Concept|SIMPLE_SEGMENT|7047,7052|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7047,7056|false|false|false|C0524470|Right hip region structure|right hip
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|7047,7062|false|false|false|C1285116|Right hip joint structure|right hip joint
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7053,7056|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7053,7056|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7053,7056|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7053,7056|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|SIMPLE_SEGMENT|7053,7056|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7053,7056|false|false|false|C1292890|Procedure on hip|hip
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|7053,7062|false|false|false|C0019558|Hip Joint|hip joint
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|7057,7062|false|false|false|C0022417;C0392905;C1269611|Articular system;Joints|joint
Anatomy|Body System|SIMPLE_SEGMENT|7057,7062|false|false|false|C0022417;C0392905;C1269611|Articular system;Joints|joint
Finding|Finding|SIMPLE_SEGMENT|7057,7062|false|false|false|C0575044|Joint problem|joint
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|7069,7074|false|false|false|C0022417;C0392905;C1269611|Articular system;Joints|joint
Anatomy|Body System|SIMPLE_SEGMENT|7069,7074|false|false|false|C0022417;C0392905;C1269611|Articular system;Joints|joint
Finding|Finding|SIMPLE_SEGMENT|7069,7074|false|false|false|C0575044|Joint problem|joint
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|7069,7080|false|false|false|C0224497|Articular space|joint space
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|7075,7080|false|false|false|C0282173|Space (Astronomy)|space
Event|Event|SIMPLE_SEGMENT|7081,7085|false|false|false|||loss
Finding|Finding|SIMPLE_SEGMENT|7081,7085|false|false|false|C5890125|Loss (adaptation)|loss
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7090,7100|false|false|false|C0015302;C1956089|External hyperostosis;Osteophyte|osteophyte
Finding|Pathologic Function|SIMPLE_SEGMENT|7090,7110|false|false|false|C5442360|Osteophyte formation|osteophyte formation
Event|Event|SIMPLE_SEGMENT|7101,7110|false|false|false|||formation
Finding|Functional Concept|SIMPLE_SEGMENT|7101,7110|false|false|false|C1522492|Formation|formation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|7101,7110|false|false|false|C0220781|Anabolism|formation
Event|Event|SIMPLE_SEGMENT|7116,7127|false|false|false|||destructive
Finding|Individual Behavior|SIMPLE_SEGMENT|7116,7127|true|false|false|C0233520|Destructive behavior|destructive
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7129,7136|false|false|false|C0262950;C4520924|Bone Tissue, Human;Skeletal bone|osseous
Anatomy|Tissue|SIMPLE_SEGMENT|7129,7136|false|false|false|C0262950;C4520924|Bone Tissue, Human;Skeletal bone|osseous
Event|Event|SIMPLE_SEGMENT|7137,7144|false|false|false|||lesions
Finding|Finding|SIMPLE_SEGMENT|7137,7144|false|false|false|C0221198|Lesion|lesions
Event|Event|SIMPLE_SEGMENT|7152,7162|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|7152,7162|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|7152,7162|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7174,7183|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7174,7183|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|7174,7183|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7188,7195|false|false|false|C0205054|Hepatic|hepatic
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7188,7206|false|false|false|C0494165|Metastatic malignant neoplasm to liver|hepatic metastases
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7196,7206|false|false|false|C0027627;C2939419|Metastatic malignant neoplasm;Neoplasm Metastasis|metastases
Event|Event|SIMPLE_SEGMENT|7196,7206|false|false|false|||metastases
Finding|Finding|SIMPLE_SEGMENT|7196,7206|false|false|false|C1513183|Metastatic Lesion|metastases
Event|Event|SIMPLE_SEGMENT|7230,7236|false|false|false|||lesion
Finding|Finding|SIMPLE_SEGMENT|7230,7236|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|SIMPLE_SEGMENT|7230,7236|false|false|false|C0221198;C1546698|Lesion|lesion
Event|Event|SIMPLE_SEGMENT|7238,7248|false|false|false|||identified
Finding|Intellectual Product|SIMPLE_SEGMENT|7256,7261|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|7262,7270|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7262,7277|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|7262,7277|false|false|false|C0489547|Hospital course|Hospital Course
Event|Event|SIMPLE_SEGMENT|7306,7315|false|false|false|||diagnosed
Finding|Functional Concept|SIMPLE_SEGMENT|7316,7326|false|true|false|C0036525;C1522484|Metastatic to;metastatic qualifier|metastatic
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7316,7333|false|true|false|C0027627;C0346957;C2939419|Disseminated Malignant Neoplasm;Metastatic malignant neoplasm;Neoplasm Metastasis|metastatic cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7327,7333|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|SIMPLE_SEGMENT|7327,7333|false|false|false|||cancer
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7337,7344|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Immunologic Factor|SIMPLE_SEGMENT|7337,7344|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7337,7344|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Event|Event|SIMPLE_SEGMENT|7337,7344|false|false|false|||unknown
Finding|Finding|SIMPLE_SEGMENT|7337,7344|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Functional Concept|SIMPLE_SEGMENT|7337,7344|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Idea or Concept|SIMPLE_SEGMENT|7337,7344|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Intellectual Product|SIMPLE_SEGMENT|7337,7344|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Event|Event|SIMPLE_SEGMENT|7354,7364|false|false|false|||presenting
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7370,7376|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|7370,7376|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|7370,7376|false|false|false|C0027497|Nausea|nausea
Event|Event|SIMPLE_SEGMENT|7378,7386|false|false|false|||vomiting
Finding|Sign or Symptom|SIMPLE_SEGMENT|7378,7386|false|false|false|C0042963|Vomiting|vomiting
Event|Event|SIMPLE_SEGMENT|7392,7397|false|false|false|||fever
Finding|Finding|SIMPLE_SEGMENT|7392,7397|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|7392,7397|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Idea or Concept|SIMPLE_SEGMENT|7409,7412|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|7409,7412|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|7416,7425|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|7416,7425|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|7433,7438|false|false|false|||Fever
Finding|Finding|SIMPLE_SEGMENT|7433,7438|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|7433,7438|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7439,7451|false|false|false|C0023518|Leukocytosis|leukocytosis
Event|Event|SIMPLE_SEGMENT|7439,7451|false|false|false|||leukocytosis
Finding|Finding|SIMPLE_SEGMENT|7439,7451|false|false|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Finding|Body Substance|SIMPLE_SEGMENT|7453,7460|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7453,7460|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7453,7460|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|7461,7470|false|false|false|||presented
Event|Event|SIMPLE_SEGMENT|7476,7481|false|false|false|||fever
Finding|Finding|SIMPLE_SEGMENT|7476,7481|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|7476,7481|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7487,7499|false|false|false|C0023518|Leukocytosis|leukocytosis
Event|Event|SIMPLE_SEGMENT|7487,7499|false|false|false|||leukocytosis
Finding|Finding|SIMPLE_SEGMENT|7487,7499|false|false|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Event|Event|SIMPLE_SEGMENT|7521,7531|false|false|false|||concerning
Event|Event|SIMPLE_SEGMENT|7536,7540|false|false|false|||post
Finding|Gene or Genome|SIMPLE_SEGMENT|7536,7540|false|false|false|C3469826;C3470073|DESI1 gene;SLC35G1 gene|post
Finding|Functional Concept|SIMPLE_SEGMENT|7542,7553|false|false|false|C0549186|Obstructed|obstructive
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|7554,7557|false|false|false|C0600500|Peptide Nucleic Acids|PNA
Event|Event|SIMPLE_SEGMENT|7554,7557|false|false|false|||PNA
Finding|Body Substance|SIMPLE_SEGMENT|7559,7566|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7559,7566|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7559,7566|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|7571,7578|false|false|false|||treated
Drug|Antibiotic|SIMPLE_SEGMENT|7589,7597|false|false|false|C0055003|cefepime|cefepime
Drug|Organic Chemical|SIMPLE_SEGMENT|7589,7597|false|false|false|C0055003|cefepime|cefepime
Event|Event|SIMPLE_SEGMENT|7598,7605|false|false|false|||azithro
Finding|Idea or Concept|SIMPLE_SEGMENT|7613,7616|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|7613,7616|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|7637,7639|false|false|false|||CT
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7640,7645|false|false|false|C0460005|Trunk structure|torso
Event|Event|SIMPLE_SEGMENT|7650,7660|false|false|false|||concerning
Finding|Idea or Concept|SIMPLE_SEGMENT|7666,7673|false|false|false|C0549178|Continuous|ongoing
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7674,7684|false|false|false|C0006826;C1306459|Malignant Neoplasms;Primary malignant neoplasm|malignancy
Event|Event|SIMPLE_SEGMENT|7674,7684|false|false|false|||malignancy
Event|Event|SIMPLE_SEGMENT|7693,7701|false|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|7693,7701|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|7693,7704|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7705,7718|true|false|false|C0677930|Primary Neoplasm|primary tumor
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7713,7718|true|false|false|C0027651|Neoplasms|tumor
Event|Event|SIMPLE_SEGMENT|7713,7718|false|false|false|||tumor
Finding|Finding|SIMPLE_SEGMENT|7713,7718|true|false|false|C1578706;C3273930|Tumor Mass|tumor
Finding|Intellectual Product|SIMPLE_SEGMENT|7713,7718|true|false|false|C1578706;C3273930|Tumor Mass|tumor
Event|Event|SIMPLE_SEGMENT|7734,7741|false|false|false|||concern
Finding|Idea or Concept|SIMPLE_SEGMENT|7734,7741|true|false|false|C2699424|Concern|concern
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7748,7757|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|SIMPLE_SEGMENT|7748,7757|false|false|false|||pneumonia
Event|Event|SIMPLE_SEGMENT|7782,7789|false|false|false|||stopped
Finding|Body Substance|SIMPLE_SEGMENT|7799,7806|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7799,7806|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7799,7806|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|7807,7811|false|false|false|||felt
Event|Event|SIMPLE_SEGMENT|7812,7816|false|false|false|||weak
Finding|Intellectual Product|SIMPLE_SEGMENT|7812,7816|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|weak
Finding|Sign or Symptom|SIMPLE_SEGMENT|7812,7816|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|weak
Event|Event|SIMPLE_SEGMENT|7821,7827|false|false|false|||unable
Finding|Finding|SIMPLE_SEGMENT|7821,7827|false|false|false|C1299582|Unable|unable
Event|Event|SIMPLE_SEGMENT|7834,7838|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|7834,7838|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|7834,7838|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|7834,7838|false|false|false|C1553498|home health encounter|home
Finding|Finding|SIMPLE_SEGMENT|7854,7859|false|false|false|C0439044|Living Alone|alone
Event|Event|SIMPLE_SEGMENT|7871,7879|false|false|false|||screened
Finding|Finding|SIMPLE_SEGMENT|7883,7891|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Finding|Functional Concept|SIMPLE_SEGMENT|7883,7891|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|7883,7891|false|false|false|C0031809|Physical Examination|physical
Finding|Intellectual Product|SIMPLE_SEGMENT|7883,7899|false|false|false|C1547999|Diagnostic Service Section ID - Physical Therapy|physical therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7883,7899|false|false|false|C0949766|Physical therapy|physical therapy
Event|Event|SIMPLE_SEGMENT|7892,7899|false|false|false|||therapy
Finding|Finding|SIMPLE_SEGMENT|7892,7899|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|SIMPLE_SEGMENT|7892,7899|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7892,7899|false|false|false|C0087111|Therapeutic procedure|therapy
Event|Event|SIMPLE_SEGMENT|7904,7914|false|false|false|||discharged
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7919,7924|false|false|false|C0034991|Rehabilitation therapy|rehab
Event|Event|SIMPLE_SEGMENT|7925,7933|false|false|false|||facility
Finding|Intellectual Product|SIMPLE_SEGMENT|7925,7933|false|false|false|C4695111|ADMIN.FACILITY|facility
Finding|Functional Concept|SIMPLE_SEGMENT|7940,7947|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|Failure
Finding|Idea or Concept|SIMPLE_SEGMENT|7940,7947|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|Failure
Finding|Individual Behavior|SIMPLE_SEGMENT|7940,7947|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|Failure
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7940,7957|false|false|false|C0015544;C2315100|Failure to Thrive;Pediatric failure to thrive|Failure to thrive
Drug|Organic Chemical|SIMPLE_SEGMENT|7951,7957|false|false|false|C2938208|Thrive|thrive
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7951,7957|false|false|false|C2938208|Thrive|thrive
Event|Event|SIMPLE_SEGMENT|7951,7957|false|false|false|||thrive
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7951,7957|false|false|false|C4760774|Transnasal humidified rapid-insufflation ventilatory exchange|thrive
Finding|Body Substance|SIMPLE_SEGMENT|7959,7966|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7959,7966|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7959,7966|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|7967,7975|false|false|false|||presents
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7992,7998|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|7992,7998|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|7992,7998|false|false|false|C0027497|Nausea|nausea
Event|Event|SIMPLE_SEGMENT|8001,8009|false|false|false|||vomiting
Finding|Sign or Symptom|SIMPLE_SEGMENT|8001,8009|false|false|false|C0042963|Vomiting|vomiting
Finding|Intellectual Product|SIMPLE_SEGMENT|8014,8018|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Event|Event|SIMPLE_SEGMENT|8022,8028|false|false|false|||intake
Finding|Functional Concept|SIMPLE_SEGMENT|8022,8028|false|true|false|C1512806|Intake|intake
Procedure|Health Care Activity|SIMPLE_SEGMENT|8022,8028|false|true|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|intake
Finding|Finding|SIMPLE_SEGMENT|8029,8035|false|true|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|8029,8035|false|true|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8045,8053|false|true|false|C1293134|Enlargement procedure|enlarged
Finding|Finding|SIMPLE_SEGMENT|8045,8059|false|true|false|C0019209|Hepatomegaly|enlarged liver
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8054,8059|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8054,8059|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8054,8059|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|SIMPLE_SEGMENT|8054,8059|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8054,8059|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|SIMPLE_SEGMENT|8054,8059|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|SIMPLE_SEGMENT|8054,8059|false|false|false|||liver
Finding|Finding|SIMPLE_SEGMENT|8054,8059|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|SIMPLE_SEGMENT|8054,8059|false|false|false|C0872387|Procedures on liver|liver
Event|Event|SIMPLE_SEGMENT|8066,8075|false|false|false|||continues
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8084,8089|false|false|false|C0021853|Intestines|bowel
Finding|Organism Function|SIMPLE_SEGMENT|8084,8099|false|false|false|C0011135|Defecation|bowel movements
Event|Event|SIMPLE_SEGMENT|8090,8099|false|false|false|||movements
Finding|Organism Function|SIMPLE_SEGMENT|8090,8099|false|false|false|C0026649|Movement|movements
Finding|Finding|SIMPLE_SEGMENT|8104,8108|false|false|false|C2828386|Pass (indicator)|pass
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8109,8112|false|false|false|C0017110;C1550641;C1704673|Gas - SpecimenType;Gas Dosage Form;Gases|gas
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|8109,8112|false|false|false|C0017110;C1550641;C1704673|Gas - SpecimenType;Gas Dosage Form;Gases|gas
Drug|Substance|SIMPLE_SEGMENT|8109,8112|false|false|false|C0017110;C1550641;C1704673|Gas - SpecimenType;Gas Dosage Form;Gases|gas
Event|Event|SIMPLE_SEGMENT|8109,8112|false|false|false|||gas
Finding|Gene or Genome|SIMPLE_SEGMENT|8109,8112|false|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|gas
Finding|Intellectual Product|SIMPLE_SEGMENT|8109,8112|false|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|gas
Finding|Molecular Function|SIMPLE_SEGMENT|8109,8112|false|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|gas
Finding|Sign or Symptom|SIMPLE_SEGMENT|8109,8112|false|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|gas
Finding|Body Substance|SIMPLE_SEGMENT|8114,8121|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|8114,8121|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|8114,8121|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8132,8139|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8132,8139|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8132,8139|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Event|Event|SIMPLE_SEGMENT|8132,8139|false|false|false|||albumin
Finding|Gene or Genome|SIMPLE_SEGMENT|8132,8139|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|albumin
Finding|Physiologic Function|SIMPLE_SEGMENT|8132,8139|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|albumin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8132,8139|false|false|false|C0201838|Albumin measurement|albumin
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|8148,8155|false|false|false|C0497010|Toxic effect of ketones|ketones
Drug|Organic Chemical|SIMPLE_SEGMENT|8148,8155|false|false|false|C0022634|Ketones|ketones
Event|Event|SIMPLE_SEGMENT|8148,8155|false|false|false|||ketones
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8148,8155|false|false|false|C0202110;C0555179|Ketone bodies measurement, quantitative;Urine ketone test|ketones
Event|Event|SIMPLE_SEGMENT|8163,8168|false|false|false|||urine
Finding|Body Substance|SIMPLE_SEGMENT|8163,8168|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|SIMPLE_SEGMENT|8163,8168|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|SIMPLE_SEGMENT|8163,8168|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8170,8176|false|false|false|C0944911||weight
Event|Event|SIMPLE_SEGMENT|8170,8176|false|false|false|||weight
Finding|Finding|SIMPLE_SEGMENT|8170,8176|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|8170,8176|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|8170,8176|false|false|false|C1305866|Weighing patient|weight
Finding|Finding|SIMPLE_SEGMENT|8170,8181|false|false|false|C1262477;C3540682|Losing Weight (question);Weight Loss|weight loss
Finding|Intellectual Product|SIMPLE_SEGMENT|8170,8181|false|false|false|C1262477;C3540682|Losing Weight (question);Weight Loss|weight loss
Event|Event|SIMPLE_SEGMENT|8177,8181|false|false|false|||loss
Finding|Finding|SIMPLE_SEGMENT|8177,8181|false|false|false|C5890125|Loss (adaptation)|loss
Finding|Finding|SIMPLE_SEGMENT|8186,8189|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|8186,8189|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Pathologic Function|SIMPLE_SEGMENT|8191,8207|false|false|false|C0085649|Peripheral edema|peripheral edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8202,8207|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|8202,8207|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|8202,8207|false|false|false|C0013604|Edema|edema
Finding|Intellectual Product|SIMPLE_SEGMENT|8224,8228|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8224,8238|false|false|false|C0162429|Malnutrition|poor nutrition
Event|Event|SIMPLE_SEGMENT|8229,8238|false|false|false|||nutrition
Finding|Finding|SIMPLE_SEGMENT|8229,8238|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|nutrition
Finding|Intellectual Product|SIMPLE_SEGMENT|8229,8238|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|nutrition
Finding|Organism Function|SIMPLE_SEGMENT|8229,8238|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|nutrition
Procedure|Research Activity|SIMPLE_SEGMENT|8229,8238|false|false|false|C0600072;C1521729|Feeding and dietary regimes;Nutritional Study|nutrition
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8229,8238|false|false|false|C0600072;C1521729|Feeding and dietary regimes;Nutritional Study|nutrition
Event|Event|SIMPLE_SEGMENT|8239,8249|false|false|false|||starvation
Finding|Finding|SIMPLE_SEGMENT|8239,8249|false|false|false|C0038187|Starvation|starvation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8251,8258|false|false|false|C0022638;C0220982|Ketoacidosis;Ketosis|ketosis
Event|Event|SIMPLE_SEGMENT|8251,8258|false|false|false|||ketosis
Event|Event|SIMPLE_SEGMENT|8260,8269|false|false|false|||Nutrition
Finding|Finding|SIMPLE_SEGMENT|8260,8269|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|Nutrition
Finding|Intellectual Product|SIMPLE_SEGMENT|8260,8269|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|Nutrition
Finding|Organism Function|SIMPLE_SEGMENT|8260,8269|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|Nutrition
Procedure|Research Activity|SIMPLE_SEGMENT|8260,8269|false|false|false|C0600072;C1521729|Feeding and dietary regimes;Nutritional Study|Nutrition
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8260,8269|false|false|false|C0600072;C1521729|Feeding and dietary regimes;Nutritional Study|Nutrition
Event|Event|SIMPLE_SEGMENT|8270,8277|false|false|false|||consult
Procedure|Health Care Activity|SIMPLE_SEGMENT|8270,8277|false|false|false|C0009818|Consultation|consult
Finding|Body Substance|SIMPLE_SEGMENT|8291,8298|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|8291,8298|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|8291,8298|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|8315,8323|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|SIMPLE_SEGMENT|8324,8328|false|false|false|||stay
Event|Event|SIMPLE_SEGMENT|8333,8344|false|false|false|||recommended
Anatomy|Tissue|SIMPLE_SEGMENT|8349,8352|false|false|false|C0001527|Adipose tissue|fat
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8349,8352|false|false|false|C0015677;C1435181;C3887682|FAT1 protein, human;Fatty acid glycerol esters;Platelet Glycoprotein 4, human|fat
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8349,8352|false|false|false|C0015677;C1435181;C3887682|FAT1 protein, human;Fatty acid glycerol esters;Platelet Glycoprotein 4, human|fat
Drug|Organic Chemical|SIMPLE_SEGMENT|8349,8352|false|false|false|C0015677;C1435181;C3887682|FAT1 protein, human;Fatty acid glycerol esters;Platelet Glycoprotein 4, human|fat
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8349,8352|false|false|false|C0015677;C1435181;C3887682|FAT1 protein, human;Fatty acid glycerol esters;Platelet Glycoprotein 4, human|fat
Finding|Gene or Genome|SIMPLE_SEGMENT|8349,8352|false|false|false|C0812278;C1366645;C1705088;C1708004;C3887682|CD36 gene;CD36 wt Allele;FAT1 gene;FAT1 wt Allele;Platelet Glycoprotein 4, human|fat
Finding|Receptor|SIMPLE_SEGMENT|8349,8352|false|false|false|C0812278;C1366645;C1705088;C1708004;C3887682|CD36 gene;CD36 wt Allele;FAT1 gene;FAT1 wt Allele;Platelet Glycoprotein 4, human|fat
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8349,8352|false|false|false|C0279453|doxorubicin/fluorouracil/triazinate protocol|fat
Drug|Food|SIMPLE_SEGMENT|8353,8370|false|false|false|C1874731|CARNATION INSTANT|Carnation Instant
Event|Event|SIMPLE_SEGMENT|8372,8381|false|false|false|||Breakfast
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|8372,8381|false|false|false|C2698559|Breakfast|Breakfast
Finding|Intellectual Product|SIMPLE_SEGMENT|8404,8411|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|8404,8411|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Finding|Sign or Symptom|SIMPLE_SEGMENT|8404,8421|false|false|false|C0740418|Chronic back pain|Chronic back pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|8412,8421|false|false|false|C0004604|Back Pain|back pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8417,8421|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|8417,8421|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|8417,8421|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|8417,8421|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Body Substance|SIMPLE_SEGMENT|8424,8431|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|8424,8431|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|8424,8431|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|8436,8445|false|false|false|||continued
Event|Event|SIMPLE_SEGMENT|8453,8457|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|8453,8457|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|8453,8457|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|8453,8457|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|8459,8469|false|false|false|C0060926|gabapentin|gabapentin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8459,8469|false|false|false|C0060926|gabapentin|gabapentin
Event|Event|SIMPLE_SEGMENT|8459,8469|false|false|false|||gabapentin
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8476,8486|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|Depression
Event|Event|SIMPLE_SEGMENT|8476,8486|false|false|false|||Depression
Finding|Functional Concept|SIMPLE_SEGMENT|8476,8486|false|false|false|C0460137;C1579931|Depression - motion|Depression
Finding|Sign or Symptom|SIMPLE_SEGMENT|8476,8486|false|false|false|C0460137;C1579931|Depression - motion|Depression
Finding|Body Substance|SIMPLE_SEGMENT|8489,8496|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|8489,8496|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|8489,8496|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|8501,8510|false|false|false|||continued
Finding|Idea or Concept|SIMPLE_SEGMENT|8514,8518|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|8514,8518|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|8514,8518|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|8519,8528|false|false|false|C0085208|bupropion|bupropion
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8519,8528|false|false|false|C0085208|bupropion|bupropion
Event|Event|SIMPLE_SEGMENT|8519,8528|false|false|false|||bupropion
Drug|Organic Chemical|SIMPLE_SEGMENT|8531,8541|false|false|false|C0074393|sertraline|sertraline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8531,8541|false|false|false|C0074393|sertraline|sertraline
Event|Event|SIMPLE_SEGMENT|8531,8541|false|false|false|||sertraline
Drug|Organic Chemical|SIMPLE_SEGMENT|8548,8552|false|false|false|C0020261|hydrochlorothiazide|HCTZ
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8548,8552|false|false|false|C0020261|hydrochlorothiazide|HCTZ
Event|Event|SIMPLE_SEGMENT|8548,8552|false|false|false|||HCTZ
Finding|Body Substance|SIMPLE_SEGMENT|8554,8561|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|8554,8561|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|8554,8561|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Organic Chemical|SIMPLE_SEGMENT|8564,8568|false|false|false|C0020261|hydrochlorothiazide|hctz
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8564,8568|false|false|false|C0020261|hydrochlorothiazide|hctz
Event|Event|SIMPLE_SEGMENT|8564,8568|false|false|false|||hctz
Event|Event|SIMPLE_SEGMENT|8573,8585|false|false|false|||discontinued
Event|Event|SIMPLE_SEGMENT|8598,8613|false|false|false|||hospitalization
Procedure|Health Care Activity|SIMPLE_SEGMENT|8598,8613|false|false|false|C0019993|Hospitalization|hospitalization
Finding|Intellectual Product|SIMPLE_SEGMENT|8621,8625|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Event|Event|SIMPLE_SEGMENT|8629,8635|false|false|false|||intake
Finding|Functional Concept|SIMPLE_SEGMENT|8629,8635|false|false|false|C1512806|Intake|intake
Procedure|Health Care Activity|SIMPLE_SEGMENT|8629,8635|false|false|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|intake
Event|Event|SIMPLE_SEGMENT|8640,8647|false|false|false|||concern
Finding|Idea or Concept|SIMPLE_SEGMENT|8640,8647|false|false|false|C2699424|Concern|concern
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8653,8664|false|false|false|C0011175;C2062903|Dehydration;dehydration (Na, H2O)|dehydration
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|8653,8664|false|false|false|C0011175;C2062903|Dehydration;dehydration (Na, H2O)|dehydration
Event|Event|SIMPLE_SEGMENT|8653,8664|false|false|false|||dehydration
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8653,8664|false|false|false|C4284399|Dehydration procedure|dehydration
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8666,8671|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Finding|Body Substance|SIMPLE_SEGMENT|8666,8671|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Finding|Finding|SIMPLE_SEGMENT|8666,8681|false|false|false|C1272641|Systemic arterial pressure|Blood pressures
Event|Event|SIMPLE_SEGMENT|8672,8681|false|false|false|||pressures
Finding|Finding|SIMPLE_SEGMENT|8672,8681|false|false|false|C0460139|Pressure (finding)|pressures
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|8672,8681|false|false|false|C0033095||pressures
Finding|Finding|SIMPLE_SEGMENT|8687,8691|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|8692,8702|false|false|false|||controlled
Drug|Organic Chemical|SIMPLE_SEGMENT|8713,8717|false|false|false|C0020261|hydrochlorothiazide|HCTZ
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8713,8717|false|false|false|C0020261|hydrochlorothiazide|HCTZ
Event|Event|SIMPLE_SEGMENT|8713,8717|false|false|false|||HCTZ
Event|Event|SIMPLE_SEGMENT|8727,8733|false|false|false|||deemed
Event|Event|SIMPLE_SEGMENT|8734,8743|false|false|false|||necessary
Event|Activity|SIMPLE_SEGMENT|8750,8755|false|false|false|C5966184|Issue (action)|issue
Event|Event|SIMPLE_SEGMENT|8750,8755|false|false|false|||issue
Finding|Finding|SIMPLE_SEGMENT|8750,8755|false|false|false|C0033213;C1706387|Issue (document);Problem|issue
Finding|Intellectual Product|SIMPLE_SEGMENT|8750,8755|false|false|false|C0033213;C1706387|Issue (document);Problem|issue
Event|Event|SIMPLE_SEGMENT|8766,8777|false|false|false|||readdressed
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8782,8785|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8782,8785|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8782,8785|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8782,8785|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|8782,8785|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|8782,8785|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|8782,8785|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8782,8785|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|8782,8785|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|8782,8785|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|8782,8785|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8791,8805|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|Hyperlipidemia
Event|Event|SIMPLE_SEGMENT|8791,8805|false|false|false|||Hyperlipidemia
Finding|Finding|SIMPLE_SEGMENT|8791,8805|false|false|false|C0428465|Serum lipids high (finding)|Hyperlipidemia
Finding|Body Substance|SIMPLE_SEGMENT|8813,8820|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|8813,8820|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|8813,8820|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|SIMPLE_SEGMENT|8823,8833|false|false|false|C0036525;C1522484|Metastatic to;metastatic qualifier|metastatic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8834,8841|false|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8834,8841|false|false|false|C1951340|Process Pharmacologic Substance|process
Event|Event|SIMPLE_SEGMENT|8834,8841|false|false|false|||process
Finding|Functional Concept|SIMPLE_SEGMENT|8834,8841|false|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|8834,8841|false|false|false|C1522240|Process|process
Drug|Organic Chemical|SIMPLE_SEGMENT|8843,8849|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|statin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8843,8849|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|statin
Event|Event|SIMPLE_SEGMENT|8843,8849|false|false|false|||statin
Finding|Gene or Genome|SIMPLE_SEGMENT|8843,8849|false|false|false|C1414273|EEF1A2 gene|statin
Event|Event|SIMPLE_SEGMENT|8855,8867|false|false|false|||discontinued
Event|Event|SIMPLE_SEGMENT|8875,8890|false|false|false|||hospitalization
Procedure|Health Care Activity|SIMPLE_SEGMENT|8875,8890|false|false|false|C0019993|Hospitalization|hospitalization
Event|Event|SIMPLE_SEGMENT|8894,8902|false|false|false|||simplify
Event|Event|SIMPLE_SEGMENT|8907,8914|false|false|false|||medical
Finding|Functional Concept|SIMPLE_SEGMENT|8907,8914|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|SIMPLE_SEGMENT|8907,8914|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|SIMPLE_SEGMENT|8907,8914|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|8907,8914|false|false|false|C0199168|Medical service|medical
Event|Event|SIMPLE_SEGMENT|8916,8923|false|false|false|||regimen
Finding|Intellectual Product|SIMPLE_SEGMENT|8916,8923|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8916,8923|false|false|false|C0040808|Treatment Protocols|regimen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8931,8939|false|false|false|C1950154|Insomnia homeopathic medication|Insomnia
Event|Event|SIMPLE_SEGMENT|8931,8939|false|false|false|||Insomnia
Finding|Sign or Symptom|SIMPLE_SEGMENT|8931,8939|false|false|false|C0917801|Sleeplessness|Insomnia
Event|Event|SIMPLE_SEGMENT|8941,8950|false|false|false|||Continued
Finding|Idea or Concept|SIMPLE_SEGMENT|8951,8955|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|8951,8955|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|8951,8955|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|8956,8965|false|false|false|C0040805|trazodone|trazodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8956,8965|false|false|false|C0040805|trazodone|trazodone
Event|Event|SIMPLE_SEGMENT|8956,8965|false|false|false|||trazodone
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|8970,8980|false|false|false|C0599156|Transition Mutation|TRANSITION
Event|Activity|SIMPLE_SEGMENT|8970,8980|false|false|false|C2700061|Transition (action)|TRANSITION
Event|Event|SIMPLE_SEGMENT|8981,8987|false|false|false|||ISSUES
Event|Event|SIMPLE_SEGMENT|8990,8994|false|false|false|||CODE
Event|Occupational Activity|SIMPLE_SEGMENT|8990,8994|false|false|false|C0009219|Coding|CODE
Finding|Intellectual Product|SIMPLE_SEGMENT|8990,8994|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|CODE
Finding|Finding|SIMPLE_SEGMENT|9002,9011|false|false|false|C0750484|Confirmation|Confirmed
Event|Activity|SIMPLE_SEGMENT|9017,9024|false|false|false|C3812666|Personal Contact|CONTACT
Event|Event|SIMPLE_SEGMENT|9017,9024|false|false|false|||CONTACT
Finding|Functional Concept|SIMPLE_SEGMENT|9017,9024|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Idea or Concept|SIMPLE_SEGMENT|9017,9024|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Intellectual Product|SIMPLE_SEGMENT|9017,9024|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|9017,9024|false|false|false|C0392367|Physical contact|CONTACT
Finding|Idea or Concept|SIMPLE_SEGMENT|9031,9037|false|false|false|C1546502|Relationship - Friend|friend
Drug|Organic Chemical|SIMPLE_SEGMENT|9047,9051|false|false|false|C0020261|hydrochlorothiazide|HCTZ
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9047,9051|false|false|false|C0020261|hydrochlorothiazide|HCTZ
Event|Event|SIMPLE_SEGMENT|9047,9051|false|false|false|||HCTZ
Event|Event|SIMPLE_SEGMENT|9052,9064|false|false|false|||discontinued
Event|Event|SIMPLE_SEGMENT|9068,9077|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|9068,9077|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|9079,9087|false|false|false|||consider
Finding|Idea or Concept|SIMPLE_SEGMENT|9079,9087|false|false|false|C0750591|consider|consider
Event|Event|SIMPLE_SEGMENT|9103,9113|false|false|false|||considered
Event|Event|SIMPLE_SEGMENT|9124,9133|false|false|false|||necessary
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9137,9140|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9137,9140|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|9137,9140|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9137,9140|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|9137,9140|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|9137,9140|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|9137,9140|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9137,9140|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|9137,9140|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|9137,9140|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|9137,9140|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Anatomy|Tissue|SIMPLE_SEGMENT|9148,9151|false|false|false|C0001527|Adipose tissue|fat
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9148,9151|false|false|false|C0015677;C1435181;C3887682|FAT1 protein, human;Fatty acid glycerol esters;Platelet Glycoprotein 4, human|fat
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9148,9151|false|false|false|C0015677;C1435181;C3887682|FAT1 protein, human;Fatty acid glycerol esters;Platelet Glycoprotein 4, human|fat
Drug|Organic Chemical|SIMPLE_SEGMENT|9148,9151|false|false|false|C0015677;C1435181;C3887682|FAT1 protein, human;Fatty acid glycerol esters;Platelet Glycoprotein 4, human|fat
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9148,9151|false|false|false|C0015677;C1435181;C3887682|FAT1 protein, human;Fatty acid glycerol esters;Platelet Glycoprotein 4, human|fat
Finding|Gene or Genome|SIMPLE_SEGMENT|9148,9151|false|false|false|C0812278;C1366645;C1705088;C1708004;C3887682|CD36 gene;CD36 wt Allele;FAT1 gene;FAT1 wt Allele;Platelet Glycoprotein 4, human|fat
Finding|Receptor|SIMPLE_SEGMENT|9148,9151|false|false|false|C0812278;C1366645;C1705088;C1708004;C3887682|CD36 gene;CD36 wt Allele;FAT1 gene;FAT1 wt Allele;Platelet Glycoprotein 4, human|fat
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9148,9151|false|false|false|C0279453|doxorubicin/fluorouracil/triazinate protocol|fat
Drug|Food|SIMPLE_SEGMENT|9152,9169|false|false|false|C1874731|CARNATION INSTANT|Carnation Instant
Event|Event|SIMPLE_SEGMENT|9170,9179|false|false|false|||Breakfast
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|9170,9179|false|false|false|C2698559|Breakfast|Breakfast
Event|Event|SIMPLE_SEGMENT|9203,9208|false|false|false|||meals
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|9203,9208|false|false|false|C1998602|Meal (occasion for eating)|meals
Event|Event|SIMPLE_SEGMENT|9211,9217|false|false|false|||Follow
Disorder|Neoplastic Process|SIMPLE_SEGMENT|9226,9234|false|false|false|C0027651|Neoplasms|oncology
Event|Event|SIMPLE_SEGMENT|9226,9234|false|false|false|||oncology
Procedure|Health Care Activity|SIMPLE_SEGMENT|9226,9234|false|false|false|C1555459|oncology services|oncology
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9247,9256|false|false|false|C0945731||diagnosis
Event|Event|SIMPLE_SEGMENT|9247,9256|false|false|false|||diagnosis
Finding|Classification|SIMPLE_SEGMENT|9247,9256|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|9247,9256|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9247,9256|false|false|false|C0011900|Diagnosis|diagnosis
Event|Event|SIMPLE_SEGMENT|9261,9271|false|false|false|||management
Event|Occupational Activity|SIMPLE_SEGMENT|9261,9271|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|SIMPLE_SEGMENT|9261,9271|false|false|false|C0376636|Disease Management|management
Disorder|Neoplastic Process|SIMPLE_SEGMENT|9276,9286|false|false|false|C0006826;C1306459|Malignant Neoplasms;Primary malignant neoplasm|malignancy
Event|Event|SIMPLE_SEGMENT|9276,9286|false|false|false|||malignancy
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9289,9300|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9289,9300|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|9289,9300|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|9289,9300|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|9289,9313|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|SIMPLE_SEGMENT|9304,9313|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|9304,9313|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9332,9342|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|9332,9342|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|9332,9347|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|SIMPLE_SEGMENT|9343,9347|false|false|false|||list
Finding|Intellectual Product|SIMPLE_SEGMENT|9343,9347|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|SIMPLE_SEGMENT|9351,9359|false|false|false|||accurate
Drug|Organic Chemical|SIMPLE_SEGMENT|9364,9372|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9364,9372|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|9364,9372|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|SIMPLE_SEGMENT|9364,9372|false|false|false|||complete
Finding|Functional Concept|SIMPLE_SEGMENT|9364,9372|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|9364,9372|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|SIMPLE_SEGMENT|9377,9386|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9377,9386|false|false|false|C0001927|albuterol|Albuterol
Finding|Functional Concept|SIMPLE_SEGMENT|9387,9394|false|false|false|C4319647|Inhaler (unit of presentation)|Inhaler
Finding|Gene or Genome|SIMPLE_SEGMENT|9411,9414|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|9415,9418|false|false|false|||SOB
Finding|Sign or Symptom|SIMPLE_SEGMENT|9415,9418|false|false|false|C0013404|Dyspnea|SOB
Drug|Organic Chemical|SIMPLE_SEGMENT|9423,9432|false|false|false|C0085208|bupropion|BuPROPion
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9423,9432|false|false|false|C0085208|bupropion|BuPROPion
Drug|Organic Chemical|SIMPLE_SEGMENT|9453,9463|false|false|false|C0060926|gabapentin|Gabapentin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9453,9463|false|false|false|C0060926|gabapentin|Gabapentin
Drug|Organic Chemical|SIMPLE_SEGMENT|9481,9491|false|false|false|C0074393|sertraline|Sertraline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9481,9491|false|false|false|C0074393|sertraline|Sertraline
Drug|Organic Chemical|SIMPLE_SEGMENT|9512,9523|false|false|false|C0074554|simvastatin|Simvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9512,9523|false|false|false|C0074554|simvastatin|Simvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|9543,9552|false|false|false|C0040805|trazodone|traZODONE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9543,9552|false|false|false|C0040805|trazodone|traZODONE
Event|Event|SIMPLE_SEGMENT|9543,9552|false|false|false|||traZODONE
Finding|Gene or Genome|SIMPLE_SEGMENT|9566,9569|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|SIMPLE_SEGMENT|9570,9575|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9570,9575|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Event|Event|SIMPLE_SEGMENT|9570,9575|false|false|false|||sleep
Finding|Organism Function|SIMPLE_SEGMENT|9570,9575|false|false|false|C0037313|Sleep|sleep
Drug|Organic Chemical|SIMPLE_SEGMENT|9580,9589|false|false|false|C0020740|ibuprofen|Ibuprofen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9580,9589|false|false|false|C0020740|ibuprofen|Ibuprofen
Finding|Gene or Genome|SIMPLE_SEGMENT|9605,9608|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9609,9613|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|9609,9613|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9609,9613|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9609,9613|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|9618,9637|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9618,9637|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Organic Chemical|SIMPLE_SEGMENT|9659,9670|false|false|false|C0061851|ondansetron|Ondansetron
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9659,9670|false|false|false|C0061851|ondansetron|Ondansetron
Finding|Gene or Genome|SIMPLE_SEGMENT|9683,9686|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9687,9693|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|9687,9693|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|9687,9693|false|false|false|C0027497|Nausea|nausea
Event|Event|SIMPLE_SEGMENT|9698,9707|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|9698,9707|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|9698,9707|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|9698,9707|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|9698,9707|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|9698,9719|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9708,9719|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9708,9719|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|9708,9719|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|9708,9719|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|9724,9733|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9724,9733|false|false|false|C0001927|albuterol|Albuterol
Finding|Functional Concept|SIMPLE_SEGMENT|9734,9741|false|false|false|C4319647|Inhaler (unit of presentation)|Inhaler
Finding|Gene or Genome|SIMPLE_SEGMENT|9758,9761|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|9762,9765|false|false|false|||SOB
Finding|Sign or Symptom|SIMPLE_SEGMENT|9762,9765|false|false|false|C0013404|Dyspnea|SOB
Drug|Organic Chemical|SIMPLE_SEGMENT|9770,9779|false|false|false|C0085208|bupropion|BuPROPion
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9770,9779|false|false|false|C0085208|bupropion|BuPROPion
Drug|Organic Chemical|SIMPLE_SEGMENT|9800,9810|false|false|false|C0060926|gabapentin|Gabapentin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9800,9810|false|false|false|C0060926|gabapentin|Gabapentin
Drug|Organic Chemical|SIMPLE_SEGMENT|9828,9838|false|false|false|C0074393|sertraline|Sertraline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9828,9838|false|false|false|C0074393|sertraline|Sertraline
Drug|Organic Chemical|SIMPLE_SEGMENT|9859,9868|false|false|false|C0040805|trazodone|traZODONE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9859,9868|false|false|false|C0040805|trazodone|traZODONE
Finding|Gene or Genome|SIMPLE_SEGMENT|9882,9885|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|SIMPLE_SEGMENT|9886,9891|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9886,9891|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Event|Event|SIMPLE_SEGMENT|9886,9891|false|false|false|||sleep
Finding|Organism Function|SIMPLE_SEGMENT|9886,9891|false|false|false|C0037313|Sleep|sleep
Drug|Organic Chemical|SIMPLE_SEGMENT|9896,9907|false|false|false|C0061851|ondansetron|Ondansetron
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9896,9907|false|false|false|C0061851|ondansetron|Ondansetron
Finding|Gene or Genome|SIMPLE_SEGMENT|9920,9923|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9924,9930|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|9924,9930|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|9924,9930|false|false|false|C0027497|Nausea|nausea
Drug|Organic Chemical|SIMPLE_SEGMENT|9935,9944|false|false|false|C0005632|bisacodyl|Bisacodyl
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9935,9944|false|false|false|C0005632|bisacodyl|Bisacodyl
Finding|Gene or Genome|SIMPLE_SEGMENT|9963,9966|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|9967,9979|false|false|false|||constipation
Finding|Sign or Symptom|SIMPLE_SEGMENT|9967,9979|false|false|false|C0009806|Constipation|constipation
Drug|Organic Chemical|SIMPLE_SEGMENT|9984,9993|false|false|false|C0030049|oxycodone|OxycoDONE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9984,9993|false|false|false|C0030049|oxycodone|OxycoDONE
Event|Event|SIMPLE_SEGMENT|9984,9993|false|false|false|||OxycoDONE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9984,9993|false|false|false|C0524222|Oxycodone measurement|OxycoDONE
Finding|Idea or Concept|SIMPLE_SEGMENT|9995,10004|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Finding|Intellectual Product|SIMPLE_SEGMENT|9995,10004|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9995,10012|false|false|false|C1708470|Immediate Release Dosage Form|Immediate Release
Event|Event|SIMPLE_SEGMENT|10005,10012|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|10005,10012|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|10005,10012|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10005,10012|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Finding|Gene or Genome|SIMPLE_SEGMENT|10027,10030|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10031,10035|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|10031,10035|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|10031,10035|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|10031,10035|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|10044,10048|false|false|false|||hold
Event|Event|SIMPLE_SEGMENT|10053,10061|false|false|false|||sedation
Finding|Finding|SIMPLE_SEGMENT|10053,10061|false|false|false|C0235195;C5400562|Sedated state;Sedation|sedation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10053,10061|false|false|false|C0344106|Sedation procedure|sedation
Event|Event|SIMPLE_SEGMENT|10070,10072|false|false|false|||RX
Drug|Organic Chemical|SIMPLE_SEGMENT|10074,10083|false|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10074,10083|false|false|false|C0030049|oxycodone|oxycodone
Event|Event|SIMPLE_SEGMENT|10074,10083|false|false|false|||oxycodone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10074,10083|false|false|false|C0524222|Oxycodone measurement|oxycodone
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10091,10097|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|SIMPLE_SEGMENT|10101,10109|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10104,10109|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|10104,10109|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|10135,10141|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|10142,10149|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|10142,10149|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|10156,10166|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10156,10166|false|false|false|C0206460|enoxaparin|Enoxaparin
Event|Event|SIMPLE_SEGMENT|10156,10166|false|false|false|||Enoxaparin
Drug|Organic Chemical|SIMPLE_SEGMENT|10156,10173|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10156,10173|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10167,10173|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|10167,10173|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10167,10173|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|10167,10173|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|10167,10173|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10167,10173|false|false|false|C0337443|Sodium measurement|Sodium
Event|Event|SIMPLE_SEGMENT|10193,10202|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|10193,10202|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10193,10202|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|10193,10202|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|10193,10202|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10193,10214|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|10193,10214|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10203,10214|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|10203,10214|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|10203,10214|false|false|false|C0184758|Patient disposition|Disposition
Finding|Finding|SIMPLE_SEGMENT|10216,10224|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|10216,10224|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Procedure|Health Care Activity|SIMPLE_SEGMENT|10216,10229|false|false|false|C0023977|long-term care|Extended Care
Event|Activity|SIMPLE_SEGMENT|10225,10229|false|false|false|C1947933|care activity|Care
Event|Event|SIMPLE_SEGMENT|10225,10229|false|false|false|||Care
Finding|Finding|SIMPLE_SEGMENT|10225,10229|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|SIMPLE_SEGMENT|10225,10229|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Event|Event|SIMPLE_SEGMENT|10232,10240|false|false|false|||Facility
Finding|Intellectual Product|SIMPLE_SEGMENT|10232,10240|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|SIMPLE_SEGMENT|10248,10257|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|10248,10257|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10248,10257|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|10248,10257|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|10248,10257|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|10248,10267|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10258,10267|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|10258,10267|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|10258,10267|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|10258,10267|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10258,10267|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|10269,10279|false|false|false|C0036525;C1522484|Metastatic to;metastatic qualifier|Metastatic
Disorder|Neoplastic Process|SIMPLE_SEGMENT|10269,10287|false|false|false|C0027627;C2939419;C2939420|Metastatic Neoplasm;Metastatic malignant neoplasm;Neoplasm Metastasis|Metastatic disease
Finding|Finding|SIMPLE_SEGMENT|10269,10287|false|false|false|C1513183|Metastatic Lesion|Metastatic disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10280,10287|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|10280,10287|false|false|false|||disease
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10291,10298|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Immunologic Factor|SIMPLE_SEGMENT|10291,10298|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10291,10298|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Event|Event|SIMPLE_SEGMENT|10291,10298|false|false|false|||unknown
Finding|Finding|SIMPLE_SEGMENT|10291,10298|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Functional Concept|SIMPLE_SEGMENT|10291,10298|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Idea or Concept|SIMPLE_SEGMENT|10291,10298|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Intellectual Product|SIMPLE_SEGMENT|10291,10298|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Event|Event|SIMPLE_SEGMENT|10308,10316|false|false|false|||Weakness
Finding|Sign or Symptom|SIMPLE_SEGMENT|10308,10316|false|false|false|C0004093;C3714552|Asthenia;Weakness|Weakness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10321,10327|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|10321,10327|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|10321,10327|false|false|false|C0027497|Nausea|nausea
Finding|Finding|SIMPLE_SEGMENT|10329,10335|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|10329,10335|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Disorder|Neoplastic Process|SIMPLE_SEGMENT|10341,10346|false|true|false|C0027651|Neoplasms|tumor
Finding|Finding|SIMPLE_SEGMENT|10341,10346|false|true|false|C1578706;C3273930|Tumor Mass|tumor
Finding|Intellectual Product|SIMPLE_SEGMENT|10341,10346|false|true|false|C1578706;C3273930|Tumor Mass|tumor
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10341,10353|false|true|false|C1449699|Tumor Burden|tumor burden
Event|Event|SIMPLE_SEGMENT|10347,10353|false|false|false|||burden
Finding|Idea or Concept|SIMPLE_SEGMENT|10347,10353|false|true|false|C2828008|Burden|burden
Event|Event|SIMPLE_SEGMENT|10357,10366|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|10357,10366|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10357,10366|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|10357,10366|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|10357,10366|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10367,10376|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10367,10376|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|10367,10376|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|10367,10376|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|10378,10384|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10378,10391|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|10378,10391|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10385,10391|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|10385,10391|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|10393,10398|false|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|10393,10398|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|10403,10411|false|false|false|||coherent
Finding|Finding|SIMPLE_SEGMENT|10403,10411|false|false|false|C4068804|Coherent|coherent
Event|Event|SIMPLE_SEGMENT|10413,10418|false|false|false|||Level
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10413,10435|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|10413,10435|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|SIMPLE_SEGMENT|10422,10435|false|false|false|||Consciousness
Finding|Finding|SIMPLE_SEGMENT|10422,10435|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|10422,10435|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10437,10442|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|10437,10442|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10437,10442|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|10437,10442|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|10437,10442|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|10437,10442|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|10437,10442|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|10447,10458|false|false|false|||interactive
Finding|Functional Concept|SIMPLE_SEGMENT|10447,10458|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|10460,10468|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|10460,10468|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|10460,10468|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10469,10475|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|10469,10475|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|10469,10475|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|10477,10487|false|false|false|||Ambulatory
Finding|Functional Concept|SIMPLE_SEGMENT|10477,10487|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|10477,10487|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|10477,10487|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|10477,10487|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|SIMPLE_SEGMENT|10490,10501|false|false|false|||Independent
Finding|Finding|SIMPLE_SEGMENT|10490,10501|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|SIMPLE_SEGMENT|10490,10501|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Event|Event|SIMPLE_SEGMENT|10506,10515|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|10506,10515|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|10506,10515|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|10506,10515|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|10506,10515|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10506,10528|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|10506,10528|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|10506,10528|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10516,10528|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|10516,10528|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|10516,10528|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Finding|Gene or Genome|SIMPLE_SEGMENT|10530,10534|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|SIMPLE_SEGMENT|10554,10562|false|false|false|||admitted
Event|Event|SIMPLE_SEGMENT|10574,10584|false|false|false|||evaluation
Finding|Idea or Concept|SIMPLE_SEGMENT|10574,10584|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|SIMPLE_SEGMENT|10574,10584|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Event|Event|SIMPLE_SEGMENT|10606,10614|false|false|false|||weakness
Finding|Sign or Symptom|SIMPLE_SEGMENT|10606,10614|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10619,10625|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|10619,10625|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|10619,10625|false|false|false|C0027497|Nausea|nausea
Event|Event|SIMPLE_SEGMENT|10640,10647|false|false|false|||markers
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10651,10660|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|10651,10660|false|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|10651,10660|false|false|false|C3714514|Infection|infection
Drug|Antibiotic|SIMPLE_SEGMENT|10691,10702|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|SIMPLE_SEGMENT|10691,10702|false|false|false|||antibiotics
Event|Event|SIMPLE_SEGMENT|10715,10719|false|false|false|||scan
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10715,10719|false|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10728,10733|false|false|false|C0460005|Trunk structure|torso
Event|Event|SIMPLE_SEGMENT|10735,10741|false|false|false|||showed
Finding|Functional Concept|SIMPLE_SEGMENT|10742,10752|false|false|false|C0036525;C1522484|Metastatic to;metastatic qualifier|metastatic
Disorder|Neoplastic Process|SIMPLE_SEGMENT|10742,10760|false|false|false|C0027627;C2939419;C2939420|Metastatic Neoplasm;Metastatic malignant neoplasm;Neoplasm Metastasis|metastatic disease
Finding|Finding|SIMPLE_SEGMENT|10742,10760|false|false|false|C1513183|Metastatic Lesion|metastatic disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10753,10760|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|10753,10760|false|false|false|||disease
Disorder|Neoplastic Process|SIMPLE_SEGMENT|10768,10774|false|true|false|C0006826|Malignant Neoplasms|cancer
Event|Event|SIMPLE_SEGMENT|10768,10774|false|false|false|||cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|10768,10792|false|false|false|C0220647|Carcinoma of unknown primary|cancer of unknown origin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10778,10785|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Immunologic Factor|SIMPLE_SEGMENT|10778,10785|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10778,10785|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Event|Event|SIMPLE_SEGMENT|10778,10785|false|false|false|||unknown
Finding|Finding|SIMPLE_SEGMENT|10778,10785|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Functional Concept|SIMPLE_SEGMENT|10778,10785|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Idea or Concept|SIMPLE_SEGMENT|10778,10785|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Intellectual Product|SIMPLE_SEGMENT|10778,10785|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Functional Concept|SIMPLE_SEGMENT|10778,10792|false|false|false|C0332240|Unknown (origin) (qualifier value)|unknown origin
Event|Event|SIMPLE_SEGMENT|10786,10792|false|false|false|||origin
Finding|Classification|SIMPLE_SEGMENT|10786,10792|false|false|false|C0079946;C1550512|National origin;Participation Type - origin|origin
Finding|Intellectual Product|SIMPLE_SEGMENT|10786,10792|false|false|false|C0079946;C1550512|National origin;Participation Type - origin|origin
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10802,10807|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10802,10807|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|SIMPLE_SEGMENT|10802,10807|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|SIMPLE_SEGMENT|10802,10807|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10802,10807|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|SIMPLE_SEGMENT|10802,10807|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|SIMPLE_SEGMENT|10802,10807|false|false|false|||liver
Finding|Finding|SIMPLE_SEGMENT|10802,10807|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|SIMPLE_SEGMENT|10802,10807|false|false|false|C0872387|Procedures on liver|liver
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10812,10817|false|false|false|C0024109|Lung|lungs
Event|Event|SIMPLE_SEGMENT|10824,10832|false|false|false|||weakness
Finding|Sign or Symptom|SIMPLE_SEGMENT|10824,10832|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10837,10843|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|10837,10843|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|10837,10843|false|false|false|C0027497|Nausea|nausea
Finding|Idea or Concept|SIMPLE_SEGMENT|10848,10859|false|false|false|C0750501|most likely|most likely
Event|Event|SIMPLE_SEGMENT|10853,10859|false|false|false|||likely
Finding|Finding|SIMPLE_SEGMENT|10853,10859|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|10853,10859|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10873,10881|false|false|false|C1293134|Enlargement procedure|enlarged
Finding|Finding|SIMPLE_SEGMENT|10873,10887|false|false|false|C0019209|Hepatomegaly|enlarged liver
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10882,10887|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10882,10887|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|SIMPLE_SEGMENT|10882,10887|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|SIMPLE_SEGMENT|10882,10887|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10882,10887|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|SIMPLE_SEGMENT|10882,10887|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|SIMPLE_SEGMENT|10882,10887|false|false|false|||liver
Finding|Finding|SIMPLE_SEGMENT|10882,10887|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|SIMPLE_SEGMENT|10882,10887|false|false|false|C0872387|Procedures on liver|liver
Event|Event|SIMPLE_SEGMENT|10899,10908|false|false|false|||scheduled
Event|Event|SIMPLE_SEGMENT|10912,10915|false|false|false|||see
Finding|Intellectual Product|SIMPLE_SEGMENT|10937,10941|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|SIMPLE_SEGMENT|10954,10960|false|false|false|||follow
Event|Event|SIMPLE_SEGMENT|10991,10998|false|false|false|||proceed
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11017,11026|false|false|false|C0945731||diagnosis
Event|Event|SIMPLE_SEGMENT|11017,11026|false|false|false|||diagnosis
Finding|Classification|SIMPLE_SEGMENT|11017,11026|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|11017,11026|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|11017,11026|false|false|false|C0011900|Diagnosis|diagnosis
Event|Event|SIMPLE_SEGMENT|11031,11040|false|false|false|||treatment
Finding|Conceptual Entity|SIMPLE_SEGMENT|11031,11040|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|SIMPLE_SEGMENT|11031,11040|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|SIMPLE_SEGMENT|11031,11040|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11031,11040|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Disorder|Neoplastic Process|SIMPLE_SEGMENT|11049,11059|false|false|false|C0006826;C1306459|Malignant Neoplasms;Primary malignant neoplasm|malignancy
Event|Event|SIMPLE_SEGMENT|11049,11059|false|false|false|||malignancy
Event|Event|SIMPLE_SEGMENT|11076,11086|false|false|false|||discharged
Event|Event|SIMPLE_SEGMENT|11092,11106|false|false|false|||rehabilitation
Finding|Finding|SIMPLE_SEGMENT|11092,11106|false|false|false|C0007237;C0034992|Encounter due to care involving use of rehabilitation procedures;Rehabilitation aspects|rehabilitation
Finding|Functional Concept|SIMPLE_SEGMENT|11092,11106|false|false|false|C0007237;C0034992|Encounter due to care involving use of rehabilitation procedures;Rehabilitation aspects|rehabilitation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11092,11106|false|false|false|C0034991|Rehabilitation therapy|rehabilitation
Event|Event|SIMPLE_SEGMENT|11107,11115|false|false|false|||facility
Finding|Intellectual Product|SIMPLE_SEGMENT|11107,11115|false|false|false|C4695111|ADMIN.FACILITY|facility
Event|Event|SIMPLE_SEGMENT|11119,11123|false|false|false|||help
Finding|Intellectual Product|SIMPLE_SEGMENT|11119,11123|false|false|false|C1552861|Help document|help
Drug|Food|SIMPLE_SEGMENT|11129,11135|false|false|false|C1875723|REGAIN|regain
Event|Event|SIMPLE_SEGMENT|11141,11149|false|false|false|||strength
Finding|Idea or Concept|SIMPLE_SEGMENT|11141,11149|false|false|false|C0808080|Strength (attribute)|strength
Event|Event|SIMPLE_SEGMENT|11163,11167|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|11163,11167|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|11163,11167|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|11163,11167|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|11174,11185|false|false|false|||anticipated
Finding|Finding|SIMPLE_SEGMENT|11174,11185|false|false|false|C3840775|Anticipated|anticipated
Event|Event|SIMPLE_SEGMENT|11205,11209|false|false|false|||LESS
Event|Event|SIMPLE_SEGMENT|11218,11222|false|false|false|||DAYS
Event|Event|SIMPLE_SEGMENT|11233,11236|false|false|false|||see
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|11241,11249|false|false|false|C3714578|Fix|attached
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11273,11283|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|11273,11283|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|11273,11283|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Finding|Intellectual Product|SIMPLE_SEGMENT|11273,11288|false|false|false|C0746470|MEDICATION LIST|medication list
Event|Event|SIMPLE_SEGMENT|11284,11288|false|false|false|||list
Finding|Intellectual Product|SIMPLE_SEGMENT|11284,11288|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|SIMPLE_SEGMENT|11301,11309|false|false|false|||pleasure
Finding|Intellectual Product|SIMPLE_SEGMENT|11301,11309|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|SIMPLE_SEGMENT|11301,11309|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|SIMPLE_SEGMENT|11317,11321|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|11317,11321|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|11317,11321|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|11317,11321|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|11317,11324|false|false|false|C1555558|care of - AddressPartType|care of
Finding|Idea or Concept|SIMPLE_SEGMENT|11336,11344|false|false|false|C1547192|Organization unit type - Hospital|hospital
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11349,11353|false|false|false|C3273412|NCK-Interacting Protein with SH3 Domain|wish
Event|Event|SIMPLE_SEGMENT|11349,11353|false|false|false|||wish
Finding|Gene or Genome|SIMPLE_SEGMENT|11349,11353|false|false|false|C1423524;C3273411|NCKIPSD gene;NCKIPSD wt Allele|wish
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11367,11371|false|false|false|C0339510|Vitelliform Macular Dystrophy|best
Event|Event|SIMPLE_SEGMENT|11367,11371|false|false|false|||best
Finding|Gene or Genome|SIMPLE_SEGMENT|11367,11371|false|false|false|C1826421;C5781213|BEST1 gene;BEST1 wt Allele|best
Procedure|Health Care Activity|SIMPLE_SEGMENT|11375,11383|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11384,11396|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|11384,11396|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|11384,11396|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

