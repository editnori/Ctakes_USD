 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|43,52|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|43,52|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|43,57|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|77,86|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|77,86|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|77,91|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|133,136|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|144,151|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|144,151|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|153,161|true|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|Allergies|185,194|true|false|false|C1717415||Allergies
Event|Event|Allergies|185,194|true|false|false|||Allergies
Finding|Pathologic Function|Allergies|185,194|true|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|Allergies|197,219|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|Allergies|205,209|true|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|Allergies|205,209|true|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|Allergies|205,219|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Event|Event|Allergies|210,219|true|false|false|||Reactions
Event|Event|Allergies|222,231|false|false|false|||Attending
Finding|Functional Concept|Allergies|222,231|false|false|false|C1999232|Attending (action)|Attending
Event|Event|Chief Complaint|257,264|false|false|false|||dyspnea
Finding|Finding|Chief Complaint|257,264|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|Chief Complaint|257,264|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|Chief Complaint|257,276|false|false|false|C0231807|Dyspnea on exertion|dyspnea on exertion
Event|Event|Chief Complaint|268,276|false|false|false|||exertion
Finding|Organism Function|Chief Complaint|268,276|false|false|false|C0015264|Exertion|exertion
Finding|Classification|Chief Complaint|280,285|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|286,294|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|286,294|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|298,316|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|307,316|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|307,316|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|307,316|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|307,316|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|307,316|false|false|false|C0184661|Interventional procedure|Procedure
Finding|Body Substance|History of Present Illness|354,361|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|354,361|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|354,361|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|371,375|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|History of Present Illness|371,375|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|History of Present Illness|376,379|false|false|false|||old
Drug|Chemical Viewed Structurally|History of Present Illness|398,405|false|false|false|C0302912|Radicals (chemistry)|radical
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|398,416|false|false|false|C0194401|Complete cystectomy|radical cystectomy
Event|Event|History of Present Illness|406,416|false|false|false|||cystectomy
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|406,416|false|false|false|C0010651|Cystectomy|cystectomy
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|428,433|false|false|false|C0020885|ileum|ileal
Disorder|Acquired Abnormality|History of Present Illness|428,441|false|false|false|C0441253|Structure of ileal conduit|ileal conduit
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|428,441|false|false|false|C0348002|Ileal conduit procedure|ileal conduit
Event|Activity|History of Present Illness|442,450|false|false|false|C1706214|Creation|creation
Event|Event|History of Present Illness|442,450|false|false|false|||creation
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|442,450|false|false|false|C0441513|Surgical construction|creation
Event|Event|History of Present Illness|464,470|false|false|false|||course
Event|Event|History of Present Illness|472,483|false|false|false|||complicated
Event|Event|History of Present Illness|487,497|false|false|false|||bacteremia
Finding|Finding|History of Present Illness|487,497|false|false|false|C0004610|Bacteremia|bacteremia
Disorder|Disease or Syndrome|History of Present Illness|502,509|false|false|false|C0000833|Abscess|abscess
Event|Event|History of Present Illness|502,509|false|false|false|||abscess
Finding|Intellectual Product|History of Present Illness|502,509|false|false|false|C1546533||abscess
Event|Event|History of Present Illness|511,514|false|false|false|||LLE
Anatomy|Body Location or Region|History of Present Illness|515,518|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|History of Present Illness|515,518|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|History of Present Illness|515,518|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|History of Present Illness|515,518|false|false|false|||DVT
Drug|Pharmacologic Substance|History of Present Illness|523,535|false|false|false|C0355642|Drugs used in migraine prophylaxis|prophylactic
Event|Event|History of Present Illness|523,535|false|false|false|||prophylactic
Finding|Functional Concept|History of Present Illness|523,535|false|false|false|C0445202|Prophylactic behavior|prophylactic
Drug|Organic Chemical|History of Present Illness|544,551|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|History of Present Illness|544,551|false|false|false|C0728963|Lovenox|lovenox
Event|Event|History of Present Illness|544,551|false|false|false|||lovenox
Event|Event|History of Present Illness|557,565|false|false|false|||presents
Event|Event|History of Present Illness|571,578|false|false|false|||dyspnea
Finding|Finding|History of Present Illness|571,578|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|History of Present Illness|571,578|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|History of Present Illness|571,590|false|false|false|C0231807|Dyspnea on exertion|dyspnea on exertion
Event|Event|History of Present Illness|582,590|false|false|false|||exertion
Finding|Organism Function|History of Present Illness|582,590|false|false|false|C0015264|Exertion|exertion
Finding|Body Substance|History of Present Illness|620,627|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|620,627|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|620,627|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|642,650|false|false|false|||admitted
Event|Occupational Activity|History of Present Illness|666,673|false|false|false|C0557854|Services|service
Finding|Idea or Concept|History of Present Illness|666,673|false|false|false|C3245478|ActInformationPrivacyReason - service|service
Disorder|Disease or Syndrome|History of Present Illness|696,704|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Event|Event|History of Present Illness|705,717|false|false|false|||exenteration
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|705,717|false|false|false|C0015258||exenteration
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|723,728|false|false|false|C0020885|ileum|ileal
Event|Event|History of Present Illness|730,737|false|false|false|||conduit
Event|Event|History of Present Illness|747,757|false|false|false|||discharged
Event|Event|History of Present Illness|761,766|false|false|false|||rehab
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|761,766|false|false|false|C0034991|Rehabilitation therapy|rehab
Drug|Pharmacologic Substance|History of Present Illness|770,782|false|false|false|C0355642|Drugs used in migraine prophylaxis|prophylactic
Event|Event|History of Present Illness|770,782|false|false|false|||prophylactic
Finding|Functional Concept|History of Present Illness|770,782|false|false|false|C0445202|Prophylactic behavior|prophylactic
Event|Event|History of Present Illness|783,789|false|false|false|||dosing
Drug|Organic Chemical|History of Present Illness|791,798|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|History of Present Illness|791,798|false|false|false|C0728963|Lovenox|lovenox
Event|Event|History of Present Illness|791,798|false|false|false|||lovenox
Finding|Idea or Concept|History of Present Illness|805,810|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|History of Present Illness|805,810|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|History of Present Illness|820,824|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|History of Present Illness|825,835|false|false|false|||readmitted
Disorder|Disease or Syndrome|History of Present Illness|850,855|false|false|false|C1258215;C4019039|Ileus;Intestinal obstruction co-occurrent and due to decreased peristalsis|ileus
Event|Event|History of Present Illness|850,855|false|false|false|||ileus
Event|Event|History of Present Illness|870,883|false|false|false|||decompression
Finding|Functional Concept|History of Present Illness|870,883|false|false|false|C1965697|Decompression - action (qualifier value)|decompression
Phenomenon|Phenomenon or Process|History of Present Illness|870,883|false|false|false|C0011117|external decompression|decompression
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|870,883|false|false|false|C0021153;C1829459|Decompression;Decompressive incision|decompression
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|885,888|false|false|false|C0027303;C1313790|NADP;TAPBP protein, human|TPN
Drug|Biologically Active Substance|History of Present Illness|885,888|false|false|false|C0027303;C1313790|NADP;TAPBP protein, human|TPN
Drug|Nucleic Acid, Nucleoside, or Nucleotide|History of Present Illness|885,888|false|false|false|C0027303;C1313790|NADP;TAPBP protein, human|TPN
Event|Event|History of Present Illness|885,888|false|false|false|||TPN
Finding|Gene or Genome|History of Present Illness|885,888|false|false|false|C1420583;C3813711|TAPBP gene;TAPBP wt Allele|TPN
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|885,888|false|false|false|C0030548|Parenteral Nutrition, Total|TPN
Event|Event|History of Present Illness|894,898|false|false|false|||grew
Disorder|Disease or Syndrome|History of Present Illness|923,926|false|false|false|C0238052|Xanthomatosis, Cerebrotendinous|CTX
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|923,926|false|false|false|C0010377;C0010583;C5574748|C-Terminal Telopeptide Type 1 Collagen, human;Crotoxin;cyclophosphamide|CTX
Drug|Biologically Active Substance|History of Present Illness|923,926|false|false|false|C0010377;C0010583;C5574748|C-Terminal Telopeptide Type 1 Collagen, human;Crotoxin;cyclophosphamide|CTX
Drug|Enzyme|History of Present Illness|923,926|false|false|false|C0010377;C0010583;C5574748|C-Terminal Telopeptide Type 1 Collagen, human;Crotoxin;cyclophosphamide|CTX
Drug|Hazardous or Poisonous Substance|History of Present Illness|923,926|false|false|false|C0010377;C0010583;C5574748|C-Terminal Telopeptide Type 1 Collagen, human;Crotoxin;cyclophosphamide|CTX
Drug|Organic Chemical|History of Present Illness|923,926|false|false|false|C0010377;C0010583;C5574748|C-Terminal Telopeptide Type 1 Collagen, human;Crotoxin;cyclophosphamide|CTX
Drug|Pharmacologic Substance|History of Present Illness|923,926|false|false|false|C0010377;C0010583;C5574748|C-Terminal Telopeptide Type 1 Collagen, human;Crotoxin;cyclophosphamide|CTX
Event|Event|History of Present Illness|923,926|false|false|false|||CTX
Finding|Gene or Genome|History of Present Illness|923,926|false|false|false|C1413864;C3539598|CYP27A1 gene;CYP27A1 wt Allele|CTX
Event|Event|History of Present Illness|931,938|false|false|false|||started
Event|Event|History of Present Illness|940,942|false|false|false|||CT
Event|Event|History of Present Illness|943,949|false|false|false|||showed
Event|Event|History of Present Illness|950,965|false|false|false|||intra-abdominal
Finding|Functional Concept|History of Present Illness|950,965|false|false|false|C1512911|Intraabdominal Route of Administration|intra-abdominal
Event|Event|History of Present Illness|967,976|false|false|false|||interloop
Finding|Gene or Genome|History of Present Illness|979,985|false|false|false|C1424587|LITAF gene|simple
Drug|Substance|History of Present Illness|986,991|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|History of Present Illness|986,991|false|false|false|||fluid
Finding|Intellectual Product|History of Present Illness|986,991|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|History of Present Illness|992,1002|false|false|false|||collection
Finding|Conceptual Entity|History of Present Illness|992,1002|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|History of Present Illness|992,1002|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|History of Present Illness|992,1002|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|History of Present Illness|992,1002|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Anatomy|Body Location or Region|History of Present Illness|1007,1010|false|false|false|C0230180|Structure of left lower quadrant of abdomen|LLQ
Drug|Substance|History of Present Illness|1011,1016|false|false|false|C1550628|Drain - SpecimenType|drain
Event|Event|History of Present Illness|1011,1016|false|false|false|||drain
Finding|Intellectual Product|History of Present Illness|1011,1016|false|false|false|C1546604|Drain Specimen Code|drain
Event|Event|History of Present Illness|1021,1027|false|false|false|||placed
Finding|Body Substance|History of Present Illness|1036,1043|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|1036,1043|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|1036,1043|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|History of Present Illness|1045,1053|false|false|false|||improved
Disorder|Disease or Syndrome|History of Present Illness|1063,1066|false|false|false|C0006430|Burning Mouth Syndrome|BMs
Event|Event|History of Present Illness|1063,1066|false|false|false|||BMs
Event|Event|History of Present Illness|1094,1104|false|false|false|||discharged
Drug|Organic Chemical|History of Present Illness|1109,1114|false|false|false|C0701042|Cipro|cipro
Drug|Pharmacologic Substance|History of Present Illness|1109,1114|false|false|false|C0701042|Cipro|cipro
Event|Event|History of Present Illness|1109,1114|false|false|false|||cipro
Drug|Organic Chemical|History of Present Illness|1115,1121|false|false|false|C0699678|Flagyl|flagyl
Drug|Pharmacologic Substance|History of Present Illness|1115,1121|false|false|false|C0699678|Flagyl|flagyl
Event|Event|History of Present Illness|1115,1121|false|false|false|||flagyl
Event|Event|History of Present Illness|1136,1146|false|false|false|||discharged
Drug|Organic Chemical|History of Present Illness|1153,1160|false|false|false|C0591139|Bactrim|Bactrim
Drug|Pharmacologic Substance|History of Present Illness|1153,1160|false|false|false|C0591139|Bactrim|Bactrim
Event|Event|History of Present Illness|1153,1160|false|false|false|||Bactrim
Event|Event|History of Present Illness|1165,1173|false|false|false|||presumed
Disorder|Disease or Syndrome|History of Present Illness|1175,1178|false|false|false|C0042029|Urinary tract infection|UTI
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1175,1178|false|false|false|C0077906|urinastatin|UTI
Drug|Pharmacologic Substance|History of Present Illness|1175,1178|false|false|false|C0077906|urinastatin|UTI
Event|Event|History of Present Illness|1175,1178|false|false|false|||UTI
Finding|Gene or Genome|History of Present Illness|1175,1178|false|false|false|C1412376;C5780748|AMBP gene;AMBP wt Allele|UTI
Event|Event|History of Present Illness|1211,1215|false|false|false|||took
Event|Event|History of Present Illness|1235,1244|false|false|false|||admission
Procedure|Health Care Activity|History of Present Illness|1235,1244|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|History of Present Illness|1254,1259|false|false|false|||noted
Finding|Finding|History of Present Illness|1268,1271|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|History of Present Illness|1268,1271|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Attribute|Clinical Attribute|History of Present Illness|1286,1291|false|false|false|C1717255||edema
Event|Event|History of Present Illness|1286,1291|false|false|false|||edema
Finding|Pathologic Function|History of Present Illness|1286,1291|false|false|false|C0013604|Edema|edema
Finding|Finding|History of Present Illness|1307,1311|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|History of Present Illness|1307,1311|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|History of Present Illness|1307,1311|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|History of Present Illness|1312,1318|false|false|false|||showed
Attribute|Clinical Attribute|History of Present Illness|1324,1328|false|false|false|C4318566|Deep Resection Margin|deep
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1324,1333|false|false|false|C0226514|Structure of deep vein|deep vein
Disorder|Disease or Syndrome|History of Present Illness|1324,1344|false|false|false|C0149871;C0340708|Deep Vein Thrombosis;Deep vein thrombosis of lower limb|deep vein thrombosis
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1329,1333|false|false|false|C0042449|Veins|vein
Finding|Pathologic Function|History of Present Illness|1329,1344|false|false|false|C0042487|Venous Thrombosis|vein thrombosis
Event|Event|History of Present Illness|1334,1344|false|false|false|||thrombosis
Finding|Pathologic Function|History of Present Illness|1334,1344|false|false|false|C0040053|Thrombosis|thrombosis
Event|Event|History of Present Illness|1352,1362|false|false|false|||duplicated
Finding|Finding|History of Present Illness|1352,1362|false|false|false|C0332597|Duplication (finding)|duplicated
Attribute|Clinical Attribute|History of Present Illness|1372,1378|false|false|false|C4522154|Distal Resection Margin|distal
Finding|Functional Concept|History of Present Illness|1379,1383|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1384,1391|false|false|false|C0015811|Femur|femoral
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1384,1397|false|false|false|C0015809|Femoral vein|femoral veins
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1392,1397|false|false|false|C0042449|Veins|veins
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1392,1397|false|false|false|C0398102|Procedure on vein|veins
Event|Event|History of Present Illness|1407,1417|false|false|false|||discharged
Drug|Organic Chemical|History of Present Illness|1423,1433|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Pharmacologic Substance|History of Present Illness|1423,1433|false|false|false|C0206460|enoxaparin|Enoxaparin
Event|Event|History of Present Illness|1423,1433|false|false|false|||Enoxaparin
Drug|Organic Chemical|History of Present Illness|1423,1440|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Pharmacologic Substance|History of Present Illness|1423,1440|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Biologically Active Substance|History of Present Illness|1434,1440|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|History of Present Illness|1434,1440|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|History of Present Illness|1434,1440|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|History of Present Illness|1434,1440|false|false|false|||Sodium
Finding|Physiologic Function|History of Present Illness|1434,1440|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|History of Present Illness|1434,1440|false|false|false|C0337443|Sodium measurement|Sodium
Event|Event|History of Present Illness|1461,1468|false|false|false|||reports
Disorder|Disease or Syndrome|History of Present Illness|1478,1481|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|1478,1481|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|History of Present Illness|1478,1481|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1478,1481|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|History of Present Illness|1478,1481|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|History of Present Illness|1478,1481|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|History of Present Illness|1478,1481|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|History of Present Illness|1478,1481|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|History of Present Illness|1478,1481|false|false|false|||PCP
Finding|Gene or Genome|History of Present Illness|1478,1481|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|History of Present Illness|1478,1481|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|History of Present Illness|1483,1490|false|false|false|||started
Finding|Intellectual Product|History of Present Illness|1519,1523|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|History of Present Illness|1540,1551|false|false|false|||improvement
Finding|Conceptual Entity|History of Present Illness|1540,1551|false|false|false|C2986411|Improvement|improvement
Event|Event|History of Present Illness|1559,1567|false|false|false|||swelling
Finding|Finding|History of Present Illness|1559,1567|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|History of Present Illness|1559,1567|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Attribute|Clinical Attribute|History of Present Illness|1577,1583|false|false|false|C4255046||report
Event|Event|History of Present Illness|1577,1583|false|false|false|||report
Finding|Intellectual Product|History of Present Illness|1577,1583|false|false|false|C0684224|Report (document)|report
Procedure|Health Care Activity|History of Present Illness|1577,1583|false|false|false|C0700287|Reporting|report
Finding|Functional Concept|History of Present Illness|1587,1593|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1606,1611|false|false|false|C0034991|Rehabilitation therapy|rehab
Event|Event|History of Present Illness|1612,1620|false|false|false|||facility
Finding|Intellectual Product|History of Present Illness|1612,1620|false|false|false|C4695111|ADMIN.FACILITY|facility
Event|Event|History of Present Illness|1631,1639|false|false|false|||negative
Finding|Classification|History of Present Illness|1631,1639|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|History of Present Illness|1631,1639|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|History of Present Illness|1631,1639|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|History of Present Illness|1631,1643|false|false|false|C0205160|Negative|negative for
Anatomy|Body Location or Region|History of Present Illness|1644,1647|true|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|History of Present Illness|1644,1647|true|false|false|C2926618||DVT
Disorder|Disease or Syndrome|History of Present Illness|1644,1647|true|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|History of Present Illness|1644,1647|true|false|false|||DVT
Finding|Body Substance|History of Present Illness|1650,1657|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|1650,1657|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|1650,1657|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|History of Present Illness|1658,1665|false|false|false|||reports
Event|Event|History of Present Illness|1675,1684|false|false|false|||recovered
Finding|Finding|History of Present Illness|1685,1689|false|false|false|C5575035|Well (answer to question)|well
Event|Event|History of Present Illness|1722,1726|false|false|false|||well
Finding|Finding|History of Present Illness|1722,1726|false|false|false|C5575035|Well (answer to question)|well
Procedure|Health Care Activity|History of Present Illness|1734,1749|false|false|false|C1456630|Assisted Living|assisted living
Event|Event|History of Present Illness|1743,1749|false|false|false|||living
Finding|Conceptual Entity|History of Present Illness|1743,1749|false|false|false|C0595998;C4520849;C4551704|Alive;Household composition;Living|living
Finding|Finding|History of Present Illness|1743,1749|false|false|false|C0595998;C4520849;C4551704|Alive;Household composition;Living|living
Finding|Intellectual Product|History of Present Illness|1750,1758|false|false|false|C4695111|ADMIN.FACILITY|facility
Finding|Intellectual Product|History of Present Illness|1770,1774|false|false|false|C1561540|Transaction counts and value totals - week|week
Finding|Gene or Genome|History of Present Illness|1775,1778|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|History of Present Illness|1789,1794|false|false|false|||began
Event|Event|History of Present Illness|1808,1815|false|false|false|||dyspnea
Finding|Finding|History of Present Illness|1808,1815|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|History of Present Illness|1808,1815|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|History of Present Illness|1808,1827|false|false|false|C0231807|Dyspnea on exertion|dyspnea on exertion
Event|Event|History of Present Illness|1819,1827|false|false|false|||exertion
Finding|Organism Function|History of Present Illness|1819,1827|false|false|false|C0015264|Exertion|exertion
Event|Event|History of Present Illness|1833,1839|false|false|false|||states
Event|Event|History of Present Illness|1863,1867|false|false|false|||able
Finding|Finding|History of Present Illness|1863,1867|false|false|false|C1299581|Able (qualifier value)|able
Event|Event|History of Present Illness|1871,1879|false|false|false|||ambulate
Drug|Biomedical or Dental Material|History of Present Illness|1882,1887|false|false|false|C1706085|Block Dosage Form|block
Event|Event|History of Present Illness|1882,1887|false|false|false|||block
Finding|Body Substance|History of Present Illness|1882,1887|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|block
Finding|Finding|History of Present Illness|1882,1887|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|block
Finding|Functional Concept|History of Present Illness|1882,1887|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|block
Event|Event|History of Present Illness|1895,1903|false|false|false|||stopping
Event|Event|History of Present Illness|1908,1913|false|false|false|||catch
Finding|Sign or Symptom|History of Present Illness|1908,1913|false|false|false|C0231617|Catch - Finding of sensory dimension of pain|catch
Event|Event|History of Present Illness|1918,1924|false|false|false|||breath
Finding|Body Substance|History of Present Illness|1918,1924|false|false|false|C0225386|Breath|breath
Finding|Intellectual Product|History of Present Illness|1946,1950|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|History of Present Illness|1964,1970|false|false|false|||unable
Finding|Finding|History of Present Illness|1964,1970|false|false|false|C1299582|Unable|unable
Event|Event|History of Present Illness|1996,2001|false|false|false|||steps
Finding|Conceptual Entity|History of Present Illness|1996,2001|false|false|false|C1261552|Step (specific stage)|steps
Procedure|Health Care Activity|History of Present Illness|1996,2001|false|false|false|C4722257|STEPS to Enhance Physical Activity|steps
Event|Event|History of Present Illness|2007,2013|false|false|false|||states
Event|Event|History of Present Illness|2026,2032|false|false|false|||become
Event|Event|History of Present Illness|2052,2061|false|false|false|||difficult
Finding|Finding|History of Present Illness|2052,2061|false|false|false|C0332218|Difficult (qualifier value)|difficult
Event|Event|History of Present Illness|2065,2073|false|false|false|||ambulate
Event|Event|History of Present Illness|2083,2090|false|false|false|||bedroom
Event|Event|History of Present Illness|2099,2107|false|false|false|||bathroom
Event|Event|History of Present Illness|2114,2121|false|false|false|||visited
Finding|Functional Concept|History of Present Illness|2136,2146|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|ambulatory
Finding|Idea or Concept|History of Present Illness|2136,2146|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|ambulatory
Finding|Intellectual Product|History of Present Illness|2136,2146|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|ambulatory
Procedure|Health Care Activity|History of Present Illness|2136,2146|false|false|false|C1561560|ambulatory encounter|ambulatory
Event|Event|History of Present Illness|2147,2157|false|false|false|||saturation
Phenomenon|Natural Phenomenon or Process|History of Present Illness|2147,2157|false|false|false|C0522534|Saturated|saturation
Event|Event|History of Present Illness|2163,2168|false|false|false|||noted
Event|Event|History of Present Illness|2202,2213|false|false|false|||tachycardia
Finding|Finding|History of Present Illness|2202,2213|false|false|false|C0039231;C3827868|Tachycardia;Tachycardia by ECG Finding|tachycardia
Event|Event|History of Present Illness|2223,2229|false|false|false|||pallor
Finding|Finding|History of Present Illness|2223,2229|false|false|false|C0241137|Pallor of skin|pallor
Event|Event|History of Present Illness|2234,2245|false|false|false|||diaphoresis
Finding|Finding|History of Present Illness|2234,2245|false|false|false|C0700590|Increased sweating|diaphoresis
Event|Event|History of Present Illness|2251,2259|false|false|false|||endorses
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2271,2274|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Pathologic Function|History of Present Illness|2271,2283|false|true|false|C0581394|Swelling of lower limb|leg swelling
Event|Event|History of Present Illness|2275,2283|false|false|false|||swelling
Finding|Finding|History of Present Illness|2275,2283|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|History of Present Illness|2275,2283|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Functional Concept|History of Present Illness|2285,2289|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Event|Event|History of Present Illness|2290,2295|false|false|false|||worse
Finding|Finding|History of Present Illness|2290,2295|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Idea or Concept|History of Present Illness|2290,2295|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Event|Event|History of Present Illness|2301,2306|false|false|false|||right
Finding|Functional Concept|History of Present Illness|2301,2306|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Event|Event|History of Present Illness|2316,2322|false|false|false|||states
Anatomy|Body Location or Region|History of Present Illness|2332,2338|false|false|false|C0039866|Thigh structure|thighs
Event|Event|History of Present Illness|2340,2344|false|false|false|||feel
Finding|Mental Process|History of Present Illness|2340,2344|false|false|false|C1527305|Feelings|feel
Event|Event|History of Present Illness|2358,2364|true|false|false|||denies
Anatomy|Body Location or Region|History of Present Illness|2380,2385|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|2380,2385|true|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|2380,2390|true|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|2380,2390|true|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|2386,2390|true|false|false|C2598155||pain
Event|Event|History of Present Illness|2386,2390|true|false|false|||pain
Finding|Functional Concept|History of Present Illness|2386,2390|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|2386,2390|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|2392,2397|true|false|false|||fever
Finding|Finding|History of Present Illness|2392,2397|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|History of Present Illness|2392,2397|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|History of Present Illness|2399,2405|true|false|false|||chills
Finding|Sign or Symptom|History of Present Illness|2399,2405|true|false|false|C0085593|Chills|chills
Attribute|Clinical Attribute|History of Present Illness|2408,2412|false|false|false|C2598155||pain
Event|Event|History of Present Illness|2408,2412|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|2408,2412|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|2408,2412|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|History of Present Illness|2418,2422|false|false|false|C4318566|Deep Resection Margin|deep
Event|Event|History of Present Illness|2423,2434|false|false|false|||inspiration
Finding|Organism Function|History of Present Illness|2423,2434|false|false|false|C0004048|Inspiration (function)|inspiration
Anatomy|Body Location or Region|History of Present Illness|2436,2445|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|History of Present Illness|2436,2450|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|History of Present Illness|2446,2450|false|false|false|C2598155||pain
Event|Event|History of Present Illness|2446,2450|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|2446,2450|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|2446,2450|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|2452,2458|false|false|false|||rashes
Finding|Sign or Symptom|History of Present Illness|2452,2458|false|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Event|Event|History of Present Illness|2460,2469|false|false|false|||dizziness
Finding|Sign or Symptom|History of Present Illness|2460,2469|false|false|false|C0012833;C0042571|Dizziness;Vertigo|dizziness
Event|Event|History of Present Illness|2472,2487|false|false|false|||lightheadedness
Finding|Sign or Symptom|History of Present Illness|2472,2487|false|false|false|C0220870|Lightheadedness|lightheadedness
Finding|Idea or Concept|History of Present Illness|2503,2510|false|false|false|C1555582|Initial (abbreviation)|initial
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2543,2548|false|false|false|C0028429||Nasal
Drug|Biomedical or Dental Material|History of Present Illness|2543,2548|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Organic Chemical|History of Present Illness|2543,2548|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Pharmacologic Substance|History of Present Illness|2543,2548|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Finding|Finding|History of Present Illness|2543,2548|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Functional Concept|History of Present Illness|2543,2548|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2549,2556|false|false|false|C1550232|Body Parts - Cannula|Cannula
Finding|Body Substance|History of Present Illness|2549,2556|false|false|false|C1546577;C1550622|Specimen Type - Cannula|Cannula
Finding|Intellectual Product|History of Present Illness|2549,2556|false|false|false|C1546577;C1550622|Specimen Type - Cannula|Cannula
Event|Event|History of Present Illness|2562,2570|false|false|false|||physical
Finding|Finding|History of Present Illness|2562,2570|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Finding|Functional Concept|History of Present Illness|2562,2570|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Procedure|Health Care Activity|History of Present Illness|2562,2570|false|false|false|C0031809|Physical Examination|physical
Finding|Finding|History of Present Illness|2562,2575|false|false|false|C1509143|physical examination (physical finding)|physical exam
Procedure|Health Care Activity|History of Present Illness|2562,2575|false|false|false|C0031809|Physical Examination|physical exam
Event|Event|History of Present Illness|2571,2575|false|false|false|||exam
Finding|Functional Concept|History of Present Illness|2571,2575|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|History of Present Illness|2571,2575|false|false|false|C0582103|Medical Examination|exam
Event|Event|History of Present Illness|2580,2588|false|false|false|||recorded
Finding|Body Substance|History of Present Illness|2592,2599|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|2592,2599|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|2592,2599|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2637,2640|false|false|false|C0023759|Lip structure|lip
Disorder|Disease or Syndrome|History of Present Illness|2637,2640|false|false|false|C0153932;C0264511|Benign neoplasm of the lip;Lymphoid interstitial pneumonia|lip
Disorder|Neoplastic Process|History of Present Illness|2637,2640|false|false|false|C0153932;C0264511|Benign neoplasm of the lip;Lymphoid interstitial pneumonia|lip
Finding|Gene or Genome|History of Present Illness|2637,2640|false|false|false|C1846919;C3889123|SMG1 gene;SMG1 wt Allele|lip
Attribute|Clinical Attribute|History of Present Illness|2641,2650|false|false|false|C5885990||breathing
Event|Event|History of Present Illness|2641,2650|false|false|false|||breathing
Finding|Finding|History of Present Illness|2641,2650|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|History of Present Illness|2641,2650|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|History of Present Illness|2641,2650|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|History of Present Illness|2641,2650|false|false|false|C1160636|respiratory system process|breathing
Event|Event|History of Present Illness|2652,2658|false|false|false|||unable
Finding|Finding|History of Present Illness|2652,2658|false|false|false|C1299582|Unable|unable
Finding|Finding|History of Present Illness|2652,2667|false|false|false|C0564216;C4722246|Unable to Speak at All;Unable to speak (finding)|unable to speak
Event|Event|History of Present Illness|2662,2667|false|false|false|||speak
Finding|Finding|History of Present Illness|2662,2667|false|false|false|C0234856;C0600116;C1547187|Does speak;Speak - language ability;Speaking (function)|speak
Finding|Idea or Concept|History of Present Illness|2662,2667|false|false|false|C0234856;C0600116;C1547187|Does speak;Speak - language ability;Speaking (function)|speak
Finding|Individual Behavior|History of Present Illness|2662,2667|false|false|false|C0234856;C0600116;C1547187|Does speak;Speak - language ability;Speaking (function)|speak
Event|Event|History of Present Illness|2676,2685|false|false|false|||sentences
Finding|Intellectual Product|History of Present Illness|2676,2685|false|false|false|C0876929|Sentence|sentences
Event|Event|History of Present Illness|2694,2702|false|false|false|||becoming
Finding|Sign or Symptom|History of Present Illness|2703,2718|false|false|false|C0013404|Dyspnea|short of breath
Finding|Body Substance|History of Present Illness|2712,2718|false|false|false|C0225386|Breath|breath
Anatomy|Anatomical Structure|History of Present Illness|2720,2728|false|false|false|C0559495|Urological stoma|urostomy
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|2720,2728|false|false|false|C0856443|Urostomy procedure|urostomy
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2729,2734|false|false|false|C0222017|Abdominal skin pouch|pouch
Anatomy|Body Location or Region|History of Present Illness|2738,2741|false|false|false|C0230178|Structure of right lower quadrant of abdomen|RLQ
Anatomy|Anatomical Structure|History of Present Illness|2743,2748|false|false|false|C1955856|Surgical Stoma|stoma
Attribute|Clinical Attribute|History of Present Illness|2759,2764|false|false|false|C1717255||edema
Event|Event|History of Present Illness|2759,2764|false|false|false|||edema
Finding|Pathologic Function|History of Present Illness|2759,2764|false|false|false|C0013604|Edema|edema
Anatomy|Body Location or Region|History of Present Illness|2778,2783|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|History of Present Illness|2778,2783|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2778,2795|false|false|false|C0023216|Lower Extremity|lower extremities
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2784,2795|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Event|Event|History of Present Illness|2806,2810|false|false|false|||labs
Lab|Laboratory or Test Result|History of Present Illness|2806,2810|false|false|false|C0587081|Laboratory test finding|labs
Event|Event|History of Present Illness|2816,2823|false|false|false|||notable
Event|Event|History of Present Illness|2835,2838|false|false|false|||Hct
Procedure|Laboratory Procedure|History of Present Illness|2835,2838|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|2835,2838|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Event|Event|History of Present Illness|2843,2846|false|false|false|||plt
Procedure|Laboratory Procedure|History of Present Illness|2843,2846|false|false|false|C0201617|Primed lymphocyte test|plt
Finding|Gene or Genome|History of Present Illness|2856,2861|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Anatomy|Cell|History of Present Illness|2873,2876|false|false|false|C0023516|Leukocytes|WBC
Disorder|Disease or Syndrome|History of Present Illness|2890,2893|false|false|false|C0267963|Exocrine pancreatic insufficiency|epi
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|2890,2893|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|epi
Drug|Biologically Active Substance|History of Present Illness|2890,2893|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|epi
Drug|Hormone|History of Present Illness|2890,2893|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|epi
Drug|Organic Chemical|History of Present Illness|2890,2893|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|epi
Drug|Pharmacologic Substance|History of Present Illness|2890,2893|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|epi
Event|Event|History of Present Illness|2890,2893|false|false|false|||epi
Finding|Gene or Genome|History of Present Illness|2890,2893|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|epi
Finding|Intellectual Product|History of Present Illness|2890,2893|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|epi
Procedure|Diagnostic Procedure|History of Present Illness|2890,2893|false|false|false|C0162734;C3641909|Echo-Planar Imaging;Electronic Portal Imaging|epi
Finding|Finding|History of Present Illness|2900,2903|false|false|false|C5848551|Neg - answer|neg
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|2908,2914|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Drug|Hormone|History of Present Illness|2908,2914|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Event|Event|History of Present Illness|2915,2921|false|false|false|||normal
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|2923,2926|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|History of Present Illness|2923,2926|false|false|false|||CTA
Finding|Gene or Genome|History of Present Illness|2923,2926|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|History of Present Illness|2923,2926|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Anatomy|Body Location or Region|History of Present Illness|2927,2932|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|2927,2932|false|false|false|C0741025|Chest problem|chest
Event|Event|History of Present Illness|2933,2939|false|false|false|||showed
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2954,2963|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|History of Present Illness|2954,2963|false|false|false|C2707265||pulmonary
Finding|Finding|History of Present Illness|2954,2963|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|History of Present Illness|2954,2972|false|false|false|C0034065|Pulmonary Embolism|pulmonary embolism
Event|Event|History of Present Illness|2964,2972|false|false|false|||embolism
Finding|Finding|History of Present Illness|2964,2972|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Finding|Pathologic Function|History of Present Illness|2964,2972|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Event|Event|History of Present Illness|2978,2986|false|false|false|||thrombus
Finding|Pathologic Function|History of Present Illness|2978,2986|false|false|false|C0087086;C0302148|Blood Clot;Thrombus|thrombus
Event|Event|History of Present Illness|2987,2991|false|false|false|||seen
Event|Event|History of Present Illness|2992,3001|false|false|false|||extending
Finding|Functional Concept|History of Present Illness|3012,3017|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|3012,3039|false|false|false|C0226054;C0923924|Right pulmonary arterial tree;Right pulmonary artery|right main pulmonary artery
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|3023,3032|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|History of Present Illness|3023,3032|false|false|false|C2707265||pulmonary
Finding|Finding|History of Present Illness|3023,3032|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|3023,3039|false|false|false|C0034052|Pulmonary artery structure|pulmonary artery
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|3033,3039|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|History of Present Illness|3033,3039|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Finding|Functional Concept|History of Present Illness|3077,3082|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Event|Event|History of Present Illness|3090,3096|false|false|false|||middle
Finding|Intellectual Product|History of Present Illness|3090,3096|false|false|false|C1552826|Table Cell Vertical Align - middle|middle
Anatomy|Body Location or Region|History of Present Illness|3102,3107|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|History of Present Illness|3102,3107|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|3102,3112|false|false|false|C0225758|Structure of lower lobe of lung|lower lobe
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|3108,3112|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|History of Present Illness|3108,3112|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|3108,3122|false|false|false|C0225752|Structure of lobe of lung|lobe pulmonary
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|3113,3122|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|History of Present Illness|3113,3122|false|false|false|C2707265||pulmonary
Finding|Finding|History of Present Illness|3113,3122|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|3124,3132|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Anatomy|Body System|History of Present Illness|3124,3132|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Event|Event|History of Present Illness|3124,3132|false|false|false|||arteries
Procedure|Health Care Activity|History of Present Illness|3124,3132|false|false|false|C0397581|Procedure on artery|arteries
Finding|Functional Concept|History of Present Illness|3137,3142|true|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|History of Present Illness|3137,3148|true|false|false|C0225808|Right side of heart|right heart
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|3143,3148|true|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|History of Present Illness|3143,3148|true|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|History of Present Illness|3143,3148|true|false|false|C0795691|HEART PROBLEM|heart
Disorder|Injury or Poisoning|History of Present Illness|3149,3155|true|false|false|C0080194|Muscle strain|strain
Event|Event|History of Present Illness|3149,3155|true|false|false|||strain
Finding|Idea or Concept|History of Present Illness|3149,3155|true|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Finding|Mental Process|History of Present Illness|3149,3155|true|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Finding|Physiologic Function|History of Present Illness|3149,3155|true|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Finding|Sign or Symptom|History of Present Illness|3149,3155|true|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Event|Event|History of Present Illness|3156,3166|true|false|false|||identified
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|3204,3213|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|History of Present Illness|3204,3213|false|false|false|C2707265||pulmonary
Finding|Finding|History of Present Illness|3204,3213|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|History of Present Illness|3204,3220|false|false|false|C0034065|Pulmonary Embolism|pulmonary emboli
Event|Event|History of Present Illness|3214,3220|false|false|false|||emboli
Finding|Finding|History of Present Illness|3214,3220|false|false|false|C1704212|Embolus|emboli
Event|Event|History of Present Illness|3221,3225|false|false|false|||seen
Event|Event|History of Present Illness|3261,3269|false|false|false|||branches
Finding|Functional Concept|History of Present Illness|3277,3281|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|History of Present Illness|3292,3297|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|History of Present Illness|3292,3297|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|3298,3303|false|false|false|C0796494|lobe|lobes
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|3317,3326|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|History of Present Illness|3317,3326|false|false|false|C2707265||pulmonary
Finding|Finding|History of Present Illness|3317,3326|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Finding|History of Present Illness|3317,3334|false|false|false|C0748164|Multiple Pulmonary Nodules|pulmonary nodules
Event|Event|History of Present Illness|3327,3334|false|false|false|||nodules
Event|Event|History of Present Illness|3339,3344|false|false|false|||noted
Event|Event|History of Present Illness|3349,3354|false|false|false|||noted
Event|Event|History of Present Illness|3395,3405|false|false|false|||spiculated
Event|Event|History of Present Illness|3410,3419|false|false|false|||measuring
Finding|Functional Concept|History of Present Illness|3439,3444|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|3439,3456|false|false|false|C4281590|Structure of middle lobe of right lung|right middle lobe
Finding|Intellectual Product|History of Present Illness|3445,3451|false|false|false|C1552826|Table Cell Vertical Align - middle|middle
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|3445,3456|false|false|false|C4281590|Structure of middle lobe of right lung|middle lobe
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|3452,3456|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|History of Present Illness|3452,3456|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Event|Event|History of Present Illness|3458,3468|false|false|false|||suspicious
Finding|Finding|History of Present Illness|3458,3483|false|false|false|C4050405|Suspicious for Malignancy|suspicious for malignancy
Disorder|Neoplastic Process|History of Present Illness|3473,3483|false|true|false|C0006826;C1306459|Malignant Neoplasms;Primary malignant neoplasm|malignancy
Event|Event|History of Present Illness|3473,3483|false|false|false|||malignancy
Procedure|Diagnostic Procedure|History of Present Illness|3501,3504|false|false|false|C0032743;C0040398|Positron-Emission Tomography;Tomography, Emission-Computed|PET
Procedure|Diagnostic Procedure|History of Present Illness|3501,3507|false|false|false|C1699633|PET/CT scan|PET-CT
Event|Event|History of Present Illness|3505,3507|false|false|false|||CT
Event|Event|History of Present Illness|3516,3529|false|false|false|||demonstration
Finding|Functional Concept|History of Present Illness|3535,3539|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|3535,3546|false|false|false|C0222601|Left breast|left breast
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|3540,3546|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|History of Present Illness|3540,3546|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Finding|Finding|History of Present Illness|3540,3546|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|3540,3546|false|false|false|C0191838|Procedures on breast|breast
Finding|Finding|History of Present Illness|3540,3554|false|false|false|C0024103|Mass in breast|breast nodules
Event|Event|History of Present Illness|3547,3554|false|false|false|||nodules
Event|Event|History of Present Illness|3566,3577|false|false|false|||correlation
Event|Event|History of Present Illness|3583,3594|false|false|false|||mammography
Procedure|Diagnostic Procedure|History of Present Illness|3583,3594|false|false|false|C0024671;C0848600|Mammography;Mammography, Female|mammography
Event|Event|History of Present Illness|3599,3609|false|false|false|||ultrasound
Finding|Functional Concept|History of Present Illness|3599,3609|false|false|false|C0220934|Ultrasonic|ultrasound
Phenomenon|Natural Phenomenon or Process|History of Present Illness|3599,3609|false|false|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|ultrasound
Procedure|Diagnostic Procedure|History of Present Illness|3599,3609|false|false|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|ultrasound
Event|Event|History of Present Illness|3613,3622|false|false|false|||suggested
Event|Event|History of Present Illness|3625,3628|false|false|false|||EKG
Finding|Intellectual Product|History of Present Illness|3625,3628|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|History of Present Illness|3625,3628|false|false|false|C1623258|Electrocardiography|EKG
Event|Event|History of Present Illness|3629,3635|false|false|false|||showed
Event|Event|History of Present Illness|3636,3639|false|false|false|||NSR
Finding|Molecular Function|History of Present Illness|3636,3639|false|false|false|C1704493;C2700623|Neutral Sidebent Rotated|NSR
Finding|Pathologic Function|History of Present Illness|3636,3639|false|false|false|C1704493;C2700623|Neutral Sidebent Rotated|NSR
Anatomy|Cell Component|History of Present Illness|3654,3657|false|false|false|C5239889|protein aggregate center|PAC
Disorder|Disease or Syndrome|History of Present Illness|3654,3657|false|false|false|C0033036|Atrial Premature Complexes|PAC
Event|Event|History of Present Illness|3654,3657|false|false|false|||PAC
Finding|Finding|History of Present Illness|3654,3657|false|false|false|C1823219;C4082832|Atrial Premature Complex by ECG Finding;PACC1 gene|PAC
Finding|Gene or Genome|History of Present Illness|3654,3657|false|false|false|C1823219;C4082832|Atrial Premature Complex by ECG Finding;PACC1 gene|PAC
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|3654,3657|false|false|false|C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol|PAC
Finding|Body Substance|History of Present Illness|3659,3666|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|3659,3666|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|3659,3666|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Organic Chemical|History of Present Illness|3694,3707|false|false|false|C0008809|ciprofloxacin|Ciprofloxacin
Drug|Pharmacologic Substance|History of Present Illness|3694,3707|false|false|false|C0008809|ciprofloxacin|Ciprofloxacin
Drug|Antibiotic|History of Present Illness|3694,3711|false|false|false|C0282104|ciprofloxacin hydrochloride|Ciprofloxacin HCl
Drug|Organic Chemical|History of Present Illness|3694,3711|false|false|false|C0282104|ciprofloxacin hydrochloride|Ciprofloxacin HCl
Disorder|Neoplastic Process|History of Present Illness|3708,3711|false|false|false|C0023443|Hairy Cell Leukemia|HCl
Drug|Immunologic Factor|History of Present Illness|3708,3711|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Inorganic Chemical|History of Present Illness|3708,3711|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Pharmacologic Substance|History of Present Illness|3708,3711|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Event|Event|History of Present Illness|3708,3711|false|false|false|||HCl
Drug|Biologically Active Substance|History of Present Illness|3733,3740|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Drug|Organic Chemical|History of Present Illness|3733,3740|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Drug|Pharmacologic Substance|History of Present Illness|3733,3740|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Event|Event|History of Present Illness|3733,3740|false|false|false|||Heparin
Event|Event|History of Present Illness|3746,3750|false|false|false|||UNIT
Drug|Biologically Active Substance|History of Present Illness|3765,3772|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Drug|Organic Chemical|History of Present Illness|3765,3772|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Drug|Pharmacologic Substance|History of Present Illness|3765,3772|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Event|Event|History of Present Illness|3765,3772|false|false|false|||Heparin
Event|Event|History of Present Illness|3776,3784|false|false|false|||Transfer
Finding|Functional Concept|History of Present Illness|3776,3784|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|Transfer
Finding|Idea or Concept|History of Present Illness|3776,3784|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|Transfer
Procedure|Health Care Activity|History of Present Illness|3776,3784|false|false|false|C4706767|Transfer (immobility management)|Transfer
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|3816,3821|false|false|false|C0028429||Nasal
Drug|Biomedical or Dental Material|History of Present Illness|3816,3821|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Organic Chemical|History of Present Illness|3816,3821|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Pharmacologic Substance|History of Present Illness|3816,3821|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Finding|Finding|History of Present Illness|3816,3821|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Functional Concept|History of Present Illness|3816,3821|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|3822,3829|false|false|false|C1550232|Body Parts - Cannula|Cannula
Finding|Body Substance|History of Present Illness|3822,3829|false|false|false|C1546577;C1550622|Specimen Type - Cannula|Cannula
Finding|Intellectual Product|History of Present Illness|3822,3829|false|false|false|C1546577;C1550622|Specimen Type - Cannula|Cannula
Event|Event|History of Present Illness|3837,3841|false|false|false|||seen
Anatomy|Anatomical Structure|History of Present Illness|3849,3854|false|false|false|C3714591|Floor (anatomic)|floor
Event|Event|History of Present Illness|3860,3867|false|false|false|||reports
Finding|Idea or Concept|History of Present Illness|3868,3879|false|false|false|C0750502|Significant|significant
Event|Event|History of Present Illness|3880,3887|false|false|false|||dyspnea
Finding|Finding|History of Present Illness|3880,3887|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|History of Present Illness|3880,3887|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Event|Event|History of Present Illness|3902,3910|false|false|false|||exertion
Finding|Organism Function|History of Present Illness|3902,3910|false|false|false|C0015264|Exertion|exertion
Event|Event|History of Present Illness|3912,3918|false|false|false|||Denies
Anatomy|Body Location or Region|History of Present Illness|3919,3924|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|3919,3924|true|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|3919,3929|true|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|3919,3929|true|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|3925,3929|true|false|false|C2598155||pain
Event|Event|History of Present Illness|3925,3929|true|false|false|||pain
Finding|Functional Concept|History of Present Illness|3925,3929|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|3925,3929|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|3931,3943|true|false|false|||palpitations
Finding|Finding|History of Present Illness|3931,3943|true|false|false|C0030252|Palpitations|palpitations
Event|Event|History of Present Illness|3946,3961|true|false|false|||lightheadedness
Finding|Sign or Symptom|History of Present Illness|3946,3961|true|false|false|C0220870|Lightheadedness|lightheadedness
Anatomy|Body Space or Junction|History of Present Illness|3975,3978|false|false|false|C0262327|rostral sulcus|ROS
Drug|Biologically Active Substance|History of Present Illness|3975,3978|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Element, Ion, or Isotope|History of Present Illness|3975,3978|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Organic Chemical|History of Present Illness|3975,3978|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Pharmacologic Substance|History of Present Illness|3975,3978|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Event|Event|History of Present Illness|3975,3978|false|false|false|||ROS
Finding|Gene or Genome|History of Present Illness|3975,3978|false|false|false|C0812281;C1709820|ROS1 gene;ROS1 wt Allele|ROS
Procedure|Health Care Activity|History of Present Illness|3975,3978|false|false|false|C0489633|Review of systems (procedure)|ROS
Event|Event|History of Present Illness|3983,3992|false|false|false|||conducted
Event|Event|History of Present Illness|4001,4009|false|false|false|||negative
Finding|Classification|History of Present Illness|4001,4009|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|History of Present Illness|4001,4009|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|History of Present Illness|4001,4009|false|false|false|C5237010|Expression Negative|negative
Finding|Idea or Concept|History of Present Illness|4020,4025|false|false|false|C1552828|Table Frame - above|above
Disorder|Disease or Syndrome|History of Present Illness|4034,4037|false|false|false|C0268529|Proline dehydrogenase deficiency|HPI
Event|Event|History of Present Illness|4034,4037|false|false|false|||HPI
Finding|Finding|History of Present Illness|4034,4037|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Finding|Molecular Function|History of Present Illness|4034,4037|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Disorder|Disease or Syndrome|Past Medical History|4063,4075|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|Past Medical History|4063,4075|false|false|false|||Hypertension
Procedure|Diagnostic Procedure|Past Medical History|4077,4089|false|false|false|C0031150|Laparoscopy|laparoscopic
Procedure|Therapeutic or Preventive Procedure|Past Medical History|4077,4105|false|false|false|C0162522|Cholecystectomy, Laparoscopic|laparoscopic cholecystectomy
Event|Event|Past Medical History|4090,4105|false|false|false|||cholecystectomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|4090,4105|false|false|false|C0008320|Cholecystectomy procedure|cholecystectomy
Finding|Functional Concept|Past Medical History|4107,4111|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|Past Medical History|4107,4116|false|false|false|C0230432;C4281599|Structure of left knee;Structure of left knee region|left knee
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|4107,4116|false|false|false|C0230432;C4281599|Structure of left knee;Structure of left knee region|left knee
Anatomy|Body Location or Region|Past Medical History|4112,4116|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|4112,4116|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Space or Junction|Past Medical History|4112,4116|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Procedure|Diagnostic Procedure|Past Medical History|4112,4116|false|false|false|C0562271|Examination of knee joint|knee
Event|Event|Past Medical History|4118,4129|false|false|false|||replacement
Finding|Functional Concept|Past Medical History|4118,4129|false|false|false|C0559956|Replacement|replacement
Procedure|Health Care Activity|Past Medical History|4118,4129|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Procedure|Therapeutic or Preventive Procedure|Past Medical History|4118,4129|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Finding|Gene or Genome|Past Medical History|4147,4150|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|Past Medical History|4152,4163|false|false|false|||laminectomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|4152,4163|false|false|false|C0022983|Laminectomy|laminectomy
Attribute|Clinical Attribute|Past Medical History|4176,4179|false|false|false|C1114365||age
Drug|Biologically Active Substance|Past Medical History|4176,4179|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|Past Medical History|4176,4179|false|false|false|C0162574|Glycation End Products, Advanced|age
Event|Event|Past Medical History|4176,4179|false|false|false|||age
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|4190,4197|false|false|false|C0042232|Vagina|vaginal
Drug|Biomedical or Dental Material|Past Medical History|4190,4197|false|false|false|C1272941|Vaginal Dosage Form|vaginal
Finding|Finding|Past Medical History|4190,4197|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Finding|Functional Concept|Past Medical History|4190,4197|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Event|Event|Past Medical History|4198,4208|false|false|false|||deliveries
Event|Event|Past Medical History|4240,4252|false|false|false|||laparoscopic
Procedure|Diagnostic Procedure|Past Medical History|4240,4252|false|false|false|C0031150|Laparoscopy|laparoscopic
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|4263,4269|false|false|false|C0030797|Pelvis|pelvic
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|4263,4280|false|false|false|C0729595|Pelvic lymph node group|pelvic lymph node
Finding|Body Substance|Past Medical History|4270,4275|false|false|false|C0024202|Lymph|lymph
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|4270,4280|false|false|false|C0024204|lymph nodes|lymph node
Event|Event|Past Medical History|4282,4292|false|false|false|||dissection
Finding|Pathologic Function|Past Medical History|4282,4292|false|false|false|C0333288|Dissecting hemorrhage|dissection
Procedure|Therapeutic or Preventive Procedure|Past Medical History|4282,4292|false|false|false|C0012737|Tissue Dissection|dissection
Event|Event|Past Medical History|4312,4324|false|false|false|||hysterectomy
Finding|Finding|Past Medical History|4312,4324|false|false|false|C1548863|Consent Type - Hysterectomy|hysterectomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|4312,4324|false|false|false|C0020699|Hysterectomy|hysterectomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|4329,4351|false|false|false|C0278321|Bilateral oophorectomy|bilateral oophorectomy
Event|Event|Past Medical History|4339,4351|false|false|false|||oophorectomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|4339,4351|false|false|false|C0029936|Ovariectomy|oophorectomy
Finding|Gene or Genome|Past Medical History|4357,4362|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Finding|Finding|Past Medical History|4357,4369|false|false|false|C0151994|Enlarged uterus|large uterus
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|4363,4369|false|false|false|C0042149;C1519876;C4266525|Mouse Uterus;Pelvis>Uterus;Uterus|uterus
Anatomy|Tissue|Past Medical History|4363,4369|false|false|false|C0042149;C1519876;C4266525|Mouse Uterus;Pelvis>Uterus;Uterus|uterus
Disorder|Disease or Syndrome|Past Medical History|4363,4369|false|false|false|C0042131;C0496919|Neoplasm of uncertain or unknown behavior of uterus;Uterine Diseases|uterus
Disorder|Neoplastic Process|Past Medical History|4363,4369|false|false|false|C0042131;C0496919|Neoplasm of uncertain or unknown behavior of uterus;Uterine Diseases|uterus
Event|Event|Past Medical History|4363,4369|false|false|false|||uterus
Procedure|Diagnostic Procedure|Past Medical History|4363,4369|false|false|false|C0869889|examination of uterus|uterus
Finding|Gene or Genome|Past Medical History|4400,4405|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Disorder|Neoplastic Process|Past Medical History|4406,4413|false|false|false|C0023267|Fibroid Tumor|fibroid
Event|Event|Past Medical History|4406,4413|false|false|false|||fibroid
Procedure|Diagnostic Procedure|Past Medical History|4418,4430|false|false|false|C0031150|Laparoscopy|Laparoscopic
Procedure|Therapeutic or Preventive Procedure|Past Medical History|4418,4449|false|false|false|C5879917|Laparoscopic radical cystectomy|Laparoscopic radical cystectomy
Drug|Chemical Viewed Structurally|Past Medical History|4431,4438|false|false|false|C0302912|Radicals (chemistry)|radical
Procedure|Therapeutic or Preventive Procedure|Past Medical History|4431,4449|false|false|false|C0194401|Complete cystectomy|radical cystectomy
Event|Event|Past Medical History|4439,4449|false|false|false|||cystectomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|4439,4449|false|false|false|C0010651|Cystectomy|cystectomy
Disorder|Disease or Syndrome|Past Medical History|4454,4462|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Event|Event|Past Medical History|4463,4474|false|false|false|||vaginectomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|4463,4474|false|false|false|C0195130|Vaginectomy|vaginectomy
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|4481,4488|false|false|false|C0042232|Vagina|vaginal
Drug|Biomedical or Dental Material|Past Medical History|4481,4488|false|false|false|C1272941|Vaginal Dosage Form|vaginal
Finding|Finding|Past Medical History|4481,4488|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Finding|Functional Concept|Past Medical History|4481,4488|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Procedure|Therapeutic or Preventive Procedure|Past Medical History|4481,4503|false|false|false|C0195196|Reconstruction of vagina|vaginal reconstruction
Event|Event|Past Medical History|4489,4503|false|false|false|||reconstruction
Procedure|Machine Activity|Past Medical History|4489,4503|false|false|false|C0020912;C0524865|Optical Image Reconstruction;Reconstructive Surgical Procedures|reconstruction
Procedure|Therapeutic or Preventive Procedure|Past Medical History|4489,4503|false|false|false|C0020912;C0524865|Optical Image Reconstruction;Reconstructive Surgical Procedures|reconstruction
Event|Event|Family Medical History|4544,4552|false|false|false|||Negative
Finding|Classification|Family Medical History|4544,4552|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Finding|Finding|Family Medical History|4544,4552|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Lab|Laboratory or Test Result|Family Medical History|4544,4552|false|false|false|C5237010|Expression Negative|Negative
Finding|Finding|Family Medical History|4544,4556|false|false|false|C0205160|Negative|Negative for
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|4557,4564|true|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|Family Medical History|4557,4564|true|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Event|Event|Family Medical History|4557,4564|true|false|false|||bladder
Procedure|Therapeutic or Preventive Procedure|Family Medical History|4557,4564|true|false|false|C0872388|Procedures on bladder|bladder
Disorder|Neoplastic Process|Family Medical History|4557,4567|true|true|false|C0005684|Malignant neoplasm of urinary bladder|bladder CA
Procedure|Health Care Activity|General Exam|4587,4596|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|General Exam|4597,4601|false|false|false|||EXAM
Finding|Functional Concept|General Exam|4597,4601|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|4597,4601|false|false|false|C0582103|Medical Examination|EXAM
Finding|Classification|General Exam|4604,4607|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Finding|Gene or Genome|General Exam|4604,4607|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Disorder|Disease or Syndrome|General Exam|4609,4612|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|4609,4612|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|4609,4612|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|4609,4612|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|4609,4612|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|General Exam|4609,4612|false|false|false|||NAD
Finding|Finding|General Exam|4609,4612|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Event|Event|General Exam|4614,4622|false|false|false|||speaking
Finding|Idea or Concept|General Exam|4628,4632|false|false|false|C1705313|Term (lexical)|word
Event|Event|General Exam|4633,4642|true|false|false|||sentences
Finding|Intellectual Product|General Exam|4633,4642|true|false|false|C0876929|Sentence|sentences
Event|Event|General Exam|4644,4650|true|false|false|||pursed
Anatomy|Body Part, Organ, or Organ Component|General Exam|4651,4654|true|false|false|C0023759|Lip structure|lip
Disorder|Disease or Syndrome|General Exam|4651,4654|true|false|false|C0153932;C0264511|Benign neoplasm of the lip;Lymphoid interstitial pneumonia|lip
Disorder|Neoplastic Process|General Exam|4651,4654|true|false|false|C0153932;C0264511|Benign neoplasm of the lip;Lymphoid interstitial pneumonia|lip
Finding|Gene or Genome|General Exam|4651,4654|true|false|false|C1846919;C3889123|SMG1 gene;SMG1 wt Allele|lip
Attribute|Clinical Attribute|General Exam|4655,4664|true|false|false|C5885990||breathing
Event|Event|General Exam|4655,4664|true|false|false|||breathing
Finding|Finding|General Exam|4655,4664|true|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|General Exam|4655,4664|true|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|General Exam|4655,4664|true|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|General Exam|4655,4664|true|false|false|C1160636|respiratory system process|breathing
Disorder|Congenital Abnormality|General Exam|4670,4686|true|false|false|C0158784|Accessory skeletal muscle|accessory muscle
Finding|Finding|General Exam|4670,4690|true|false|false|C1821466|Use of accessory muscles|accessory muscle use
Anatomy|Body Part, Organ, or Organ Component|General Exam|4680,4686|true|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|General Exam|4680,4686|true|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Event|Event|General Exam|4687,4690|true|false|false|||use
Finding|Functional Concept|General Exam|4687,4690|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|General Exam|4687,4690|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Event|Event|General Exam|4692,4697|true|false|false|||lying
Disorder|Disease or Syndrome|General Exam|4701,4704|true|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Event|Event|General Exam|4701,4704|true|false|false|||bed
Finding|Intellectual Product|General Exam|4701,4704|true|false|false|C2346952|Bachelor of Education|bed
Anatomy|Body Part, Organ, or Organ Component|General Exam|4706,4710|false|false|false|C0015392|Eye|Eyes
Attribute|Clinical Attribute|General Exam|4706,4710|false|false|false|C5848506||Eyes
Event|Event|General Exam|4712,4716|false|false|false|||EOMI
Event|Event|General Exam|4726,4735|false|false|false|||anicteric
Finding|Finding|General Exam|4726,4735|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Location or Region|General Exam|4739,4742|false|false|false|C0150934;C0175196|Ear, nose and throat;Structure of entorhinal cortex|ENT
Anatomy|Body Part, Organ, or Organ Component|General Exam|4739,4742|false|false|false|C0150934;C0175196|Ear, nose and throat;Structure of entorhinal cortex|ENT
Finding|Gene or Genome|General Exam|4739,4742|false|false|false|C0262471;C1417861;C3889152|ENT problem;NT5E gene;NT5E wt Allele|ENT
Finding|Sign or Symptom|General Exam|4739,4742|false|false|false|C0262471;C1417861;C3889152|ENT problem;NT5E gene;NT5E wt Allele|ENT
Anatomy|Body Part, Organ, or Organ Component|General Exam|4744,4747|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|General Exam|4744,4747|false|false|false|C0026987|Myelofibrosis|MMM
Event|Event|General Exam|4744,4747|false|false|false|||MMM
Event|Event|General Exam|4752,4757|false|false|false|||clear
Finding|Idea or Concept|General Exam|4752,4757|false|false|false|C1550016|Remote control command - Clear|clear
Event|Event|General Exam|4771,4774|true|false|false|||RRR
Event|Event|General Exam|4779,4782|true|false|false|||MRG
Finding|Gene or Genome|General Exam|4779,4782|true|false|false|C1422304|MAS1L gene|MRG
Drug|Food|General Exam|4789,4795|true|false|false|C5890763||pulses
Event|Event|General Exam|4789,4795|true|false|false|||pulses
Finding|Physiologic Function|General Exam|4789,4795|true|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|4789,4795|true|false|false|C0034107|Pulse taking|pulses
Attribute|Clinical Attribute|General Exam|4800,4805|false|false|false|C1717255||edema
Event|Event|General Exam|4800,4805|false|false|false|||edema
Finding|Pathologic Function|General Exam|4800,4805|false|false|false|C0013604|Edema|edema
Event|Event|General Exam|4824,4835|true|false|false|||compression
Finding|Functional Concept|General Exam|4824,4835|true|false|false|C0332459;C4551657|Compressed structure|compression
Phenomenon|Natural Phenomenon or Process|General Exam|4824,4835|true|false|false|C0728907|Compression|compression
Procedure|Machine Activity|General Exam|4824,4835|true|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Procedure|Therapeutic or Preventive Procedure|General Exam|4824,4835|true|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Event|Event|General Exam|4836,4845|true|false|false|||stockings
Event|Activity|General Exam|4849,4854|true|false|false|C1882509|put - instruction imperative|place
Event|Event|General Exam|4849,4854|true|false|false|||place
Finding|Functional Concept|General Exam|4849,4854|true|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|General Exam|4849,4854|true|false|false|C1533810||place
Event|Event|General Exam|4859,4862|true|false|false|||JVD
Finding|Finding|General Exam|4859,4862|true|false|false|C0425687|Jugular venous engorgement|JVD
Attribute|Clinical Attribute|General Exam|4865,4869|true|false|false|C0231832|Respiratory rate|Resp
Disorder|Disease or Syndrome|General Exam|4865,4869|true|false|false|C0851355|Respiratory, thoracic and mediastinal disorders|Resp
Event|Event|General Exam|4865,4869|true|false|false|||Resp
Event|Event|General Exam|4878,4884|true|false|false|||effort
Finding|Organism Function|General Exam|4878,4884|true|false|false|C0015264|Exertion|effort
Disorder|Congenital Abnormality|General Exam|4889,4905|true|false|false|C0158784|Accessory skeletal muscle|accessory muscle
Finding|Finding|General Exam|4889,4909|true|false|false|C1821466|Use of accessory muscles|accessory muscle use
Anatomy|Body Part, Organ, or Organ Component|General Exam|4899,4905|true|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|General Exam|4899,4905|true|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Event|Event|General Exam|4906,4909|true|false|false|||use
Finding|Functional Concept|General Exam|4906,4909|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|General Exam|4906,4909|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Anatomy|Body Part, Organ, or Organ Component|General Exam|4911,4916|true|false|false|C0024109|Lung|lungs
Drug|Amino Acid, Peptide, or Protein|General Exam|4917,4920|true|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|General Exam|4917,4920|true|false|false|||CTA
Finding|Gene or Genome|General Exam|4917,4920|true|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|General Exam|4917,4920|true|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Disorder|Disease or Syndrome|General Exam|4929,4937|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Event|Event|General Exam|4938,4950|false|false|false|||auscultation
Procedure|Diagnostic Procedure|General Exam|4938,4950|false|false|false|C0004339|Auscultation|auscultation
Disorder|Disease or Syndrome|General Exam|4957,4961|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|General Exam|4957,4961|false|false|false|||soft
Anatomy|Anatomical Structure|General Exam|4976,4984|true|false|false|C0559495|Urological stoma|Urostomy
Procedure|Therapeutic or Preventive Procedure|General Exam|4976,4984|true|false|false|C0856443|Urostomy procedure|Urostomy
Finding|Finding|General Exam|4976,4989|true|false|false|C4053891|Urostomy Site|Urostomy site
Anatomy|Body Location or Region|General Exam|4985,4989|true|false|false|C1515974|Anatomic Site|site
Finding|Intellectual Product|General Exam|4985,4989|true|false|false|C1546778||site
Event|Event|General Exam|4999,5005|true|false|false|||appear
Event|Event|General Exam|5006,5014|true|false|false|||infected
Finding|Finding|General Exam|5006,5014|true|true|false|C0439663|Infected|infected
Disorder|Congenital Abnormality|General Exam|5016,5019|true|false|false|C0022681|Medullary sponge kidney|MSK
Disorder|Disease or Syndrome|General Exam|5016,5019|true|false|false|C0022681|Medullary sponge kidney|MSK
Event|Event|General Exam|5016,5019|true|false|false|||MSK
Finding|Gene or Genome|General Exam|5016,5019|true|false|false|C1420279|SIK1 gene|MSK
Finding|Idea or Concept|General Exam|5024,5035|true|false|false|C0750502|Significant|significant
Disorder|Acquired Abnormality|General Exam|5036,5044|true|false|false|C0022821;C0022822;C0265673|Acquired kyphosis;Congenital kyphosis;Kyphosis deformity of spine|kyphosis
Disorder|Anatomical Abnormality|General Exam|5036,5044|true|false|false|C0022821;C0022822;C0265673|Acquired kyphosis;Congenital kyphosis;Kyphosis deformity of spine|kyphosis
Disorder|Congenital Abnormality|General Exam|5036,5044|true|false|false|C0022821;C0022822;C0265673|Acquired kyphosis;Congenital kyphosis;Kyphosis deformity of spine|kyphosis
Event|Event|General Exam|5036,5044|true|false|false|||kyphosis
Finding|Finding|General Exam|5036,5044|true|false|false|C2115817|kyphosis|kyphosis
Disorder|Disease or Syndrome|General Exam|5058,5067|true|false|false|C0039103|Synovitis|synovitis
Event|Event|General Exam|5058,5067|true|false|false|||synovitis
Anatomy|Body System|General Exam|5070,5074|false|false|false|C1123023;C4520765|Skin;Skin, Human|Skin
Disorder|Disease or Syndrome|General Exam|5070,5074|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Disorder|Neoplastic Process|General Exam|5070,5074|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Finding|Body Substance|General Exam|5070,5074|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Finding|Intellectual Product|General Exam|5070,5074|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Disorder|Disease or Syndrome|General Exam|5087,5091|true|false|false|C5779629|Eruption of skin (disorder)|rash
Event|Event|General Exam|5087,5091|true|false|false|||rash
Finding|Pathologic Function|General Exam|5087,5091|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|General Exam|5087,5091|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Event|Event|General Exam|5096,5104|true|false|false|||jaundice
Finding|Finding|General Exam|5096,5104|true|false|false|C0022346;C2010848;C2203646|Icterus;jaundice;yellow skin or eyes (symptom)|jaundice
Finding|Sign or Symptom|General Exam|5096,5104|true|false|false|C0022346;C2010848;C2203646|Icterus;jaundice;yellow skin or eyes (symptom)|jaundice
Event|Event|General Exam|5114,5119|false|false|false|||AAOx3
Anatomy|Body Location or Region|General Exam|5124,5130|true|false|false|C0015450|Face|facial
Disorder|Disease or Syndrome|General Exam|5124,5136|true|false|false|C0427055|Facial Paresis|facial droop
Finding|Finding|General Exam|5124,5136|true|false|false|C4022719|Unilateral facial palsy|facial droop
Event|Event|General Exam|5131,5136|true|false|false|||droop
Disorder|Mental or Behavioral Dysfunction|General Exam|5139,5144|false|false|false|C0004936;C1306597|Mental disorders;Psychiatric problem|Psych
Event|Event|General Exam|5139,5144|false|false|false|||Psych
Event|Event|General Exam|5151,5156|false|false|false|||range
Finding|Intellectual Product|General Exam|5151,5156|false|false|false|C3542016|Concept model range (foundation metadata concept)|range
Event|Event|General Exam|5160,5166|false|false|false|||affect
Finding|Mental Process|General Exam|5160,5166|false|false|false|C0001721|Affect (mental function)|affect
Procedure|Health Care Activity|General Exam|5160,5166|false|false|false|C2237113|assessment of affect|affect
Finding|Body Substance|General Exam|5169,5178|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|5169,5178|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|5169,5178|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|5169,5178|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|General Exam|5179,5183|false|false|false|||EXAM
Finding|Functional Concept|General Exam|5179,5183|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|5179,5183|false|false|false|C0582103|Medical Examination|EXAM
Event|Event|General Exam|5185,5191|false|false|false|||vitals
Finding|Classification|General Exam|5218,5221|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Finding|Gene or Genome|General Exam|5218,5221|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Event|Event|General Exam|5223,5228|true|false|false|||Lying
Finding|Individual Behavior|General Exam|5223,5228|true|false|false|C0600261|Telling untruths|Lying
Disorder|Disease or Syndrome|General Exam|5232,5235|true|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Finding|Intellectual Product|General Exam|5232,5235|true|false|false|C2346952|Bachelor of Education|bed
Finding|Idea or Concept|General Exam|5242,5250|true|false|false|C0750489|apparent|apparent
Event|Event|General Exam|5251,5259|true|false|false|||distress
Finding|Finding|General Exam|5251,5259|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|General Exam|5251,5259|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|General Exam|5260,5265|true|false|false|C1512338|HEENT|HEENT
Event|Event|General Exam|5267,5276|false|false|false|||Anicteric
Finding|Finding|General Exam|5267,5276|false|false|false|C0205180|Anicteric|Anicteric
Anatomy|Body Part, Organ, or Organ Component|General Exam|5278,5281|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|General Exam|5278,5281|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body System|General Exam|5282,5296|false|false|false|C0007226;C3887460|Cardiovascular;Cardiovascular system|Cardiovascular
Event|Event|General Exam|5298,5301|true|false|false|||RRR
Finding|Functional Concept|General Exam|5320,5325|true|false|false|C1552823|Table Cell Horizontal Align - right|right
Disorder|Disease or Syndrome|General Exam|5332,5337|true|false|false|C3714496|Chronic obstructive pulmonary disease of horses|heave
Event|Event|General Exam|5332,5337|true|false|false|||heave
Finding|Organ or Tissue Function|General Exam|5344,5352|false|false|false|C0039155|Systole|systolic
Finding|Finding|General Exam|5344,5359|false|false|false|C0232257|Systolic Murmurs|systolic murmur
Event|Event|General Exam|5353,5359|false|false|false|||murmur
Finding|Finding|General Exam|5353,5359|false|false|false|C0018808|Heart murmur|murmur
Anatomy|Body Part, Organ, or Organ Component|General Exam|5361,5370|false|false|false|C0024109|Lung|Pulmonary
Attribute|Clinical Attribute|General Exam|5361,5370|false|false|false|C2707265||Pulmonary
Finding|Finding|General Exam|5361,5370|false|false|false|C4522268|Pulmonary (intended site)|Pulmonary
Anatomy|Body Location or Region|General Exam|5372,5376|false|false|false|C0024109;C4037972|Chest>Lung;Lung|Lung
Anatomy|Body Part, Organ, or Organ Component|General Exam|5372,5376|false|false|false|C0024109;C4037972|Chest>Lung;Lung|Lung
Disorder|Disease or Syndrome|General Exam|5372,5376|false|false|false|C0024115|Lung diseases|Lung
Finding|Finding|General Exam|5372,5376|false|false|false|C0740941|Lung Problem|Lung
Event|Event|General Exam|5377,5383|false|false|false|||fields
Event|Event|General Exam|5384,5389|false|false|false|||clear
Finding|Idea or Concept|General Exam|5384,5389|false|false|false|C1550016|Remote control command - Clear|clear
Event|Event|General Exam|5393,5405|false|false|false|||auscultation
Procedure|Diagnostic Procedure|General Exam|5393,5405|false|false|false|C0004339|Auscultation|auscultation
Event|Event|General Exam|5422,5430|true|false|false|||crackles
Finding|Finding|General Exam|5422,5430|true|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Event|Event|General Exam|5434,5442|true|false|false|||wheezing
Finding|Sign or Symptom|General Exam|5434,5442|true|false|false|C0043144|Wheezing|wheezing
Disorder|Disease or Syndrome|General Exam|5449,5453|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|General Exam|5449,5453|false|false|false|||Soft
Event|Event|General Exam|5455,5464|false|false|false|||distended
Finding|Finding|General Exam|5455,5464|false|false|false|C0700124|Dilated|distended
Event|Event|General Exam|5466,5475|false|false|false|||nontender
Anatomy|Body Part, Organ, or Organ Component|General Exam|5477,5482|false|false|false|C0021853|Intestines|bowel
Finding|Finding|General Exam|5477,5489|false|false|false|C0232693|Bowel sounds|bowel sounds
Event|Event|General Exam|5483,5489|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|General Exam|5483,5489|false|false|false|C0037709||sounds
Finding|Finding|General Exam|5490,5497|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|General Exam|5490,5497|false|false|false|C0150312;C0449450|Present;Presentation|present
Anatomy|Anatomical Structure|General Exam|5499,5507|false|false|false|C0559495|Urological stoma|urostomy
Procedure|Therapeutic or Preventive Procedure|General Exam|5499,5507|false|false|false|C0856443|Urostomy procedure|urostomy
Event|Activity|General Exam|5512,5517|false|false|false|C1882509|put - instruction imperative|place
Event|Event|General Exam|5512,5517|false|false|false|||place
Finding|Functional Concept|General Exam|5512,5517|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|General Exam|5512,5517|false|false|false|C1533810||place
Anatomy|Body Part, Organ, or Organ Component|General Exam|5519,5530|false|false|false|C0015385;C0278454|All extremities;Limb structure|Extremities
Attribute|Clinical Attribute|General Exam|5535,5540|true|false|false|C1717255||edema
Event|Event|General Exam|5535,5540|true|false|false|||edema
Finding|Pathologic Function|General Exam|5535,5540|true|false|false|C0013604|Edema|edema
Finding|Functional Concept|General Exam|5549,5553|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|General Exam|5549,5557|false|false|false|C0230416;C0230443|Left lower extremity;Structure of left lower leg|left leg
Anatomy|Body Part, Organ, or Organ Component|General Exam|5554,5557|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Event|Event|General Exam|5566,5572|false|false|false|||larger
Event|Event|General Exam|5578,5583|false|false|false|||right
Finding|Functional Concept|General Exam|5578,5583|false|true|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|General Exam|5585,5588|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Event|Event|General Exam|5590,5594|false|false|false|||warm
Finding|Finding|General Exam|5590,5594|false|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|General Exam|5590,5594|false|false|false|C0687712|warming process|warm
Finding|Finding|General Exam|5596,5600|false|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|5601,5609|false|false|false|||perfused
Finding|Functional Concept|General Exam|5615,5620|false|false|false|C1513492|motor movement|motor
Finding|Finding|General Exam|5615,5629|false|false|false|C5551447|Motor function (finding)|motor function
Phenomenon|Biologic Function|General Exam|5615,5629|false|false|false|C0234130|Motor function (observable entity)|motor function
Event|Event|General Exam|5621,5629|false|false|false|||function
Finding|Finding|General Exam|5621,5629|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|General Exam|5621,5629|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|General Exam|5621,5629|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|General Exam|5621,5629|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Event|Event|General Exam|5630,5636|false|false|false|||intact
Finding|Finding|General Exam|5630,5636|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Functional Concept|General Exam|5642,5646|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|General Exam|5648,5653|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|5648,5653|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|General Exam|5648,5657|false|false|false|C1140621;C4299093|Leg;Lower extremity>Lower leg|lower leg
Anatomy|Body Part, Organ, or Organ Component|General Exam|5654,5657|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Event|Event|General Exam|5661,5668|false|false|false|||wrapped
Event|Event|General Exam|5693,5697|false|false|false|||LABS
Lab|Laboratory or Test Result|General Exam|5693,5697|false|false|false|C0587081|Laboratory test finding|LABS
Procedure|Health Care Activity|General Exam|5726,5735|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Lab|Laboratory or Test Result|General Exam|5736,5740|false|false|false|C0587081|Laboratory test finding|labs
Drug|Biologically Active Substance|General Exam|5756,5763|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|General Exam|5756,5763|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|General Exam|5756,5763|false|false|false|C0017725|glucose|GLUCOSE
Event|Event|General Exam|5756,5763|false|false|false|||GLUCOSE
Lab|Laboratory or Test Result|General Exam|5756,5763|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|General Exam|5756,5763|false|false|false|C0337438|Glucose measurement|GLUCOSE
Drug|Biologically Active Substance|General Exam|5769,5773|false|false|false|C0041942|urea|UREA
Drug|Organic Chemical|General Exam|5769,5773|false|false|false|C0041942|urea|UREA
Drug|Pharmacologic Substance|General Exam|5769,5773|false|false|false|C0041942|urea|UREA
Event|Event|General Exam|5769,5773|false|false|false|||UREA
Procedure|Laboratory Procedure|General Exam|5769,5773|false|false|false|C0523961|Urea measurement|UREA
Drug|Biologically Active Substance|General Exam|5790,5796|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Element, Ion, or Isotope|General Exam|5790,5796|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Pharmacologic Substance|General Exam|5790,5796|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Event|Event|General Exam|5790,5796|false|false|false|||SODIUM
Finding|Physiologic Function|General Exam|5790,5796|false|false|false|C4553025|Sodium metabolic function|SODIUM
Procedure|Laboratory Procedure|General Exam|5790,5796|false|false|false|C0337443|Sodium measurement|SODIUM
Drug|Biologically Active Substance|General Exam|5802,5811|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Element, Ion, or Isotope|General Exam|5802,5811|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Food|General Exam|5802,5811|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Inorganic Chemical|General Exam|5802,5811|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Pharmacologic Substance|General Exam|5802,5811|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Event|Event|General Exam|5802,5811|false|false|false|||POTASSIUM
Finding|Physiologic Function|General Exam|5802,5811|false|false|false|C4553027|Potassium metabolic function|POTASSIUM
Procedure|Laboratory Procedure|General Exam|5802,5811|false|false|false|C0202194|Potassium measurement|POTASSIUM
Drug|Element, Ion, or Isotope|General Exam|5816,5824|false|false|false|C0008203;C0596019|Chlorides;chloride ion|CHLORIDE
Event|Event|General Exam|5816,5824|false|false|false|||CHLORIDE
Finding|Physiologic Function|General Exam|5816,5824|false|false|false|C4553021|Chloride metabolic function|CHLORIDE
Procedure|Laboratory Procedure|General Exam|5816,5824|false|false|false|C0201952|Chloride measurement|CHLORIDE
Drug|Biologically Active Substance|General Exam|5834,5837|false|false|false|C0007012|carbon dioxide|CO2
Drug|Inorganic Chemical|General Exam|5834,5837|false|false|false|C0007012|carbon dioxide|CO2
Event|Event|General Exam|5834,5837|false|false|false|||CO2
Finding|Finding|General Exam|5834,5837|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Finding|Gene or Genome|General Exam|5834,5837|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Drug|Element, Ion, or Isotope|General Exam|5841,5846|false|false|false|C0003075|Anions|ANION
Attribute|Clinical Attribute|General Exam|5841,5850|false|false|false|C0003074|Anion Gap|ANION GAP
Lab|Laboratory or Test Result|General Exam|5841,5850|false|false|false|C1509129|Anion gap result|ANION GAP
Procedure|Laboratory Procedure|General Exam|5841,5850|false|false|false|C0201889;C2189246|Anion gap measurement;blood anion gap (lab test)|ANION GAP
Drug|Amino Acid, Peptide, or Protein|General Exam|5847,5850|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Drug|Biologically Active Substance|General Exam|5847,5850|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Event|Event|General Exam|5847,5850|false|false|false|||GAP
Finding|Gene or Genome|General Exam|5847,5850|false|false|false|C1419277;C2984552|RASA1 gene;RASA1 wt Allele|GAP
Drug|Amino Acid, Peptide, or Protein|General Exam|5896,5902|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Drug|Hormone|General Exam|5896,5902|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Event|Event|General Exam|5896,5902|false|false|false|||proBNP
Anatomy|Cell|General Exam|5921,5924|false|false|false|C0023516|Leukocytes|WBC
Event|Event|General Exam|5921,5924|false|false|false|||WBC
Anatomy|Cell|General Exam|5929,5932|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|5929,5932|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|5929,5932|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|5939,5942|false|false|false|C0019046|Hemoglobin|HGB
Drug|Biologically Active Substance|General Exam|5939,5942|false|false|false|C0019046|Hemoglobin|HGB
Event|Event|General Exam|5939,5942|false|false|false|||HGB
Finding|Gene or Genome|General Exam|5939,5942|false|false|false|C1424337|CYGB gene|HGB
Lab|Laboratory or Test Result|General Exam|5939,5942|false|false|false|C0019029|Hemoglobin concentration|HGB
Procedure|Laboratory Procedure|General Exam|5948,5951|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|General Exam|5948,5951|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Disorder|Virus|General Exam|5958,5961|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|5958,5961|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|5958,5961|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|5958,5961|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|5958,5961|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|5966,5969|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|5966,5969|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|5966,5969|false|false|false|||MCH
Finding|Gene or Genome|General Exam|5966,5969|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|5966,5969|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|5966,5969|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|5975,5979|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|5975,5979|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Event|Event|General Exam|6021,6024|false|false|false|||PLT
Procedure|Laboratory Procedure|General Exam|6021,6024|false|false|false|C0201617|Primed lymphocyte test|PLT
Disorder|Neoplastic Process|General Exam|6054,6057|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|General Exam|6054,6057|false|false|false|||PTT
Procedure|Laboratory Procedure|General Exam|6054,6057|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Finding|Body Substance|General Exam|6068,6077|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|General Exam|6068,6077|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|General Exam|6068,6077|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|General Exam|6068,6077|false|false|false|C0030685|Patient Discharge|Discharge
Lab|Laboratory or Test Result|General Exam|6078,6082|false|false|false|C0587081|Laboratory test finding|labs
Disorder|Disease or Syndrome|General Exam|6096,6101|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|6096,6101|false|false|false|||BLOOD
Finding|Body Substance|General Exam|6096,6101|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|6102,6105|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|6112,6115|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|6112,6115|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|6112,6115|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|6122,6125|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|6122,6125|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|6122,6125|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|6122,6125|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|6131,6134|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|6131,6134|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|6142,6145|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|6142,6145|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|6142,6145|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|6142,6145|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|6142,6145|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|6149,6152|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|6149,6152|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|6149,6152|false|false|false|||MCH
Finding|Gene or Genome|General Exam|6149,6152|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|6149,6152|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|6149,6152|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|6158,6162|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|6158,6162|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|6190,6193|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|6210,6215|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|6210,6215|false|false|false|||BLOOD
Finding|Body Substance|General Exam|6210,6215|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|6210,6223|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|6210,6223|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|6210,6223|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|6216,6223|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|6216,6223|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|6216,6223|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|6216,6223|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|6216,6223|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|6216,6223|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|6267,6271|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|6267,6271|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|6267,6271|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|6296,6301|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|6296,6301|false|false|false|||BLOOD
Finding|Body Substance|General Exam|6296,6301|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|6296,6309|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|General Exam|6302,6309|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|6302,6309|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|6302,6309|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|6302,6309|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|6302,6309|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|General Exam|6302,6309|false|false|false|||Calcium
Finding|Physiologic Function|General Exam|6302,6309|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|6302,6309|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|General Exam|6343,6348|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|6343,6348|false|false|false|||BLOOD
Finding|Body Substance|General Exam|6343,6348|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|6375,6378|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Biologically Active Substance|General Exam|6375,6378|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Hormone|General Exam|6375,6378|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Pharmacologic Substance|General Exam|6375,6378|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Finding|Gene or Genome|General Exam|6375,6378|false|false|false|C1334121;C1336604;C1705002|IL5 gene;TERF1 gene;TERF1 wt Allele|TRF
Disorder|Disease or Syndrome|General Exam|6396,6401|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|6396,6401|false|false|false|||BLOOD
Finding|Body Substance|General Exam|6396,6401|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|6396,6406|false|false|false|C0853169|Blood iron measurement|BLOOD Iron
Drug|Biologically Active Substance|General Exam|6402,6406|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Element, Ion, or Isotope|General Exam|6402,6406|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Pharmacologic Substance|General Exam|6402,6406|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Event|Event|General Exam|6402,6406|false|false|false|||Iron
Procedure|Laboratory Procedure|General Exam|6402,6406|false|false|false|C0337439|Iron measurement|Iron
Event|Event|General Exam|6412,6424|false|false|false|||MICROBIOLOGY
Finding|Functional Concept|General Exam|6412,6424|false|false|false|C0025953;C1571921;C4049106|Microbiological;Microbiology - Laboratory Class;Microbiology Diagnostic Service Section ID|MICROBIOLOGY
Finding|Intellectual Product|General Exam|6412,6424|false|false|false|C0025953;C1571921;C4049106|Microbiological;Microbiology - Laboratory Class;Microbiology Diagnostic Service Section ID|MICROBIOLOGY
Procedure|Laboratory Procedure|General Exam|6412,6424|false|false|false|C0085672|Microbiology procedure|MICROBIOLOGY
Finding|Body Substance|General Exam|6464,6469|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|6464,6469|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|6464,6469|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Idea or Concept|General Exam|6501,6506|false|false|false|C1546485|Diagnosis Type - Final|FINAL
Finding|Intellectual Product|General Exam|6501,6513|false|false|false|C0460114|Final report|FINAL REPORT
Attribute|Clinical Attribute|General Exam|6507,6513|false|false|false|C4255046||REPORT
Event|Event|General Exam|6507,6513|false|false|false|||REPORT
Finding|Intellectual Product|General Exam|6507,6513|false|false|false|C0684224|Report (document)|REPORT
Procedure|Health Care Activity|General Exam|6507,6513|false|false|false|C0700287|Reporting|REPORT
Finding|Body Substance|General Exam|6522,6527|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|6522,6527|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|6522,6527|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Procedure|Laboratory Procedure|General Exam|6522,6535|false|false|false|C0430404|Urine culture|URINE CULTURE
Drug|Biomedical or Dental Material|General Exam|6528,6535|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|General Exam|6528,6535|false|false|false|||CULTURE
Finding|Functional Concept|General Exam|6528,6535|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|General Exam|6528,6535|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|General Exam|6528,6535|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|General Exam|6537,6542|false|false|false|||Final
Finding|Idea or Concept|General Exam|6537,6542|false|false|false|C1546485|Diagnosis Type - Final|Final
Event|Event|General Exam|6555,6560|false|false|false|||MIXED
Anatomy|Cell|General Exam|6584,6590|false|false|false|C1947989|Colony (cells or organisms)|COLONY
Event|Event|General Exam|6599,6609|false|false|false|||CONSISTENT
Finding|Idea or Concept|General Exam|6599,6609|false|false|false|C0332290|Consistent with|CONSISTENT
Anatomy|Body System|General Exam|6616,6620|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|General Exam|6616,6620|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|General Exam|6616,6620|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|General Exam|6616,6620|false|false|false|||SKIN
Finding|Body Substance|General Exam|6616,6620|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|General Exam|6616,6620|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Event|Event|General Exam|6630,6631|false|false|false|||/
Anatomy|Body Part, Organ, or Organ Component|General Exam|6634,6641|false|false|false|C0017420;C0559522|Genital system;Genitalia|GENITAL
Anatomy|Body System|General Exam|6634,6641|false|false|false|C0017420;C0559522|Genital system;Genitalia|GENITAL
Finding|Body Substance|General Exam|6634,6641|false|false|false|C1546649;C1550642|Specimen Type - Genital|GENITAL
Finding|Intellectual Product|General Exam|6634,6641|false|false|false|C1546649;C1550642|Specimen Type - Genital|GENITAL
Event|Event|General Exam|6642,6655|false|false|false|||CONTAMINATION
Finding|Idea or Concept|General Exam|6642,6655|false|false|false|C2349974|Contamination|CONTAMINATION
Phenomenon|Human-caused Phenomenon or Process|General Exam|6642,6655|false|false|false|C0259846|adulteration|CONTAMINATION
Event|Event|General Exam|6677,6679|false|false|false|||SP
Finding|Functional Concept|General Exam|6735,6744|false|false|false|C1285553|Interprets|INTERPRET
Event|Event|General Exam|6745,6752|false|false|false|||RESULTS
Event|Event|General Exam|6758,6765|false|false|false|||CAUTION
Event|Event|General Exam|6799,6812|false|false|false|||SENSITIVITIES
Finding|Finding|General Exam|6799,6812|false|false|false|C0427965|Antimicrobial susceptibility|SENSITIVITIES
Disorder|Neoplastic Process|General Exam|6814,6817|false|false|false|C2732473|Ductal Carcinoma In Situ with Microinvasion|MIC
Drug|Hazardous or Poisonous Substance|General Exam|6814,6817|false|false|false|C0066256|methyl isocyanate|MIC
Drug|Organic Chemical|General Exam|6814,6817|false|false|false|C0066256|methyl isocyanate|MIC
Event|Event|General Exam|6814,6817|false|false|false|||MIC
Procedure|Laboratory Procedure|General Exam|6814,6817|false|false|false|C0281162;C0427978|Minimum Inhibitory Concentration Test;cisplatin/ifosfamide/mitomycin protocol|MIC
Procedure|Therapeutic or Preventive Procedure|General Exam|6814,6817|false|false|false|C0281162;C0427978|Minimum Inhibitory Concentration Test;cisplatin/ifosfamide/mitomycin protocol|MIC
Event|Event|General Exam|6832,6835|false|false|false|||MCG
Event|Event|General Exam|6962,6964|false|false|false|||SP
Drug|Antibiotic|General Exam|7000,7010|false|false|false|C0002680;C2095775|ampicillin;ampicillins|AMPICILLIN
Drug|Organic Chemical|General Exam|7000,7010|false|false|false|C0002680;C2095775|ampicillin;ampicillins|AMPICILLIN
Drug|Organic Chemical|General Exam|7031,7045|false|false|false|C0028156|nitrofurantoin|NITROFURANTOIN
Drug|Pharmacologic Substance|General Exam|7031,7045|false|false|false|C0028156|nitrofurantoin|NITROFURANTOIN
Disorder|Injury or Poisoning|General Exam|7062,7074|false|false|false|C0481114|Tetracyclines causing adverse effects in therapeutic use|TETRACYCLINE
Drug|Antibiotic|General Exam|7062,7074|false|false|false|C0039644;C1744619|Tetracycline Antibiotics;tetracycline|TETRACYCLINE
Drug|Organic Chemical|General Exam|7062,7074|false|false|false|C0039644;C1744619|Tetracycline Antibiotics;tetracycline|TETRACYCLINE
Event|Event|General Exam|7062,7074|false|false|false|||TETRACYCLINE
Drug|Amino Acid, Peptide, or Protein|General Exam|7093,7103|false|false|false|C0042313|vancomycin|VANCOMYCIN
Drug|Antibiotic|General Exam|7093,7103|false|false|false|C0042313|vancomycin|VANCOMYCIN
Event|Event|General Exam|7093,7103|false|false|false|||VANCOMYCIN
Procedure|Laboratory Procedure|General Exam|7093,7103|false|false|false|C0489941|Vancomycin measurement|VANCOMYCIN
Event|Event|General Exam|7125,7132|false|false|false|||IMAGING
Finding|Finding|General Exam|7125,7132|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|General Exam|7125,7132|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Event|Event|General Exam|7164,7167|false|false|false|||CXR
Procedure|Diagnostic Procedure|General Exam|7164,7167|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|General Exam|7168,7178|false|false|false|||IMPRESSION
Finding|Intellectual Product|General Exam|7168,7178|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|General Exam|7168,7178|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Event|Event|General Exam|7186,7196|true|false|false|||congestion
Finding|Pathologic Function|General Exam|7186,7196|true|false|false|C0700148|Congestion|congestion
Disorder|Disease or Syndrome|General Exam|7205,7210|true|false|false|C0398650|Immune thrombocytopenic purpura|frank
Attribute|Clinical Attribute|General Exam|7211,7216|true|false|false|C1717255||edema
Event|Event|General Exam|7211,7216|true|false|false|||edema
Finding|Pathologic Function|General Exam|7211,7216|true|false|false|C0013604|Edema|edema
Event|Event|General Exam|7234,7239|true|false|false|||signs
Finding|Finding|General Exam|7234,7239|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|General Exam|7234,7239|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Disorder|Disease or Syndrome|General Exam|7243,7252|true|false|false|C0032285|Pneumonia|pneumonia
Event|Event|General Exam|7243,7252|true|false|false|||pneumonia
Drug|Amino Acid, Peptide, or Protein|General Exam|7259,7262|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|General Exam|7259,7262|false|false|false|||CTA
Finding|Gene or Genome|General Exam|7259,7262|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|General Exam|7259,7262|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Anatomy|Body Location or Region|General Exam|7263,7268|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|General Exam|7263,7268|false|false|false|C0741025|Chest problem|chest
Event|Event|General Exam|7269,7275|false|false|false|||showed
Anatomy|Body Part, Organ, or Organ Component|General Exam|7290,7299|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|General Exam|7290,7299|false|false|false|C2707265||pulmonary
Finding|Finding|General Exam|7290,7299|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|General Exam|7290,7308|false|false|false|C0034065|Pulmonary Embolism|pulmonary embolism
Event|Event|General Exam|7300,7308|false|false|false|||embolism
Finding|Finding|General Exam|7300,7308|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Finding|Pathologic Function|General Exam|7300,7308|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Event|Event|General Exam|7314,7322|false|false|false|||thrombus
Finding|Pathologic Function|General Exam|7314,7322|false|false|false|C0087086;C0302148|Blood Clot;Thrombus|thrombus
Event|Event|General Exam|7323,7327|false|false|false|||seen
Event|Event|General Exam|7328,7337|false|false|false|||extending
Finding|Functional Concept|General Exam|7348,7353|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|General Exam|7348,7375|false|false|false|C0226054;C0923924|Right pulmonary arterial tree;Right pulmonary artery|right main pulmonary artery
Anatomy|Body Part, Organ, or Organ Component|General Exam|7359,7368|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|General Exam|7359,7368|false|false|false|C2707265||pulmonary
Finding|Finding|General Exam|7359,7368|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Anatomy|Body Part, Organ, or Organ Component|General Exam|7359,7375|false|false|false|C0034052|Pulmonary artery structure|pulmonary artery
Anatomy|Body Part, Organ, or Organ Component|General Exam|7369,7375|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|General Exam|7369,7375|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Finding|Functional Concept|General Exam|7413,7418|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Event|Event|General Exam|7426,7432|false|false|false|||middle
Finding|Intellectual Product|General Exam|7426,7432|false|false|false|C1552826|Table Cell Vertical Align - middle|middle
Anatomy|Body Location or Region|General Exam|7438,7443|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|7438,7443|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|General Exam|7438,7448|false|false|false|C0225758|Structure of lower lobe of lung|lower lobe
Anatomy|Body Part, Organ, or Organ Component|General Exam|7444,7448|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|General Exam|7444,7448|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Anatomy|Body Part, Organ, or Organ Component|General Exam|7444,7458|false|false|false|C0225752|Structure of lobe of lung|lobe pulmonary
Anatomy|Body Part, Organ, or Organ Component|General Exam|7449,7458|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|General Exam|7449,7458|false|false|false|C2707265||pulmonary
Finding|Finding|General Exam|7449,7458|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Anatomy|Body Part, Organ, or Organ Component|General Exam|7460,7468|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Anatomy|Body System|General Exam|7460,7468|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Event|Event|General Exam|7460,7468|false|false|false|||arteries
Procedure|Health Care Activity|General Exam|7460,7468|false|false|false|C0397581|Procedure on artery|arteries
Finding|Functional Concept|General Exam|7473,7478|true|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|General Exam|7473,7484|true|false|false|C0225808|Right side of heart|right heart
Anatomy|Body Part, Organ, or Organ Component|General Exam|7479,7484|true|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|General Exam|7479,7484|true|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|General Exam|7479,7484|true|false|false|C0795691|HEART PROBLEM|heart
Disorder|Injury or Poisoning|General Exam|7485,7491|true|false|false|C0080194|Muscle strain|strain
Event|Event|General Exam|7485,7491|true|false|false|||strain
Finding|Idea or Concept|General Exam|7485,7491|true|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Finding|Mental Process|General Exam|7485,7491|true|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Finding|Physiologic Function|General Exam|7485,7491|true|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Finding|Sign or Symptom|General Exam|7485,7491|true|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Event|Event|General Exam|7492,7502|true|false|false|||identified
Anatomy|Body Part, Organ, or Organ Component|General Exam|7540,7549|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|General Exam|7540,7549|false|false|false|C2707265||pulmonary
Finding|Finding|General Exam|7540,7549|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|General Exam|7540,7556|false|false|false|C0034065|Pulmonary Embolism|pulmonary emboli
Event|Event|General Exam|7550,7556|false|false|false|||emboli
Finding|Finding|General Exam|7550,7556|false|false|false|C1704212|Embolus|emboli
Event|Event|General Exam|7557,7561|false|false|false|||seen
Event|Event|General Exam|7597,7605|false|false|false|||branches
Finding|Functional Concept|General Exam|7613,7617|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|General Exam|7628,7633|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|7628,7633|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|General Exam|7634,7639|false|false|false|C0796494|lobe|lobes
Anatomy|Body Part, Organ, or Organ Component|General Exam|7653,7662|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|General Exam|7653,7662|false|false|false|C2707265||pulmonary
Finding|Finding|General Exam|7653,7662|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Finding|General Exam|7653,7670|false|false|false|C0748164|Multiple Pulmonary Nodules|pulmonary nodules
Event|Event|General Exam|7663,7670|false|false|false|||nodules
Event|Event|General Exam|7675,7680|false|false|false|||noted
Event|Event|General Exam|7685,7690|false|false|false|||noted
Event|Event|General Exam|7731,7741|false|false|false|||spiculated
Event|Event|General Exam|7746,7755|false|false|false|||measuring
Finding|Functional Concept|General Exam|7775,7780|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|General Exam|7775,7792|false|false|false|C4281590|Structure of middle lobe of right lung|right middle lobe
Finding|Intellectual Product|General Exam|7781,7787|false|false|false|C1552826|Table Cell Vertical Align - middle|middle
Anatomy|Body Part, Organ, or Organ Component|General Exam|7781,7792|false|false|false|C4281590|Structure of middle lobe of right lung|middle lobe
Anatomy|Body Part, Organ, or Organ Component|General Exam|7788,7792|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|General Exam|7788,7792|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Event|Event|General Exam|7794,7804|false|false|false|||suspicious
Finding|Finding|General Exam|7794,7819|false|false|false|C4050405|Suspicious for Malignancy|suspicious for malignancy
Disorder|Neoplastic Process|General Exam|7809,7819|false|true|false|C0006826;C1306459|Malignant Neoplasms;Primary malignant neoplasm|malignancy
Event|Event|General Exam|7809,7819|false|false|false|||malignancy
Procedure|Diagnostic Procedure|General Exam|7837,7840|false|false|false|C0032743;C0040398|Positron-Emission Tomography;Tomography, Emission-Computed|PET
Procedure|Diagnostic Procedure|General Exam|7837,7843|false|false|false|C1699633|PET/CT scan|PET-CT
Event|Event|General Exam|7841,7843|false|false|false|||CT
Event|Event|General Exam|7852,7865|false|false|false|||demonstration
Finding|Functional Concept|General Exam|7871,7875|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|General Exam|7871,7882|false|false|false|C0222601|Left breast|left breast
Anatomy|Body Part, Organ, or Organ Component|General Exam|7876,7882|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|General Exam|7876,7882|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Finding|Finding|General Exam|7876,7882|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|General Exam|7876,7882|false|false|false|C0191838|Procedures on breast|breast
Finding|Finding|General Exam|7876,7890|false|false|false|C0024103|Mass in breast|breast nodules
Event|Event|General Exam|7883,7890|false|false|false|||nodules
Event|Event|General Exam|7902,7913|false|false|false|||correlation
Event|Event|General Exam|7919,7930|false|false|false|||mammography
Procedure|Diagnostic Procedure|General Exam|7919,7930|false|false|false|C0024671;C0848600|Mammography;Mammography, Female|mammography
Event|Event|General Exam|7935,7945|false|false|false|||ultrasound
Finding|Functional Concept|General Exam|7935,7945|false|false|false|C0220934|Ultrasonic|ultrasound
Phenomenon|Natural Phenomenon or Process|General Exam|7935,7945|false|false|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|ultrasound
Procedure|Diagnostic Procedure|General Exam|7935,7945|false|false|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|ultrasound
Event|Event|General Exam|7949,7958|false|false|false|||suggested
Finding|Intellectual Product|Impression|7985,7993|false|false|false|C1552654|Parameterized Data Type - Interval|Interval
Event|Event|Impression|7994,8005|false|false|false|||progression
Finding|Functional Concept|Impression|7994,8005|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Finding|Pathologic Function|Impression|7994,8005|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Attribute|Clinical Attribute|Impression|8009,8013|false|false|false|C4318566|Deep Resection Margin|deep
Anatomy|Body Part, Organ, or Organ Component|Impression|8009,8018|false|false|false|C0226514|Structure of deep vein|deep vein
Disorder|Disease or Syndrome|Impression|8009,8029|false|false|false|C0149871;C0340708|Deep Vein Thrombosis;Deep vein thrombosis of lower limb|deep vein thrombosis
Anatomy|Body Part, Organ, or Organ Component|Impression|8014,8018|false|false|false|C0042449|Veins|vein
Finding|Pathologic Function|Impression|8014,8029|false|false|false|C0042487|Venous Thrombosis|vein thrombosis
Event|Event|Impression|8019,8029|false|false|false|||thrombosis
Finding|Pathologic Function|Impression|8019,8029|false|false|false|C0040053|Thrombosis|thrombosis
Finding|Functional Concept|Impression|8037,8041|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|Impression|8043,8048|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|Impression|8043,8048|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|Impression|8043,8058|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|Impression|8049,8058|false|false|false|C0015385|Limb structure|extremity
Finding|Functional Concept|Impression|8065,8074|false|false|false|C1947917|Occluded|occlusive
Disorder|Acquired Abnormality|Impression|8065,8083|false|false|false|C0333203|Occlusive thrombus|occlusive thrombus
Event|Event|Impression|8075,8083|false|false|false|||thrombus
Finding|Pathologic Function|Impression|8075,8083|false|false|false|C0087086;C0302148|Blood Clot;Thrombus|thrombus
Event|Event|Impression|8084,8093|false|false|false|||involving
Anatomy|Body Part, Organ, or Organ Component|Impression|8106,8113|false|false|false|C0015811|Femur|femoral
Anatomy|Body Part, Organ, or Organ Component|Impression|8106,8118|false|false|false|C0015809|Femoral vein|femoral vein
Anatomy|Body Part, Organ, or Organ Component|Impression|8114,8118|false|false|false|C0042449|Veins|vein
Event|Event|Impression|8136,8145|false|false|false|||involving
Attribute|Clinical Attribute|Impression|8158,8164|false|false|false|C4522154|Distal Resection Margin|distal
Anatomy|Body Part, Organ, or Organ Component|Impression|8166,8173|false|false|false|C0015811|Femur|femoral
Anatomy|Body Part, Organ, or Organ Component|Impression|8166,8178|false|false|false|C0015809|Femoral vein|femoral vein
Anatomy|Body Part, Organ, or Organ Component|Impression|8174,8178|false|false|false|C0042449|Veins|vein
Finding|Functional Concept|Impression|8190,8200|false|false|false|C1524062|Additional|additional
Event|Event|Impression|8214,8222|false|false|false|||thrombus
Finding|Pathologic Function|Impression|8214,8222|false|false|false|C0087086;C0302148|Blood Clot;Thrombus|thrombus
Attribute|Clinical Attribute|Impression|8231,8235|false|false|false|C4318566|Deep Resection Margin|deep
Anatomy|Body Part, Organ, or Organ Component|Impression|8231,8248|false|false|false|C0226841|Structure of profunda femoris vein|deep femoral vein
Anatomy|Body Part, Organ, or Organ Component|Impression|8236,8243|false|false|false|C0015811|Femur|femoral
Anatomy|Body Part, Organ, or Organ Component|Impression|8236,8248|false|false|false|C0015809|Femoral vein|femoral vein
Anatomy|Body Part, Organ, or Organ Component|Impression|8244,8248|false|false|false|C0042449|Veins|vein
Finding|Functional Concept|Impression|8255,8259|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Functional Concept|Impression|8260,8266|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Finding|Intellectual Product|Impression|8260,8266|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Anatomy|Body Part, Organ, or Organ Component|Impression|8267,8274|false|false|false|C0015811|Femur|femoral
Anatomy|Body Location or Region|Impression|8279,8288|false|false|false|C0442037|popliteal|popliteal
Anatomy|Body Part, Organ, or Organ Component|Impression|8279,8294|false|false|false|C0032652|Structure of popliteal vein|popliteal veins
Anatomy|Body Part, Organ, or Organ Component|Impression|8289,8294|false|false|false|C0042449|Veins|veins
Procedure|Therapeutic or Preventive Procedure|Impression|8289,8294|false|false|false|C0398102|Procedure on vein|veins
Event|Event|Impression|8300,8306|false|false|false|||patent
Finding|Intellectual Product|Impression|8300,8306|false|false|false|C0030650|Legal patent|patent
Anatomy|Body Location or Region|Impression|8325,8329|true|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|Impression|8325,8329|true|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|Impression|8330,8335|true|false|false|C0042449|Veins|veins
Event|Event|Impression|8330,8335|true|false|false|||veins
Procedure|Therapeutic or Preventive Procedure|Impression|8330,8335|true|false|false|C0398102|Procedure on vein|veins
Event|Event|Impression|8345,8355|true|false|false|||visualized
Event|Event|Impression|8367,8376|true|false|false|||overlying
Drug|Biomedical or Dental Material|Impression|8377,8385|true|false|false|C1705365|Dressing Dosage Form|dressing
Event|Event|Impression|8377,8385|true|false|false|||dressing
Finding|Daily or Recreational Activity|Impression|8377,8385|true|false|false|C0518459;C1305428|Ability to dress|dressing
Finding|Finding|Impression|8377,8385|true|false|false|C0518459;C1305428|Ability to dress|dressing
Procedure|Health Care Activity|Impression|8377,8385|true|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Procedure|Therapeutic or Preventive Procedure|Impression|8377,8385|true|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Event|Event|Impression|8400,8408|true|false|false|||evidence
Finding|Idea or Concept|Impression|8400,8408|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Impression|8400,8411|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Attribute|Clinical Attribute|Impression|8412,8416|true|false|false|C4318566|Deep Resection Margin|deep
Anatomy|Body Part, Organ, or Organ Component|Impression|8417,8423|true|false|false|C0042449|Veins|venous
Event|Event|Impression|8425,8435|true|false|false|||thrombosis
Finding|Pathologic Function|Impression|8425,8435|true|false|false|C0040053|Thrombosis|thrombosis
Finding|Functional Concept|Impression|8443,8448|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|Impression|8443,8464|false|false|false|C0230415|Right lower extremity|right lower extremity
Anatomy|Body Location or Region|Impression|8449,8454|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|Impression|8449,8454|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|Impression|8449,8464|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|Impression|8455,8464|false|false|false|C0015385|Limb structure|extremity
Event|Event|Impression|8471,8474|false|false|false|||TTE
Procedure|Diagnostic Procedure|Impression|8471,8474|false|false|false|C0430462|Transthoracic echocardiography|TTE
Event|Event|Impression|8476,8487|false|false|false|||Conclusions
Finding|Idea or Concept|Impression|8476,8487|false|false|false|C1707478|Conclusion|Conclusions
Finding|Functional Concept|Impression|8492,8496|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Impression|8492,8503|false|false|false|C0225860|Left atrial structure|left atrium
Anatomy|Body Part, Organ, or Organ Component|Impression|8497,8503|false|false|false|C0018792|Heart Atrium|atrium
Event|Event|Impression|8507,8513|false|false|false|||normal
Finding|Functional Concept|Impression|8537,8542|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|Impression|8543,8549|false|false|false|C0018792|Heart Atrium|atrial
Event|Event|Impression|8551,8559|false|false|false|||pressure
Finding|Finding|Impression|8551,8559|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|Impression|8551,8559|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|Impression|8551,8559|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|Impression|8551,8559|false|false|false|C0033095||pressure
Finding|Functional Concept|Impression|8573,8577|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|Impression|8573,8594|false|false|false|C0504053|Wall of left ventricle|Left ventricular wall
Anatomy|Body Part, Organ, or Organ Component|Impression|8578,8589|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Part, Organ, or Organ Component|Impression|8578,8594|false|false|false|C0507618|Wall of ventricle|ventricular wall
Finding|Finding|Impression|8578,8604|false|false|false|C2024242|cardiac evaluation of ventricular wall thickness|ventricular wall thickness
Event|Event|Impression|8595,8604|false|false|false|||thickness
Anatomy|Body Space or Junction|Impression|8606,8612|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|Impression|8606,8612|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|Impression|8606,8612|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Finding|Organ or Tissue Function|Impression|8631,8639|false|false|false|C0039155|Systole|systolic
Event|Event|Impression|8640,8648|false|false|false|||function
Finding|Finding|Impression|8640,8648|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|Impression|8640,8648|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|Impression|8640,8648|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|Impression|8640,8648|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Event|Event|Impression|8653,8659|false|false|false|||normal
Attribute|Clinical Attribute|Impression|8661,8665|false|false|false|C0428772|Left ventricular ejection fraction|LVEF
Event|Event|Impression|8661,8665|false|false|false|||LVEF
Procedure|Diagnostic Procedure|Impression|8661,8665|false|false|false|C3837267|LVEF (procedure)|LVEF
Procedure|Diagnostic Procedure|Impression|8673,8680|false|false|false|C0554756|Doppler studies|Doppler
Event|Event|Impression|8681,8691|false|false|false|||parameters
Finding|Finding|Impression|8681,8691|false|false|false|C0449381|Observation parameter|parameters
Event|Event|Impression|8701,8711|false|false|false|||consistent
Finding|Idea or Concept|Impression|8701,8711|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|Impression|8701,8716|false|false|false|C0332290|Consistent with|consistent with
Finding|Classification|Impression|8712,8722|false|false|false|C0441800|Grade|with Grade
Finding|Classification|Impression|8717,8722|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|Grade
Finding|Finding|Impression|8717,8722|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|Grade
Finding|Finding|Impression|8717,8724|false|false|false|C0475269;C0687695;C4049998|Clavien-Dindo Grade I;Grade 1 (qualifier value);Tumor grade G1|Grade I
Finding|Intellectual Product|Impression|8717,8724|false|false|false|C0475269;C0687695;C4049998|Clavien-Dindo Grade I;Grade 1 (qualifier value);Tumor grade G1|Grade I
Finding|Intellectual Product|Impression|8726,8730|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Functional Concept|Impression|8732,8736|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Impression|8738,8749|false|false|false|C0018827|Heart Ventricle|ventricular
Attribute|Clinical Attribute|Impression|8750,8759|false|false|false|C0012000|Diastole|diastolic
Finding|Pathologic Function|Impression|8750,8771|false|false|false|C0520863|Diastolic dysfunction|diastolic dysfunction
Disorder|Disease or Syndrome|Impression|8760,8771|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Event|Event|Impression|8760,8771|false|false|false|||dysfunction
Finding|Conceptual Entity|Impression|8760,8771|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|Impression|8760,8771|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|Impression|8760,8771|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|Impression|8773,8778|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Part, Organ, or Organ Component|Impression|8779,8790|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Part, Organ, or Organ Component|Impression|8791,8798|false|false|false|C0935616|chamber [body part]|chamber
Event|Event|Impression|8809,8813|false|false|false|||free
Finding|Functional Concept|Impression|8809,8813|false|false|false|C0332296|Free of (attribute)|free
Attribute|Clinical Attribute|Impression|8814,8825|false|false|false|C1980023|Wall motion|wall motion
Event|Event|Impression|8819,8825|false|false|false|||motion
Phenomenon|Natural Phenomenon or Process|Impression|8819,8825|false|false|false|C0026597|Motion|motion
Event|Event|Impression|8830,8836|false|false|false|||normal
Anatomy|Body Part, Organ, or Organ Component|Impression|8842,8848|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|Impression|8842,8854|false|false|false|C0003501;C4533215|Aortic valve structure;Chest>Aortic valve|aortic valve
Anatomy|Body Part, Organ, or Organ Component|Impression|8849,8854|false|false|false|C1186983|Anatomical valve|valve
Event|Event|Impression|8876,8885|false|false|false|||thickened
Anatomy|Body Part, Organ, or Organ Component|Impression|8904,8910|true|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|Impression|8904,8916|true|false|false|C0003501;C4533215|Aortic valve structure;Chest>Aortic valve|aortic valve
Disorder|Congenital Abnormality|Impression|8904,8925|true|false|false|C5193127;C5700069|AORTIC VALVE DISEASE 3;Stenosis of aorta|aortic valve stenosis
Disorder|Disease or Syndrome|Impression|8904,8925|true|false|false|C5193127;C5700069|AORTIC VALVE DISEASE 3;Stenosis of aorta|aortic valve stenosis
Finding|Pathologic Function|Impression|8904,8925|true|false|false|C0003507|Aortic Valve Stenosis|aortic valve stenosis
Anatomy|Body Part, Organ, or Organ Component|Impression|8911,8916|true|false|false|C1186983|Anatomical valve|valve
Event|Event|Impression|8917,8925|true|false|false|||stenosis
Finding|Pathologic Function|Impression|8917,8925|true|false|false|C1261287|Stenosis|stenosis
Disorder|Disease or Syndrome|Impression|8936,8956|false|false|false|C0026266|Mitral Valve Insufficiency|mitral regurgitation
Event|Event|Impression|8943,8956|false|false|false|||regurgitation
Finding|Finding|Impression|8943,8956|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|Impression|8943,8956|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|Impression|8943,8956|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Event|Event|Impression|8960,8964|false|false|false|||seen
Finding|Intellectual Product|Impression|8975,8979|false|false|false|C1547225|Mild Severity of Illness Code|mild
Anatomy|Body Part, Organ, or Organ Component|Impression|8980,8989|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Impression|8980,8989|false|false|false|C2707265||pulmonary
Finding|Finding|Impression|8980,8989|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Anatomy|Body Part, Organ, or Organ Component|Impression|8991,8997|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|Impression|8991,8997|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Finding|Organ or Tissue Function|Impression|8998,9006|false|false|false|C0039155|Systole|systolic
Disorder|Disease or Syndrome|Impression|8998,9019|false|false|false|C0221155|Systolic Hypertension|systolic hypertension
Disorder|Disease or Syndrome|Impression|9007,9019|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|Impression|9007,9019|false|false|false|||hypertension
Event|Event|Impression|9027,9030|false|false|false|||CXR
Procedure|Diagnostic Procedure|Impression|9027,9030|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|Impression|9044,9052|false|false|false|||Compared
Anatomy|Body Location or Region|Impression|9056,9061|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Impression|9056,9061|false|false|false|C0741025|Chest problem|chest
Event|Event|Impression|9062,9073|false|false|false|||radiographs
Procedure|Diagnostic Procedure|Impression|9062,9073|false|false|false|C1306645|Plain x-ray|radiographs
Anatomy|Body Part, Organ, or Organ Component|Impression|9092,9097|false|false|false|C0018787;C4037974|Chest>Heart;Heart|Heart
Disorder|Neoplastic Process|Impression|9092,9097|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|Heart
Finding|Sign or Symptom|Impression|9092,9097|false|false|false|C0795691|HEART PROBLEM|Heart
Finding|Finding|Impression|9092,9102|false|false|false|C0744689|heart size|Heart size
Anatomy|Body Part, Organ, or Organ Component|Impression|9116,9121|false|false|false|C0024109|Lung|Lungs
Event|Event|Impression|9130,9135|false|false|false|||clear
Finding|Idea or Concept|Impression|9130,9135|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Tissue|Impression|9141,9148|true|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|Impression|9141,9148|true|false|false|C0032226|Pleural Diseases|pleural
Disorder|Congenital Abnormality|Impression|9150,9161|true|false|false|C0000768|Congenital Abnormality|abnormality
Event|Event|Impression|9150,9161|true|false|false|||abnormality
Finding|Finding|Impression|9150,9161|true|false|false|C1704258|Abnormality|abnormality
Event|Event|Impression|9165,9173|true|false|false|||evidence
Finding|Idea or Concept|Impression|9165,9173|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Impression|9165,9176|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Drug|Pharmacologic Substance|Impression|9177,9184|true|false|false|C0719205|Central brand of multivitamin with minerals|central
Drug|Vitamin|Impression|9177,9184|true|false|false|C0719205|Central brand of multivitamin with minerals|central
Event|Event|Impression|9177,9184|true|false|false|||central
Procedure|Laboratory Procedure|Impression|9177,9184|true|false|false|C1879652|Central Minus|central
Finding|Body Substance|Impression|9177,9190|true|false|false|C1179479|Central lymph|central lymph
Finding|Body Substance|Impression|9185,9190|false|false|false|C0024202|Lymph|lymph
Anatomy|Body Part, Organ, or Organ Component|Impression|9185,9195|false|false|false|C0024204|lymph nodes|lymph node
Disorder|Disease or Syndrome|Impression|9185,9207|false|false|false|C0497156|Lymphadenopathy|lymph node enlargement
Finding|Sign or Symptom|Impression|9185,9207|false|false|false|C4282165|Swollen Lymph Node|lymph node enlargement
Disorder|Anatomical Abnormality|Impression|9196,9207|false|false|false|C2711450|Enlargement (morphologic abnormality)|enlargement
Event|Event|Impression|9196,9207|false|false|false|||enlargement
Finding|Pathologic Function|Impression|9196,9207|false|false|false|C0020564|Hypertrophy|enlargement
Procedure|Therapeutic or Preventive Procedure|Impression|9196,9207|false|false|false|C1293134|Enlargement procedure|enlargement
Drug|Chemical Viewed Structurally|Hospital Course|9270,9277|false|false|false|C0302912|Radicals (chemistry)|radical
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9270,9288|false|false|false|C0194401|Complete cystectomy|radical cystectomy
Event|Event|Hospital Course|9278,9288|false|false|false|||cystectomy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9278,9288|false|false|false|C0010651|Cystectomy|cystectomy
Event|Event|Hospital Course|9293,9303|false|false|false|||omplicated
Finding|Finding|Hospital Course|9307,9317|false|false|false|C0004610|Bacteremia|bacteremia
Disorder|Disease or Syndrome|Hospital Course|9323,9330|false|false|false|C0000833|Abscess|abscess
Event|Event|Hospital Course|9323,9330|false|false|false|||abscess
Finding|Intellectual Product|Hospital Course|9323,9330|false|false|false|C1546533||abscess
Event|Event|Hospital Course|9332,9335|false|false|false|||LLE
Anatomy|Body Location or Region|Hospital Course|9336,9339|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Hospital Course|9336,9339|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Hospital Course|9336,9339|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|Hospital Course|9336,9339|false|false|false|||DVT
Drug|Organic Chemical|Hospital Course|9360,9367|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|Hospital Course|9360,9367|false|false|false|C0728963|Lovenox|lovenox
Event|Event|Hospital Course|9360,9367|false|false|false|||lovenox
Event|Event|Hospital Course|9372,9380|false|false|false|||presents
Event|Event|Hospital Course|9387,9394|false|false|false|||dyspnea
Finding|Finding|Hospital Course|9387,9394|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|Hospital Course|9387,9394|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|Hospital Course|9387,9406|false|false|false|C0231807|Dyspnea on exertion|dyspnea on exertion
Event|Event|Hospital Course|9398,9406|false|false|false|||exertion
Finding|Organism Function|Hospital Course|9398,9406|false|false|false|C0015264|Exertion|exertion
Event|Event|Hospital Course|9411,9418|false|false|false|||dyspnea
Finding|Finding|Hospital Course|9411,9418|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|Hospital Course|9411,9418|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|Hospital Course|9411,9430|false|false|false|C0231807|Dyspnea on exertion|dyspnea on exertion
Event|Event|Hospital Course|9422,9430|false|false|false|||exertion
Finding|Organism Function|Hospital Course|9422,9430|false|false|false|C0015264|Exertion|exertion
Event|Event|Hospital Course|9435,9440|false|false|false|||found
Finding|Gene or Genome|Hospital Course|9450,9455|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Event|Event|Hospital Course|9463,9474|false|false|false|||progression
Finding|Functional Concept|Hospital Course|9463,9474|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Finding|Pathologic Function|Hospital Course|9463,9474|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Anatomy|Body Location or Region|Hospital Course|9478,9481|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Hospital Course|9478,9481|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Hospital Course|9478,9481|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|Hospital Course|9478,9481|false|false|false|||DVT
Anatomy|Body Location or Region|Hospital Course|9489,9492|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Hospital Course|9489,9492|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Hospital Course|9489,9492|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Finding|Finding|Hospital Course|9494,9500|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Idea or Concept|Hospital Course|9494,9500|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Event|Event|Hospital Course|9501,9504|false|false|false|||due
Finding|Functional Concept|Hospital Course|9501,9504|false|true|false|C0678226;C3146286|Due;Due to|due
Finding|Idea or Concept|Hospital Course|9501,9504|false|true|false|C0678226;C3146286|Due;Due to|due
Finding|Functional Concept|Hospital Course|9501,9507|false|true|false|C0678226|Due to|due to
Event|Event|Hospital Course|9508,9522|false|false|false|||undertreatment
Procedure|Health Care Activity|Hospital Course|9508,9522|false|true|false|C5828474|Undertreatment|undertreatment
Anatomy|Body Location or Region|Hospital Course|9536,9539|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Hospital Course|9536,9539|false|true|false|C2926618||DVT
Disorder|Disease or Syndrome|Hospital Course|9536,9539|false|true|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|Hospital Course|9536,9539|false|false|false|||DVT
Drug|Pharmacologic Substance|Hospital Course|9546,9558|false|false|false|C0355642|Drugs used in migraine prophylaxis|prophylactic
Event|Event|Hospital Course|9546,9558|false|false|false|||prophylactic
Finding|Functional Concept|Hospital Course|9546,9558|false|false|false|C0445202|Prophylactic behavior|prophylactic
Event|Event|Hospital Course|9559,9565|false|false|false|||dosing
Drug|Organic Chemical|Hospital Course|9569,9576|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|Hospital Course|9569,9576|false|false|false|C0728963|Lovenox|lovenox
Event|Event|Hospital Course|9569,9576|false|false|false|||lovenox
Event|Event|Hospital Course|9584,9595|true|false|false|||underdosing
Drug|Organic Chemical|Hospital Course|9599,9606|true|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|Hospital Course|9599,9606|true|false|false|C0728963|Lovenox|lovenox
Event|Event|Hospital Course|9599,9606|true|false|false|||lovenox
Event|Event|Hospital Course|9622,9629|true|false|false|||thought
Event|Event|Hospital Course|9636,9645|true|false|false|||treatment
Finding|Conceptual Entity|Hospital Course|9636,9645|true|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Hospital Course|9636,9645|true|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Hospital Course|9636,9645|true|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9636,9645|true|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Finding|Finding|Hospital Course|9636,9653|true|false|false|C0162643;C0438286;C1547544|Absent response to treatment;Charge Type Reason - Treatment Failure;treatment failure|treatment failure
Finding|Idea or Concept|Hospital Course|9636,9653|true|false|false|C0162643;C0438286;C1547544|Absent response to treatment;Charge Type Reason - Treatment Failure;treatment failure|treatment failure
Event|Event|Hospital Course|9646,9653|true|false|false|||failure
Finding|Functional Concept|Hospital Course|9646,9653|true|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|Hospital Course|9646,9653|true|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|Hospital Course|9646,9653|true|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9658,9661|true|false|false|C3498924|lamina IVC|IVC
Procedure|Diagnostic Procedure|Hospital Course|9658,9661|true|false|false|C4085887|Inspiratory Vital Capacity Test|IVC
Event|Event|Hospital Course|9662,9668|false|false|false|||filter
Finding|Body Substance|Hospital Course|9662,9668|false|false|false|C1522664;C1546637;C1550638;C1704449|Filter (function);Specimen Type - Filter;filter information process|filter
Finding|Conceptual Entity|Hospital Course|9662,9668|false|false|false|C1522664;C1546637;C1550638;C1704449|Filter (function);Specimen Type - Filter;filter information process|filter
Finding|Intellectual Product|Hospital Course|9662,9668|false|false|false|C1522664;C1546637;C1550638;C1704449|Filter (function);Specimen Type - Filter;filter information process|filter
Event|Event|Hospital Course|9674,9682|false|false|false|||deferred
Event|Event|Hospital Course|9695,9700|true|false|false|||signs
Finding|Finding|Hospital Course|9695,9700|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Hospital Course|9695,9700|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Hospital Course|9704,9709|true|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|Hospital Course|9704,9715|true|false|false|C0225808|Right side of heart|right heart
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9710,9715|true|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Hospital Course|9710,9715|true|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Hospital Course|9710,9715|true|false|false|C0795691|HEART PROBLEM|heart
Disorder|Injury or Poisoning|Hospital Course|9716,9722|true|false|false|C0080194|Muscle strain|strain
Event|Event|Hospital Course|9716,9722|true|false|false|||strain
Finding|Idea or Concept|Hospital Course|9716,9722|true|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Finding|Mental Process|Hospital Course|9716,9722|true|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Finding|Physiologic Function|Hospital Course|9716,9722|true|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Finding|Sign or Symptom|Hospital Course|9716,9722|true|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Event|Event|Hospital Course|9726,9733|true|false|false|||imaging
Finding|Finding|Hospital Course|9726,9733|true|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|Hospital Course|9726,9733|true|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Event|Event|Hospital Course|9736,9739|false|false|false|||EKG
Finding|Intellectual Product|Hospital Course|9736,9739|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|Hospital Course|9736,9739|false|false|false|C1623258|Electrocardiography|EKG
Event|Event|Hospital Course|9741,9745|false|false|false|||exam
Finding|Functional Concept|Hospital Course|9741,9745|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|Hospital Course|9741,9745|false|false|false|C0582103|Medical Examination|exam
Event|Event|Hospital Course|9747,9750|true|false|false|||TTE
Procedure|Diagnostic Procedure|Hospital Course|9747,9750|true|false|false|C0430462|Transthoracic echocardiography|TTE
Event|Event|Hospital Course|9751,9757|true|false|false|||showed
Event|Event|Hospital Course|9761,9769|true|false|false|||evidence
Finding|Idea or Concept|Hospital Course|9761,9769|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Hospital Course|9761,9772|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Finding|Functional Concept|Hospital Course|9773,9778|true|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|Hospital Course|9773,9784|true|false|false|C0225808|Right side of heart|right heart
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9779,9784|true|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Hospital Course|9779,9784|true|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Hospital Course|9779,9784|true|false|false|C0795691|HEART PROBLEM|heart
Disorder|Injury or Poisoning|Hospital Course|9785,9791|true|false|false|C0080194|Muscle strain|strain
Event|Event|Hospital Course|9785,9791|true|false|false|||strain
Finding|Idea or Concept|Hospital Course|9785,9791|true|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Finding|Mental Process|Hospital Course|9785,9791|true|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Finding|Physiologic Function|Hospital Course|9785,9791|true|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Finding|Sign or Symptom|Hospital Course|9785,9791|true|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Event|Event|Hospital Course|9802,9809|false|false|false|||treated
Drug|Biologically Active Substance|Hospital Course|9817,9824|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|Hospital Course|9817,9824|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|Hospital Course|9817,9824|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Event|Event|Hospital Course|9817,9824|false|false|false|||heparin
Disorder|Neoplastic Process|Hospital Course|9825,9828|false|false|false|C1135868|Gestational Trophoblastic Neoplasms|gtt
Drug|Biomedical or Dental Material|Hospital Course|9825,9828|false|false|false|C0991568|Drops - Drug Form|gtt
Event|Event|Hospital Course|9825,9828|false|false|false|||gtt
Procedure|Laboratory Procedure|Hospital Course|9825,9828|false|false|false|C0017741|Glucose tolerance test|gtt
Finding|Intellectual Product|Hospital Course|9830,9834|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|Hospital Course|9835,9847|false|false|false|||transitioned
Event|Event|Hospital Course|9851,9860|false|false|false|||treatment
Finding|Conceptual Entity|Hospital Course|9851,9860|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Hospital Course|9851,9860|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Hospital Course|9851,9860|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9851,9860|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Event|Event|Hospital Course|9861,9865|false|false|false|||dose
Drug|Organic Chemical|Hospital Course|9867,9874|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|Hospital Course|9867,9874|false|false|false|C0728963|Lovenox|lovenox
Disorder|Neoplastic Process|Hospital Course|9881,9891|false|false|false|C0006826;C1306459|Malignant Neoplasms;Primary malignant neoplasm|malignancy
Event|Event|Hospital Course|9881,9891|false|false|false|||malignancy
Event|Event|Hospital Course|9903,9913|false|false|false|||thrombosis
Finding|Pathologic Function|Hospital Course|9903,9913|false|false|false|C0040053|Thrombosis|thrombosis
Event|Event|Hospital Course|9917,9922|false|false|false|||noted
Drug|Organic Chemical|Hospital Course|9926,9930|false|false|false|C0009074|clotrimazole|CLOT
Drug|Pharmacologic Substance|Hospital Course|9926,9930|false|false|false|C0009074|clotrimazole|CLOT
Event|Event|Hospital Course|9926,9930|false|false|false|||CLOT
Finding|Pathologic Function|Hospital Course|9926,9930|false|false|false|C0302148|Blood Clot|CLOT
Event|Event|Hospital Course|9932,9937|false|false|false|||trial
Procedure|Research Activity|Hospital Course|9932,9937|false|false|false|C0008976|Clinical Trials|trial
Event|Event|Hospital Course|9952,9963|false|false|false|||symptomatic
Finding|Functional Concept|Hospital Course|9952,9963|false|false|false|C0231220|Symptomatic|symptomatic
Drug|Biologically Active Substance|Hospital Course|9977,9983|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|Hospital Course|9977,9983|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|Hospital Course|9977,9983|false|false|false|C0030054|oxygen|oxygen
Event|Event|Hospital Course|9977,9983|false|false|false|||oxygen
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9977,9983|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Event|Event|Hospital Course|9985,10000|false|false|false|||supplementation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9985,10000|false|false|false|C0242297|Dietary Supplementation|supplementation
Event|Event|Hospital Course|10009,10017|false|false|false|||improved
Event|Event|Hospital Course|10025,10040|false|false|false|||hospitalization
Procedure|Health Care Activity|Hospital Course|10025,10040|false|false|false|C0019993|Hospitalization|hospitalization
Drug|Biologically Active Substance|Hospital Course|10055,10061|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|Hospital Course|10055,10061|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|Hospital Course|10055,10061|false|false|false|C0030054|oxygen|oxygen
Event|Event|Hospital Course|10055,10061|false|false|false|||oxygen
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10055,10061|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Event|Event|Hospital Course|10065,10074|false|false|false|||tolerated
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10079,10088|false|false|false|C0024109|Lung|Pulmonary
Attribute|Clinical Attribute|Hospital Course|10079,10088|false|false|false|C2707265||Pulmonary
Finding|Finding|Hospital Course|10079,10088|false|false|false|C4522268|Pulmonary (intended site)|Pulmonary
Finding|Finding|Hospital Course|10079,10096|false|false|false|C0748164|Multiple Pulmonary Nodules|Pulmonary nodules
Event|Event|Hospital Course|10089,10096|false|false|false|||nodules
Event|Event|Hospital Course|10115,10121|false|false|false|||masses
Event|Event|Hospital Course|10132,10137|false|false|false|||noted
Event|Event|Hospital Course|10142,10144|false|false|false|||CT
Anatomy|Body Location or Region|Hospital Course|10176,10180|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10176,10180|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Hospital Course|10176,10180|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Hospital Course|10176,10180|false|false|false|C0740941|Lung Problem|lung
Disorder|Neoplastic Process|Hospital Course|10176,10191|false|true|false|C0242379|Malignant neoplasm of lung|lung malignancy
Disorder|Neoplastic Process|Hospital Course|10181,10191|false|true|false|C0006826;C1306459|Malignant Neoplasms;Primary malignant neoplasm|malignancy
Event|Event|Hospital Course|10181,10191|false|false|false|||malignancy
Event|Event|Hospital Course|10195,10199|false|false|false|||mets
Finding|Gene or Genome|Hospital Course|10195,10199|false|false|false|C0812270;C1705694|ETV3 gene;ETV3 wt Allele|mets
Phenomenon|Natural Phenomenon or Process|Hospital Course|10202,10209|false|false|false|C1705970|Electrical Current|Current
Event|Event|Hospital Course|10210,10212|false|false|false|||CT
Event|Event|Hospital Course|10213,10219|false|false|false|||showed
Finding|Intellectual Product|Hospital Course|10220,10226|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|Hospital Course|10227,10234|false|false|false|||nodules
Disorder|Disease or Syndrome|Hospital Course|10235,10240|false|false|false|C1410088|Still|still
Disorder|Neoplastic Process|Hospital Course|10257,10267|false|false|false|C0006826;C1306459|Malignant Neoplasms;Primary malignant neoplasm|malignancy
Event|Event|Hospital Course|10257,10267|false|false|false|||malignancy
Event|Event|Hospital Course|10277,10286|false|false|false|||evaluated
Anatomy|Body Location or Region|Hospital Course|10294,10302|false|false|false|C0817096|Chest|thoracic
Disorder|Disease or Syndrome|Hospital Course|10294,10302|false|false|false|C5779551|Dissecting Thoracic Aortic Aneurysm|thoracic
Event|Event|Hospital Course|10313,10324|false|false|false|||recommended
Event|Event|Hospital Course|10328,10334|false|false|false|||biopsy
Finding|Finding|Hospital Course|10328,10334|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Finding|Intellectual Product|Hospital Course|10328,10334|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Procedure|Diagnostic Procedure|Hospital Course|10328,10334|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Procedure|Health Care Activity|Hospital Course|10328,10334|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Event|Event|Hospital Course|10339,10351|false|false|false|||surveillance
Event|Occupational Activity|Hospital Course|10339,10351|false|false|false|C0684245|legal surveillance|surveillance
Finding|Functional Concept|Hospital Course|10339,10351|false|false|false|C0220920|surveillance aspects|surveillance
Procedure|Health Care Activity|Hospital Course|10339,10351|false|false|false|C0733511|Medical Surveillance|surveillance
Phenomenon|Natural Phenomenon or Process|Hospital Course|10363,10370|false|false|false|C1705970|Electrical Current|current
Anatomy|Body Location or Region|Hospital Course|10375,10378|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Hospital Course|10375,10378|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Hospital Course|10375,10378|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Finding|Classification|Hospital Course|10384,10390|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Hospital Course|10384,10390|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Hospital Course|10384,10390|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Hospital Course|10384,10390|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Body Substance|Hospital Course|10399,10406|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|10399,10406|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|10399,10406|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|10407,10414|false|false|false|||decided
Event|Event|Hospital Course|10419,10431|false|false|false|||surveillance
Event|Occupational Activity|Hospital Course|10419,10431|false|false|false|C0684245|legal surveillance|surveillance
Finding|Functional Concept|Hospital Course|10419,10431|false|false|false|C0220920|surveillance aspects|surveillance
Procedure|Health Care Activity|Hospital Course|10419,10431|false|false|false|C0733511|Medical Surveillance|surveillance
Finding|Finding|Hospital Course|10441,10445|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Hospital Course|10441,10445|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Hospital Course|10441,10445|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|Hospital Course|10457,10463|false|false|false|||follow
Finding|Intellectual Product|Hospital Course|10476,10488|false|false|false|C1547426|Location Service Code - Primary Care|primary care
Procedure|Health Care Activity|Hospital Course|10476,10488|false|false|false|C0033137|Primary Health Care|primary care
Attribute|Clinical Attribute|Hospital Course|10476,10497|false|false|false|C2735025||primary care provider
Finding|Idea or Concept|Hospital Course|10476,10497|false|false|false|C1547431|Primary Care Provider - Provider role|primary care provider
Event|Activity|Hospital Course|10484,10488|false|false|false|C1947933|care activity|care
Event|Event|Hospital Course|10484,10488|false|false|false|||care
Finding|Finding|Hospital Course|10484,10488|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Hospital Course|10484,10488|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Functional Concept|Hospital Course|10489,10497|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|provider
Finding|Intellectual Product|Hospital Course|10489,10497|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|provider
Disorder|Disease or Syndrome|Hospital Course|10516,10519|false|false|false|C0042029|Urinary tract infection|UTI
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10516,10519|false|false|false|C0077906|urinastatin|UTI
Drug|Pharmacologic Substance|Hospital Course|10516,10519|false|false|false|C0077906|urinastatin|UTI
Event|Event|Hospital Course|10516,10519|false|false|false|||UTI
Finding|Gene or Genome|Hospital Course|10516,10519|false|false|false|C1412376;C5780748|AMBP gene;AMBP wt Allele|UTI
Event|Event|Hospital Course|10528,10533|false|false|false|||noted
Anatomy|Cell|Hospital Course|10549,10552|false|false|false|C0023516|Leukocytes|WBC
Event|Event|Hospital Course|10549,10552|false|false|false|||WBC
Finding|Mental Process|Hospital Course|10560,10567|false|false|false|C0542559|contextual factors|setting
Anatomy|Anatomical Structure|Hospital Course|10581,10589|false|false|false|C0559495|Urological stoma|urostomy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10581,10589|false|false|false|C0856443|Urostomy procedure|urostomy
Event|Event|Hospital Course|10590,10597|false|false|false|||growing
Disorder|Disease or Syndrome|Hospital Course|10629,10641|false|false|false|C0023518|Leukocytosis|leukocytosis
Event|Event|Hospital Course|10629,10641|false|false|false|||leukocytosis
Finding|Finding|Hospital Course|10629,10641|false|false|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Event|Event|Hospital Course|10647,10656|false|false|false|||proceeded
Event|Event|Hospital Course|10662,10671|false|false|false|||treatment
Finding|Conceptual Entity|Hospital Course|10662,10671|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Hospital Course|10662,10671|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Hospital Course|10662,10671|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10662,10671|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Event|Event|Hospital Course|10681,10688|false|false|false|||started
Finding|Finding|Hospital Course|10689,10694|false|false|false|C3714655|On IV|on IV
Drug|Antibiotic|Hospital Course|10695,10705|false|false|false|C0002680;C2095775|ampicillin;ampicillins|Ampicillin
Drug|Organic Chemical|Hospital Course|10695,10705|false|false|false|C0002680;C2095775|ampicillin;ampicillins|Ampicillin
Event|Event|Hospital Course|10695,10705|false|false|false|||Ampicillin
Event|Event|Hospital Course|10711,10723|false|false|false|||transitioned
Drug|Organic Chemical|Hospital Course|10727,10735|false|false|false|C0591750|Macrobid|macrobid
Drug|Pharmacologic Substance|Hospital Course|10727,10735|false|false|false|C0591750|Macrobid|macrobid
Event|Event|Hospital Course|10746,10757|false|false|false|||sensitivies
Disorder|Disease or Syndrome|Hospital Course|10759,10771|false|false|false|C0023518|Leukocytosis|Leukocytosis
Event|Event|Hospital Course|10759,10771|false|false|false|||Leukocytosis
Finding|Finding|Hospital Course|10759,10771|false|false|false|C0750426|Blood leukocyte number above reference range|Leukocytosis
Event|Event|Hospital Course|10773,10781|false|false|false|||improved
Drug|Antibiotic|Hospital Course|10785,10796|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|Hospital Course|10785,10796|false|false|false|||antibiotics
Event|Event|Hospital Course|10809,10817|false|false|false|||complete
Finding|Idea or Concept|Hospital Course|10822,10825|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|10822,10825|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|10826,10832|false|false|false|||course
Finding|Idea or Concept|Hospital Course|10834,10837|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|10834,10837|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Idea or Concept|Hospital Course|10847,10850|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|10847,10850|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Finding|Hospital Course|10847,10852|false|false|false|C3842672|Day 7|day 7
Disorder|Disease or Syndrome|Hospital Course|10874,10880|false|false|false|C0002871|Anemia|Anemia
Event|Event|Hospital Course|10874,10880|false|false|false|||Anemia
Event|Event|Hospital Course|10885,10890|true|false|false|||signs
Finding|Finding|Hospital Course|10885,10890|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Hospital Course|10885,10890|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Event|Event|Hospital Course|10894,10902|true|false|false|||bleeding
Finding|Pathologic Function|Hospital Course|10894,10902|true|false|false|C0019080|Hemorrhage|bleeding
Event|Event|Hospital Course|10907,10916|true|false|false|||hemolysis
Finding|Cell Function|Hospital Course|10907,10916|true|false|false|C0019054;C1553188;C2937287;C2945560|Hemolysis (biological function);Hemolysis (disorder);Hemolysis (finding)|hemolysis
Finding|Finding|Hospital Course|10907,10916|true|false|false|C0019054;C1553188;C2937287;C2945560|Hemolysis (biological function);Hemolysis (disorder);Hemolysis (finding)|hemolysis
Finding|Pathologic Function|Hospital Course|10907,10916|true|false|false|C0019054;C1553188;C2937287;C2945560|Hemolysis (biological function);Hemolysis (disorder);Hemolysis (finding)|hemolysis
Event|Event|Hospital Course|10922,10929|false|false|false|||dropped
Event|Event|Hospital Course|10933,10938|false|false|false|||nadir
Event|Event|Hospital Course|10947,10953|false|false|false|||stable
Finding|Intellectual Product|Hospital Course|10947,10953|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|Hospital Course|10957,10966|false|false|false|||discharge
Finding|Body Substance|Hospital Course|10957,10966|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|10957,10966|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|10957,10966|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|10957,10966|false|false|false|C0030685|Patient Discharge|discharge
Drug|Biologically Active Substance|Hospital Course|10975,10979|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Element, Ion, or Isotope|Hospital Course|10975,10979|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Pharmacologic Substance|Hospital Course|10975,10979|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Event|Event|Hospital Course|10975,10979|false|false|false|||Iron
Procedure|Laboratory Procedure|Hospital Course|10975,10979|false|false|false|C0337439|Iron measurement|Iron
Event|Event|Hospital Course|10981,10988|false|false|false|||studies
Procedure|Research Activity|Hospital Course|10981,10988|false|false|false|C0947630|Scientific Study|studies
Event|Event|Hospital Course|10989,10999|false|false|false|||consistent
Finding|Idea or Concept|Hospital Course|10989,10999|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|Hospital Course|10989,11004|false|false|false|C0332290|Consistent with|consistent with
Finding|Finding|Hospital Course|11005,11011|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|11005,11011|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Finding|Hospital Course|11012,11023|false|true|false|C3811910|combination - answer to question|combination
Drug|Biologically Active Substance|Hospital Course|11024,11028|false|true|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|Hospital Course|11024,11028|false|true|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|Hospital Course|11024,11028|false|true|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Procedure|Laboratory Procedure|Hospital Course|11024,11028|false|true|false|C0337439|Iron measurement|iron
Disorder|Disease or Syndrome|Hospital Course|11024,11039|false|true|false|C0162316;C0240066|Iron deficiency;Iron deficiency anemia|iron deficiency
Disorder|Disease or Syndrome|Hospital Course|11029,11039|false|true|false|C0162429|Malnutrition|deficiency
Event|Event|Hospital Course|11029,11039|false|false|false|||deficiency
Finding|Functional Concept|Hospital Course|11029,11039|false|true|false|C0011155|Deficiency|deficiency
Disorder|Disease or Syndrome|Hospital Course|11041,11047|false|false|false|C0002871|Anemia|anemia
Event|Event|Hospital Course|11041,11047|false|false|false|||anemia
Disorder|Disease or Syndrome|Hospital Course|11052,11058|false|false|false|C0002871|Anemia|anemia
Event|Event|Hospital Course|11052,11058|false|false|false|||anemia
Disorder|Disease or Syndrome|Hospital Course|11052,11077|false|false|false|C0002873|Anemia of chronic disease|anemia of chronic disease
Finding|Intellectual Product|Hospital Course|11062,11069|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Hospital Course|11062,11069|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|Hospital Course|11062,11077|false|false|false|C0008679|Chronic disease|chronic disease
Disorder|Disease or Syndrome|Hospital Course|11070,11077|false|false|false|C0012634|Disease|disease
Event|Event|Hospital Course|11070,11077|false|false|false|||disease
Finding|Finding|Hospital Course|11083,11086|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Hospital Course|11083,11086|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Finding|Hospital Course|11083,11091|false|false|false|C0860975|Iron low|low iron
Drug|Biologically Active Substance|Hospital Course|11087,11091|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|Hospital Course|11087,11091|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|Hospital Course|11087,11091|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Event|Event|Hospital Course|11087,11091|false|false|false|||iron
Procedure|Laboratory Procedure|Hospital Course|11087,11091|false|false|false|C0337439|Iron measurement|iron
Event|Event|Hospital Course|11096,11104|false|false|false|||elevated
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11106,11114|false|false|false|C0015879|Ferritin|ferritin
Drug|Biologically Active Substance|Hospital Course|11106,11114|false|false|false|C0015879|Ferritin|ferritin
Drug|Pharmacologic Substance|Hospital Course|11106,11114|false|false|false|C0015879|Ferritin|ferritin
Event|Event|Hospital Course|11106,11114|false|false|false|||ferritin
Procedure|Laboratory Procedure|Hospital Course|11106,11114|false|false|false|C0373607|Ferritin measurement|ferritin
Finding|Finding|Hospital Course|11119,11122|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Hospital Course|11119,11122|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Event|Event|Hospital Course|11123,11127|false|false|false|||TIBC
Lab|Laboratory or Test Result|Hospital Course|11123,11127|false|false|false|C0036835|Total Iron-Binding Capacity result|TIBC
Procedure|Laboratory Procedure|Hospital Course|11123,11127|false|false|false|C1283048|Total iron binding capacity measurement|TIBC
Event|Event|Hospital Course|11135,11144|false|false|false|||recommend
Event|Event|Hospital Course|11145,11153|false|false|false|||checking
Event|Event|Hospital Course|11164,11174|false|false|false|||outpatient
Finding|Classification|Hospital Course|11164,11174|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|11164,11174|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|Hospital Course|11179,11183|false|false|false|||work
Event|Occupational Activity|Hospital Course|11179,11183|false|false|false|C0043227|Work|work
Procedure|Diagnostic Procedure|Hospital Course|11179,11186|false|false|false|C0750430|Work-up|work-up
Event|Event|Hospital Course|11190,11196|false|false|false|||needed
Event|Event|Hospital Course|11205,11213|false|false|false|||swelling
Finding|Finding|Hospital Course|11205,11213|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|Hospital Course|11205,11213|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Event|Event|Hospital Course|11222,11236|false|false|false|||multifactorial
Finding|Finding|Hospital Course|11222,11236|false|false|false|C1837655|Multifactorial|multifactorial
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11247,11253|false|false|false|C0042449|Veins|venous
Event|Event|Hospital Course|11255,11268|false|false|false|||insufficiency
Finding|Functional Concept|Hospital Course|11255,11268|false|false|false|C0231179|Insufficiency|insufficiency
Finding|Finding|Hospital Course|11273,11277|false|false|false|C5575035|Well (answer to question)|well
Anatomy|Body Location or Region|Hospital Course|11291,11294|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Hospital Course|11291,11294|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Hospital Course|11291,11294|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|Hospital Course|11291,11294|false|false|false|||DVT
Event|Event|Hospital Course|11300,11309|false|false|false|||responded
Event|Event|Hospital Course|11317,11321|false|false|false|||well
Finding|Finding|Hospital Course|11317,11321|false|false|false|C5575035|Well (answer to question)|well
Event|Event|Hospital Course|11327,11338|false|false|false|||compression
Finding|Functional Concept|Hospital Course|11327,11338|false|false|false|C0332459;C4551657|Compressed structure|compression
Phenomenon|Natural Phenomenon or Process|Hospital Course|11327,11338|false|false|false|C0728907|Compression|compression
Procedure|Machine Activity|Hospital Course|11327,11338|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11327,11338|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Event|Event|Hospital Course|11339,11348|false|false|false|||stockings
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11359,11366|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|Hospital Course|11359,11366|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11359,11366|false|false|false|C0872388|Procedures on bladder|bladder
Disorder|Neoplastic Process|Hospital Course|11359,11373|false|false|false|C0005684;C0005695;C0699885|Bladder Neoplasm;Carcinoma of bladder;Malignant neoplasm of urinary bladder|bladder cancer
Disorder|Neoplastic Process|Hospital Course|11367,11373|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Hospital Course|11367,11373|false|false|false|||cancer
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11383,11388|false|false|false|C0401496|Transurethral resection of neoplasm of bladder|TURBT
Finding|Finding|Hospital Course|11390,11394|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|Hospital Course|11390,11394|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|Hospital Course|11390,11394|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Classification|Hospital Course|11395,11400|true|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Finding|Finding|Hospital Course|11395,11400|true|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Anatomy|Cell Component|Hospital Course|11401,11404|true|false|false|C1167383|membrane attack complex location|TCC
Disorder|Disease or Syndrome|Hospital Course|11401,11404|true|false|false|C1861305|TARSAL-CARPAL COALITION SYNDROME|TCC
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11401,11404|true|false|false|C0077072;C5552697|Membrane Attack Complex;triclocarban|TCC
Drug|Biologically Active Substance|Hospital Course|11401,11404|true|false|false|C0077072;C5552697|Membrane Attack Complex;triclocarban|TCC
Drug|Organic Chemical|Hospital Course|11401,11404|true|false|false|C0077072;C5552697|Membrane Attack Complex;triclocarban|TCC
Drug|Pharmacologic Substance|Hospital Course|11401,11404|true|false|false|C0077072;C5552697|Membrane Attack Complex;triclocarban|TCC
Event|Event|Hospital Course|11401,11404|true|false|false|||TCC
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11414,11420|true|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|Hospital Course|11414,11420|true|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Event|Event|Hospital Course|11421,11431|true|false|false|||identified
Finding|Intellectual Product|Hospital Course|11434,11438|false|false|false|C1720594|Then - dosing instruction fragment|Then
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11447,11453|false|false|false|C0030797|Pelvis|pelvic
Procedure|Diagnostic Procedure|Hospital Course|11447,11457|false|false|false|C0203201|Magnetic Resonance Imaging (MRI) of Pelvis|pelvic MRI
Event|Event|Hospital Course|11454,11457|false|false|false|||MRI
Finding|Gene or Genome|Hospital Course|11454,11457|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|Hospital Course|11454,11457|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|Hospital Course|11454,11457|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Event|Event|Hospital Course|11458,11464|false|false|false|||showed
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11466,11473|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|Hospital Course|11466,11473|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11466,11473|false|false|false|C0872388|Procedures on bladder|bladder
Finding|Finding|Hospital Course|11466,11478|false|false|false|C0238775|Mass of urinary bladder|bladder mass
Finding|Finding|Hospital Course|11474,11478|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|Hospital Course|11474,11478|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Hospital Course|11474,11478|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Disorder|Neoplastic Process|Hospital Course|11479,11487|false|false|false|C1269955|Tumor Cell Invasion|invasion
Event|Event|Hospital Course|11479,11487|false|false|false|||invasion
Finding|Pathologic Function|Hospital Course|11479,11487|false|false|false|C2699153|Cell Invasion|invasion
Disorder|Disease or Syndrome|Hospital Course|11501,11505|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Anatomy|Body Location or Region|Hospital Course|11501,11512|false|false|false|C0225317;C4532079|Neck+Chest>Soft tissue;soft tissue|soft tissue
Anatomy|Tissue|Hospital Course|11501,11512|false|false|false|C0225317;C4532079|Neck+Chest>Soft tissue;soft tissue|soft tissue
Anatomy|Tissue|Hospital Course|11506,11512|false|false|false|C0040300|Body tissue|tissue
Finding|Intellectual Product|Hospital Course|11506,11512|false|false|false|C1547928|Tissue Specimen Code|tissue
Disorder|Disease or Syndrome|Hospital Course|11514,11522|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11523,11530|false|false|false|C0042232|Vagina|vaginal
Drug|Biomedical or Dental Material|Hospital Course|11523,11530|false|false|false|C1272941|Vaginal Dosage Form|vaginal
Finding|Finding|Hospital Course|11523,11530|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Finding|Functional Concept|Hospital Course|11523,11530|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Event|Event|Hospital Course|11540,11545|false|false|false|||right
Finding|Functional Concept|Hospital Course|11540,11545|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Event|Event|Hospital Course|11554,11560|false|false|false|||lesion
Finding|Finding|Hospital Course|11554,11560|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|Hospital Course|11554,11560|false|false|false|C0221198;C1546698|Lesion|lesion
Event|Event|Hospital Course|11581,11588|false|false|false|||robotic
Event|Event|Hospital Course|11590,11593|false|false|false|||TAH
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11590,11593|false|false|false|C0404079|Total abdominal hysterectomy|TAH
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11594,11597|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Drug|Hazardous or Poisonous Substance|Hospital Course|11594,11597|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Drug|Pharmacologic Substance|Hospital Course|11594,11597|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Event|Event|Hospital Course|11594,11597|false|false|false|||BSO
Disorder|Disease or Syndrome|Hospital Course|11599,11602|false|false|false|C0396060|Congenital laryngeal adductor palsy|lap
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11599,11602|false|false|false|C1870042|ACP2 protein, human|lap
Drug|Enzyme|Hospital Course|11599,11602|false|false|false|C1870042|ACP2 protein, human|lap
Event|Event|Hospital Course|11599,11602|false|false|false|||lap
Finding|Finding|Hospital Course|11599,11602|false|false|false|C0456170;C1412132;C1413323;C1423544;C1424863;C1425522;C2827449;C3540509;C5575443;C5890955|ACP2 gene;ACP2 wt Allele;CEBPB gene;CEBPB wt Allele;CENPJ gene;LAP3 gene;LAP3 wt Allele;Left atrial pressure;PICALM gene;PICALM wt Allele|lap
Finding|Gene or Genome|Hospital Course|11599,11602|false|false|false|C0456170;C1412132;C1413323;C1423544;C1424863;C1425522;C2827449;C3540509;C5575443;C5890955|ACP2 gene;ACP2 wt Allele;CEBPB gene;CEBPB wt Allele;CENPJ gene;LAP3 gene;LAP3 wt Allele;Left atrial pressure;PICALM gene;PICALM wt Allele|lap
Procedure|Diagnostic Procedure|Hospital Course|11599,11602|false|false|false|C0031150|Laparoscopy|lap
Drug|Chemical Viewed Structurally|Hospital Course|11603,11610|false|false|false|C0302912|Radicals (chemistry)|radical
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11603,11621|false|false|false|C0194401|Complete cystectomy|radical cystectomy
Event|Event|Hospital Course|11611,11621|false|false|false|||cystectomy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11611,11621|false|false|false|C0010651|Cystectomy|cystectomy
Disorder|Disease or Syndrome|Hospital Course|11626,11634|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Event|Event|Hospital Course|11635,11646|false|false|false|||vaginectomy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11635,11646|false|false|false|C0195130|Vaginectomy|vaginectomy
Event|Event|Hospital Course|11653,11662|false|false|false|||pathology
Finding|Functional Concept|Hospital Course|11653,11662|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Finding|Pathologic Function|Hospital Course|11653,11662|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Procedure|Laboratory Procedure|Hospital Course|11653,11662|false|false|false|C0919386|Pathology procedure|pathology
Event|Event|Hospital Course|11663,11670|false|false|false|||showing
Finding|Finding|Hospital Course|11671,11675|false|false|false|C1711132|pT2b TNM Finding|pT2b
Event|Event|Hospital Course|11686,11693|false|false|false|||margins
Event|Event|Hospital Course|11694,11702|false|false|false|||negative
Finding|Classification|Hospital Course|11694,11702|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|11694,11702|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|11694,11702|false|false|false|C5237010|Expression Negative|negative
Disorder|Disease or Syndrome|Hospital Course|11707,11711|true|false|false|C0270724|Infantile Neuroaxonal Dystrophy|plan
Event|Event|Hospital Course|11707,11711|true|false|false|||plan
Finding|Functional Concept|Hospital Course|11707,11711|true|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Intellectual Product|Hospital Course|11707,11711|true|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Mental Process|Hospital Course|11707,11711|true|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Event|Event|Hospital Course|11729,11736|true|false|false|||therapy
Finding|Finding|Hospital Course|11729,11736|true|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|Hospital Course|11729,11736|true|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11729,11736|true|false|false|C0087111|Therapeutic procedure|therapy
Finding|Finding|Hospital Course|11745,11749|true|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Hospital Course|11745,11749|true|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Hospital Course|11745,11749|true|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Body Substance|Hospital Course|11767,11774|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|11767,11774|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|11767,11774|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|11778,11782|false|false|false|||safe
Finding|Intellectual Product|Hospital Course|11778,11782|false|false|false|C4684764|SAFE-Biopharma Standard|safe
Event|Event|Hospital Course|11786,11795|false|false|false|||discharge
Finding|Body Substance|Hospital Course|11786,11795|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|11786,11795|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|11786,11795|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|11786,11795|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|Hospital Course|11819,11824|false|false|false|||spent
Event|Event|Hospital Course|11829,11838|false|false|false|||discharge
Finding|Body Substance|Hospital Course|11829,11838|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|11829,11838|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|11829,11838|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|11829,11838|false|false|false|C0030685|Patient Discharge|discharge
Finding|Idea or Concept|Hospital Course|11839,11842|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|11839,11842|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Occupational Activity|Hospital Course|11843,11853|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|Hospital Course|11843,11853|false|false|false|C0376636|Disease Management|management
Event|Event|Hospital Course|11854,11862|false|false|false|||services
Event|Occupational Activity|Hospital Course|11854,11862|false|false|false|C0557854|Services|services
Procedure|Health Care Activity|Hospital Course|11854,11862|false|false|false|C1704289|Clinical Service|services
Finding|Idea or Concept|Hospital Course|11865,11877|false|false|false|C1548597|Marketing basis - Transitional|Transitional
Event|Event|Hospital Course|11878,11884|false|false|false|||issues
Event|Event|Hospital Course|11897,11901|false|false|false|||need
Event|Event|Hospital Course|11902,11908|false|false|false|||follow
Anatomy|Body Location or Region|Hospital Course|11912,11917|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|11912,11917|false|false|false|C0741025|Chest problem|chest
Procedure|Diagnostic Procedure|Hospital Course|11912,11920|false|false|false|C0202823|Chest CT|chest CT
Event|Event|Hospital Course|11918,11920|false|false|false|||CT
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11925,11934|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Hospital Course|11925,11934|false|false|false|C2707265||pulmonary
Finding|Finding|Hospital Course|11925,11934|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Finding|Hospital Course|11925,11942|false|false|false|C0748164|Multiple Pulmonary Nodules|pulmonary nodules
Event|Event|Hospital Course|11935,11942|false|false|false|||nodules
Drug|Organic Chemical|Hospital Course|11967,11975|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Hospital Course|11967,11975|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Hospital Course|11967,11975|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Finding|Functional Concept|Hospital Course|11967,11975|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|11967,11975|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|11978,11981|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|11978,11981|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|11982,11988|false|false|false|||course
Disorder|Disease or Syndrome|Hospital Course|11993,11996|false|false|false|C0042029|Urinary tract infection|UTI
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11993,11996|false|false|false|C0077906|urinastatin|UTI
Drug|Pharmacologic Substance|Hospital Course|11993,11996|false|false|false|C0077906|urinastatin|UTI
Event|Event|Hospital Course|11993,11996|false|false|false|||UTI
Finding|Gene or Genome|Hospital Course|11993,11996|false|false|false|C1412376;C5780748|AMBP gene;AMBP wt Allele|UTI
Drug|Organic Chemical|Hospital Course|12002,12010|false|false|false|C0591750|Macrobid|macrobid
Drug|Pharmacologic Substance|Hospital Course|12002,12010|false|false|false|C0591750|Macrobid|macrobid
Event|Event|Hospital Course|12002,12010|false|false|false|||macrobid
Event|Event|Hospital Course|12012,12015|false|false|false|||day
Finding|Idea or Concept|Hospital Course|12012,12015|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|12012,12015|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Finding|Hospital Course|12012,12017|false|false|false|C3842672|Day 7|day 7
Drug|Biologically Active Substance|Hospital Course|12034,12040|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|Hospital Course|12034,12040|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|Hospital Course|12034,12040|false|false|false|C0030054|oxygen|oxygen
Procedure|Therapeutic or Preventive Procedure|Hospital Course|12034,12040|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Finding|Finding|Hospital Course|12034,12048|false|false|false|C1546419|Ambulatory Status - Oxygen therapy|oxygen therapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|12034,12048|false|false|false|C0184633;C3665674|Oxygen Therapy Care;Warburg Therapy|oxygen therapy
Event|Event|Hospital Course|12041,12048|false|false|false|||therapy
Finding|Finding|Hospital Course|12041,12048|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|Hospital Course|12041,12048|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|12041,12048|false|false|false|C0087111|Therapeutic procedure|therapy
Finding|Finding|Hospital Course|12053,12057|false|false|false|C0043084|Weaning|wean
Event|Event|Hospital Course|12061,12070|false|false|false|||tolerated
Drug|Substance|Hospital Course|12074,12082|false|false|false|C0721534|Maintain brand of benzocaine|maintain
Event|Activity|Hospital Course|12074,12082|false|false|false|C0024501|Maintenance|maintain
Event|Event|Hospital Course|12087,12090|false|false|false|||sat
Event|Event|Hospital Course|12107,12112|false|false|false|||check
Anatomy|Cell Component|Hospital Course|12113,12116|false|false|false|C2263086|Nuclear cap binding complex location|CBC
Event|Event|Hospital Course|12113,12116|false|false|false|||CBC
Procedure|Laboratory Procedure|Hospital Course|12113,12116|false|false|false|C0009555|Complete Blood Count|CBC
Event|Event|Hospital Course|12127,12133|false|false|false|||ensure
Event|Event|Hospital Course|12134,12143|false|false|false|||stability
Event|Event|Hospital Course|12156,12167|false|false|false|||demonstrate
Event|Event|Hospital Course|12168,12178|false|false|false|||resolution
Finding|Conceptual Entity|Hospital Course|12168,12178|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolution
Finding|Pathologic Function|Hospital Course|12168,12178|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolution
Disorder|Disease or Syndrome|Hospital Course|12182,12194|false|false|false|C0023518|Leukocytosis|leukocytosis
Event|Event|Hospital Course|12182,12194|false|false|false|||leukocytosis
Finding|Finding|Hospital Course|12182,12194|false|false|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Disorder|Disease or Syndrome|Hospital Course|12197,12200|false|false|false|C0162531|Hereditary Coproporphyria|HCP
Event|Event|Hospital Course|12197,12200|false|false|false|||HCP
Finding|Gene or Genome|Hospital Course|12197,12200|false|false|false|C1335283;C1412376;C1413681;C1705637;C5780748|AMBP gene;AMBP wt Allele;CPOX gene;PTPN6 gene;PTPN6 wt Allele|HCP
Finding|Gene or Genome|Hospital Course|12202,12205|false|false|false|C1420310|SON gene|son
Attribute|Clinical Attribute|Hospital Course|12222,12233|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|12222,12233|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|12222,12233|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|12222,12233|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|12222,12246|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|12237,12246|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|12237,12246|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|Hospital Course|12265,12275|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Hospital Course|12265,12275|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|Hospital Course|12265,12280|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|Hospital Course|12276,12280|false|false|false|||list
Finding|Intellectual Product|Hospital Course|12276,12280|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|Hospital Course|12288,12298|false|false|false|||inaccurate
Event|Event|Hospital Course|12303,12311|false|false|false|||requires
Event|Event|Hospital Course|12320,12333|false|false|false|||investigation
Finding|Intellectual Product|Hospital Course|12320,12333|false|false|false|C1552578|Act Class - investigation|investigation
Procedure|Health Care Activity|Hospital Course|12320,12333|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|investigation
Drug|Organic Chemical|Hospital Course|12338,12351|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|12338,12351|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Hospital Course|12338,12351|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|12338,12351|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Organic Chemical|Hospital Course|12370,12378|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|12370,12378|false|false|false|C1692318|docusate|Docusate
Event|Event|Hospital Course|12370,12378|false|false|false|||Docusate
Drug|Organic Chemical|Hospital Course|12370,12385|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|Hospital Course|12370,12385|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|Hospital Course|12379,12385|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|12379,12385|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|12379,12385|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|12379,12385|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|12379,12385|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|12379,12385|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|Hospital Course|12396,12399|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12396,12399|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|12396,12399|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|12396,12399|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|12396,12399|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|12404,12414|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Pharmacologic Substance|Hospital Course|12404,12414|false|false|false|C0206460|enoxaparin|Enoxaparin
Event|Event|Hospital Course|12404,12414|false|false|false|||Enoxaparin
Drug|Organic Chemical|Hospital Course|12404,12421|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Pharmacologic Substance|Hospital Course|12404,12421|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Biologically Active Substance|Hospital Course|12415,12421|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|12415,12421|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|12415,12421|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|12415,12421|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|12415,12421|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|12415,12421|false|false|false|C0337443|Sodium measurement|Sodium
Event|Event|Hospital Course|12438,12443|false|false|false|||Start
Finding|Idea or Concept|Hospital Course|12462,12466|false|false|false|C1552851|next - HtmlLinkType|Next
Event|Event|Hospital Course|12467,12474|false|false|false|||Routine
Finding|Idea or Concept|Hospital Course|12467,12474|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Finding|Intellectual Product|Hospital Course|12467,12474|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Procedure|Laboratory Procedure|Hospital Course|12467,12474|false|false|false|C1979801|Routine coag|Routine
Event|Occupational Activity|Hospital Course|12475,12489|false|false|false|C0001554|Administration occupational activities|Administration
Procedure|Therapeutic or Preventive Procedure|Hospital Course|12475,12489|false|false|false|C1533734|Administration (procedure)|Administration
Finding|Finding|Hospital Course|12490,12494|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Finding|Idea or Concept|Hospital Course|12490,12494|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Finding|Intellectual Product|Hospital Course|12490,12494|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12499,12512|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Hormone|Hospital Course|12499,12512|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Organic Chemical|Hospital Course|12499,12512|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Pharmacologic Substance|Hospital Course|12499,12512|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Event|Event|Hospital Course|12499,12512|false|false|false|||Levothyroxine
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12499,12519|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Hormone|Hospital Course|12499,12519|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Pharmacologic Substance|Hospital Course|12499,12519|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Biologically Active Substance|Hospital Course|12513,12519|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|12513,12519|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|12513,12519|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|12513,12519|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|12513,12519|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|12513,12519|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Organic Chemical|Hospital Course|12541,12553|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|12541,12553|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|Hospital Course|12571,12579|false|false|false|C0126174|losartan|Losartan
Drug|Pharmacologic Substance|Hospital Course|12571,12579|false|false|false|C0126174|losartan|Losartan
Event|Event|Hospital Course|12571,12579|false|false|false|||Losartan
Drug|Organic Chemical|Hospital Course|12571,12589|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Pharmacologic Substance|Hospital Course|12571,12589|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Biologically Active Substance|Hospital Course|12580,12589|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|Hospital Course|12580,12589|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|Hospital Course|12580,12589|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|Hospital Course|12580,12589|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|Hospital Course|12580,12589|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Event|Event|Hospital Course|12580,12589|false|false|false|||Potassium
Finding|Physiologic Function|Hospital Course|12580,12589|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|Hospital Course|12580,12589|false|false|false|C0202194|Potassium measurement|Potassium
Drug|Organic Chemical|Hospital Course|12609,12618|false|false|false|C0030049|oxycodone|OxyCODONE
Drug|Pharmacologic Substance|Hospital Course|12609,12618|false|false|false|C0030049|oxycodone|OxyCODONE
Event|Event|Hospital Course|12609,12618|false|false|false|||OxyCODONE
Procedure|Laboratory Procedure|Hospital Course|12609,12618|false|false|false|C0524222|Oxycodone measurement|OxyCODONE
Finding|Idea or Concept|Hospital Course|12620,12629|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Finding|Intellectual Product|Hospital Course|12620,12629|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Drug|Biomedical or Dental Material|Hospital Course|12620,12637|false|false|false|C1708470|Immediate Release Dosage Form|Immediate Release
Event|Event|Hospital Course|12630,12637|false|false|false|||Release
Finding|Functional Concept|Hospital Course|12630,12637|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|12630,12637|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|12630,12637|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Finding|Gene or Genome|Hospital Course|12651,12654|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|12655,12659|false|false|false|C2598155||Pain
Event|Event|Hospital Course|12655,12659|false|false|false|||Pain
Finding|Functional Concept|Hospital Course|12655,12659|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Hospital Course|12655,12659|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Finding|Hospital Course|12662,12670|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|Hospital Course|12662,12670|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Drug|Organic Chemical|Hospital Course|12676,12685|false|false|false|C0024002|lorazepam|LORazepam
Drug|Pharmacologic Substance|Hospital Course|12676,12685|false|false|false|C0024002|lorazepam|LORazepam
Disorder|Mental or Behavioral Dysfunction|Hospital Course|12697,12700|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12697,12700|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|12697,12700|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|12697,12700|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|12697,12700|false|false|false|C1332410|BID gene|BID
Finding|Gene or Genome|Hospital Course|12701,12704|false|false|false|C1422467|CIAO3 gene|PRN
Disorder|Mental or Behavioral Dysfunction|Hospital Course|12705,12712|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|Hospital Course|12705,12712|false|false|false|||anxiety
Finding|Sign or Symptom|Hospital Course|12705,12712|false|false|false|C0860603|Anxiety symptoms|anxiety
Drug|Organic Chemical|Hospital Course|12717,12722|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|Hospital Course|12717,12722|false|false|false|C3489575|sennosides, USP|Senna
Disorder|Mental or Behavioral Dysfunction|Hospital Course|12733,12736|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12733,12736|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|12733,12736|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|12733,12736|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|12733,12736|false|false|false|C1332410|BID gene|BID
Event|Event|Hospital Course|12741,12750|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|12741,12750|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|12741,12750|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|12741,12750|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|12741,12750|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|12741,12762|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|12751,12762|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|12751,12762|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|12751,12762|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|12751,12762|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|12768,12782|false|false|false|C0028156|nitrofurantoin|Nitrofurantoin
Drug|Pharmacologic Substance|Hospital Course|12768,12782|false|false|false|C0028156|nitrofurantoin|Nitrofurantoin
Drug|Organic Chemical|Hospital Course|12792,12800|false|false|false|C0591750|Macrobid|MacroBID
Drug|Pharmacologic Substance|Hospital Course|12792,12800|false|false|false|C0591750|Macrobid|MacroBID
Finding|Idea or Concept|Hospital Course|12823,12826|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|12823,12826|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|12834,12844|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Pharmacologic Substance|Hospital Course|12834,12844|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Organic Chemical|Hospital Course|12834,12851|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Pharmacologic Substance|Hospital Course|12834,12851|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Biologically Active Substance|Hospital Course|12845,12851|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|12845,12851|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|12845,12851|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|12845,12851|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|12845,12851|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|12845,12851|false|false|false|C0337443|Sodium measurement|Sodium
Event|Event|Hospital Course|12867,12872|false|false|false|||Start
Finding|Idea or Concept|Hospital Course|12899,12903|false|false|false|C1552851|next - HtmlLinkType|Next
Finding|Idea or Concept|Hospital Course|12904,12911|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Finding|Intellectual Product|Hospital Course|12904,12911|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Procedure|Laboratory Procedure|Hospital Course|12904,12911|false|false|false|C1979801|Routine coag|Routine
Event|Event|Hospital Course|12912,12926|false|false|false|||Administration
Event|Occupational Activity|Hospital Course|12912,12926|false|false|false|C0001554|Administration occupational activities|Administration
Procedure|Therapeutic or Preventive Procedure|Hospital Course|12912,12926|false|false|false|C1533734|Administration (procedure)|Administration
Finding|Finding|Hospital Course|12928,12932|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Finding|Idea or Concept|Hospital Course|12928,12932|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Finding|Intellectual Product|Hospital Course|12928,12932|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Drug|Organic Chemical|Hospital Course|12939,12948|false|false|false|C0024002|lorazepam|LORazepam
Drug|Pharmacologic Substance|Hospital Course|12939,12948|false|false|false|C0024002|lorazepam|LORazepam
Finding|Gene or Genome|Hospital Course|12964,12967|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Pharmacologic Substance|Hospital Course|12968,12976|false|false|false|C1950154|Insomnia homeopathic medication|insomnia
Event|Event|Hospital Course|12968,12976|false|false|false|||insomnia
Finding|Sign or Symptom|Hospital Course|12968,12976|false|false|false|C0917801|Sleeplessness|insomnia
Event|Event|Hospital Course|12978,12980|false|false|false|||RX
Drug|Organic Chemical|Hospital Course|12982,12991|false|false|false|C0024002|lorazepam|lorazepam
Drug|Pharmacologic Substance|Hospital Course|12982,12991|false|false|false|C0024002|lorazepam|lorazepam
Event|Event|Hospital Course|12982,12991|false|false|false|||lorazepam
Drug|Biomedical or Dental Material|Hospital Course|13014,13017|false|false|false|C0039225|Tablet Dosage Form|tab
Event|Event|Hospital Course|13014,13017|false|false|false|||tab
Finding|Functional Concept|Hospital Course|13018,13026|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|13021,13026|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|13021,13026|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Gene or Genome|Hospital Course|13031,13034|false|false|false|C1422467|CIAO3 gene|prn
Event|Activity|Hospital Course|13035,13039|false|false|false|C1880359|Dispense (activity)|Disp
Event|Event|Hospital Course|13035,13039|false|false|false|||Disp
Finding|Gene or Genome|Hospital Course|13035,13039|false|false|false|C2828567|PRSS30P gene|Disp
Drug|Biomedical or Dental Material|Hospital Course|13045,13051|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|13052,13059|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|13052,13059|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|13068,13081|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|13068,13081|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Hospital Course|13068,13081|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|13068,13081|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Organic Chemical|Hospital Course|13102,13114|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|13102,13114|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|Hospital Course|13134,13142|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|13134,13142|false|false|false|C1692318|docusate|Docusate
Event|Event|Hospital Course|13134,13142|false|false|false|||Docusate
Drug|Organic Chemical|Hospital Course|13134,13149|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|Hospital Course|13134,13149|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|Hospital Course|13143,13149|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|13143,13149|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|13143,13149|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|13143,13149|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|13143,13149|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|13143,13149|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|Hospital Course|13160,13163|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|13160,13163|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|13160,13163|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|13160,13163|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|13160,13163|false|false|false|C1332410|BID gene|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|13170,13183|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Hormone|Hospital Course|13170,13183|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Organic Chemical|Hospital Course|13170,13183|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Pharmacologic Substance|Hospital Course|13170,13183|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Amino Acid, Peptide, or Protein|Hospital Course|13170,13190|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Hormone|Hospital Course|13170,13190|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Pharmacologic Substance|Hospital Course|13170,13190|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Biologically Active Substance|Hospital Course|13184,13190|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|13184,13190|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|13184,13190|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|13184,13190|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|13184,13190|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|13184,13190|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Organic Chemical|Hospital Course|13214,13223|false|false|false|C0030049|oxycodone|OxyCODONE
Drug|Pharmacologic Substance|Hospital Course|13214,13223|false|false|false|C0030049|oxycodone|OxyCODONE
Event|Event|Hospital Course|13214,13223|false|false|false|||OxyCODONE
Procedure|Laboratory Procedure|Hospital Course|13214,13223|false|false|false|C0524222|Oxycodone measurement|OxyCODONE
Finding|Idea or Concept|Hospital Course|13225,13234|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Finding|Intellectual Product|Hospital Course|13225,13234|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Drug|Biomedical or Dental Material|Hospital Course|13225,13242|false|false|false|C1708470|Immediate Release Dosage Form|Immediate Release
Event|Event|Hospital Course|13235,13242|false|false|false|||Release
Finding|Functional Concept|Hospital Course|13235,13242|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|13235,13242|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|13235,13242|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Finding|Gene or Genome|Hospital Course|13256,13259|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|13260,13264|false|false|false|C2598155||Pain
Finding|Functional Concept|Hospital Course|13260,13264|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Hospital Course|13260,13264|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Finding|Hospital Course|13268,13276|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|Hospital Course|13268,13276|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Event|Event|Hospital Course|13278,13280|false|false|false|||RX
Drug|Organic Chemical|Hospital Course|13282,13291|false|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|Hospital Course|13282,13291|false|false|false|C0030049|oxycodone|oxycodone
Event|Event|Hospital Course|13282,13291|false|false|false|||oxycodone
Procedure|Laboratory Procedure|Hospital Course|13282,13291|false|false|false|C0524222|Oxycodone measurement|oxycodone
Drug|Biomedical or Dental Material|Hospital Course|13299,13305|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|13309,13317|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|13312,13317|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|13312,13317|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Gene or Genome|Hospital Course|13322,13325|false|false|false|C1422467|CIAO3 gene|prn
Drug|Biomedical or Dental Material|Hospital Course|13335,13341|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|13335,13341|false|false|false|||Tablet
Event|Event|Hospital Course|13343,13350|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|13343,13350|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|13359,13364|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|Hospital Course|13359,13364|false|false|false|C3489575|sennosides, USP|Senna
Disorder|Mental or Behavioral Dysfunction|Hospital Course|13375,13378|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|13375,13378|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|13375,13378|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|13375,13378|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|13375,13378|false|false|false|C1332410|BID gene|BID
Event|Event|Hospital Course|13384,13393|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|13384,13393|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|13384,13393|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|13384,13393|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|13384,13393|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|13384,13405|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|13384,13405|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|13394,13405|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|13394,13405|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|13394,13405|false|false|false|C0184758|Patient disposition|Disposition
Finding|Finding|Hospital Course|13407,13415|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|13407,13415|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Procedure|Health Care Activity|Hospital Course|13407,13420|false|false|false|C0023977|long-term care|Extended Care
Event|Activity|Hospital Course|13416,13420|false|false|false|C1947933|care activity|Care
Event|Event|Hospital Course|13416,13420|false|false|false|||Care
Finding|Finding|Hospital Course|13416,13420|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Hospital Course|13416,13420|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Event|Event|Hospital Course|13423,13431|false|false|false|||Facility
Finding|Intellectual Product|Hospital Course|13423,13431|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|Hospital Course|13439,13448|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|13439,13448|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|13439,13448|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|13439,13448|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|13439,13448|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|13439,13458|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|13449,13458|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|13449,13458|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|13449,13458|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|13449,13458|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|13449,13458|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Mental Process|Discharge Condition|13486,13492|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|13486,13499|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|13486,13499|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|13493,13499|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|13493,13499|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|13501,13506|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|13501,13506|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|13511,13519|false|false|false|||coherent
Finding|Finding|Discharge Condition|13511,13519|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|13521,13526|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|13521,13543|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|13521,13543|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|13530,13543|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|13530,13543|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|13530,13543|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|13545,13550|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|13545,13550|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|13545,13550|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|13545,13550|false|false|false|||Alert
Finding|Finding|Discharge Condition|13545,13550|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|13545,13550|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|13545,13550|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|13555,13566|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|13555,13566|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|13568,13576|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|13568,13576|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|13568,13576|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|13577,13583|false|false|false|C5889824||Status
Event|Event|Discharge Condition|13577,13583|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|13577,13583|false|false|false|C1546481|What subject filter - Status|Status
Disorder|Disease or Syndrome|Discharge Condition|13592,13595|false|false|false|C3159311|BORNHOLM EYE DISEASE|Bed
Event|Event|Discharge Condition|13592,13595|false|false|false|||Bed
Finding|Intellectual Product|Discharge Condition|13592,13595|false|false|false|C2346952|Bachelor of Education|Bed
Event|Event|Discharge Condition|13601,13611|false|false|false|||assistance
Finding|Social Behavior|Discharge Condition|13601,13611|false|false|false|C0018896|Helping Behavior|assistance
Event|Event|Discharge Condition|13625,13635|false|false|false|||wheelchair
Finding|Finding|Discharge Condition|13625,13635|false|false|false|C2135586;C4321408|Wheelchair Usually Used;has wheelchair at home (history)|wheelchair
Event|Event|Discharge Instructions|13681,13689|false|false|false|||pleasure
Finding|Intellectual Product|Discharge Instructions|13681,13689|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|Discharge Instructions|13681,13689|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|Discharge Instructions|13697,13701|false|false|false|C1947933|care activity|care
Event|Event|Discharge Instructions|13697,13701|false|false|false|||care
Finding|Finding|Discharge Instructions|13697,13701|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|13697,13701|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Event|Event|Discharge Instructions|13719,13728|false|false|false|||admission
Procedure|Health Care Activity|Discharge Instructions|13719,13728|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|Discharge Instructions|13746,13754|false|false|false|||admitted
Drug|Organic Chemical|Discharge Instructions|13761,13765|false|false|false|C0009074|clotrimazole|clot
Drug|Pharmacologic Substance|Discharge Instructions|13761,13765|false|false|false|C0009074|clotrimazole|clot
Event|Event|Discharge Instructions|13761,13765|false|false|false|||clot
Finding|Pathologic Function|Discharge Instructions|13761,13765|false|false|false|C0302148|Blood Clot|clot
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|13774,13779|false|false|false|C0024109|Lung|lungs
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|13785,13788|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Event|Event|Discharge Instructions|13799,13806|false|false|false|||treated
Disorder|Disease or Syndrome|Discharge Instructions|13814,13819|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Discharge Instructions|13814,13819|false|false|false|||blood
Finding|Body Substance|Discharge Instructions|13814,13819|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Event|Discharge Instructions|13820,13827|false|false|false|||thinner
Event|Event|Discharge Instructions|13838,13842|false|false|false|||need
Event|Event|Discharge Instructions|13847,13855|false|false|false|||continue
Disorder|Disease or Syndrome|Discharge Instructions|13860,13865|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Discharge Instructions|13860,13865|false|false|false|||blood
Finding|Body Substance|Discharge Instructions|13860,13865|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Event|Discharge Instructions|13866,13873|false|false|false|||thinner
Event|Event|Discharge Instructions|13889,13896|false|false|false|||treated
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|13903,13910|false|false|false|C0042027|Urinary tract|urinary
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|13912,13917|false|false|false|C1185740|Tract|tract
Disorder|Disease or Syndrome|Discharge Instructions|13918,13927|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|Discharge Instructions|13918,13927|false|false|false|||infection
Finding|Pathologic Function|Discharge Instructions|13918,13927|false|false|false|C3714514|Infection|infection
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|13938,13947|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Discharge Instructions|13938,13947|false|false|false|C2707265||pulmonary
Finding|Finding|Discharge Instructions|13938,13947|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Finding|Discharge Instructions|13938,13955|false|false|false|C0748164|Multiple Pulmonary Nodules|pulmonary nodules
Event|Event|Discharge Instructions|13948,13955|false|false|false|||nodules
Event|Event|Discharge Instructions|13968,13974|false|false|false|||follow
Finding|Intellectual Product|Discharge Instructions|13989,14001|false|false|false|C1547426|Location Service Code - Primary Care|primary care
Procedure|Health Care Activity|Discharge Instructions|13989,14001|false|false|false|C0033137|Primary Health Care|primary care
Event|Activity|Discharge Instructions|13997,14001|false|false|false|C1947933|care activity|care
Event|Event|Discharge Instructions|13997,14001|false|false|false|||care
Finding|Finding|Discharge Instructions|13997,14001|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|13997,14001|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|14002,14008|false|false|false|C2348314|Doctor - Title|doctor
Procedure|Health Care Activity|Discharge Instructions|14013,14021|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|14022,14034|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|14022,14034|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|14022,14034|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

