 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|22,26
No|27,29
:|29,30
_|33,34
_|34,35
_|35,36
<EOL>|36,37
<EOL>|38,39
Admission|39,48
Date|49,53
:|53,54
_|56,57
_|57,58
_|58,59
Discharge|73,82
Date|83,87
:|87,88
_|91,92
_|92,93
_|93,94
<EOL>|94,95
<EOL>|96,97
Date|97,101
of|102,104
Birth|105,110
:|110,111
_|113,114
_|114,115
_|115,116
Sex|129,132
:|132,133
F|136,137
<EOL>|137,138
<EOL>|139,140
Service|140,147
:|147,148
MEDICINE|149,157
<EOL>|157,158
<EOL>|159,160
No|172,174
Known|175,180
Allergies|181,190
/|191,192
Adverse|193,200
Drug|201,205
Reactions|206,215
<EOL>|215,216
<EOL>|217,218
Attending|218,227
:|227,228
_|229,230
_|230,231
_|231,232
.|232,233
<EOL>|233,234
<EOL>|235,236
dyspnea|253,260
on|261,263
exertion|264,272
<EOL>|272,273
<EOL>|274,275
Major|275,280
Surgical|281,289
or|290,292
Invasive|293,301
Procedure|302,311
:|311,312
<EOL>|312,313
None|313,317
<EOL>|317,318
<EOL>|318,319
<EOL>|320,321
_|349,350
_|350,351
_|351,352
with|353,357
a|358,359
history|360,367
of|368,370
of|371,373
HTN|374,377
,|377,378
CAD|379,382
s|383,384
/|384,385
p|385,386
DES|387,390
with|391,395
ischemic|396,404
MR|405,407
and|408,411
<EOL>|412,413
systolic|413,421
dysfunction|422,433
,|433,434
_|435,436
_|436,437
_|437,438
on|439,441
torsemide|442,451
,|451,452
hx|453,455
of|456,458
DVT|459,462
,|462,463
who|464,467
presents|468,476
<EOL>|477,478
with|478,482
4|483,484
days|485,489
of|490,492
dyspnea|493,500
on|501,503
exertion|504,512
,|512,513
leg|514,517
swelling|518,526
,|526,527
and|528,531
10|532,534
weight|535,541
<EOL>|542,543
gain|543,547
.|547,548
<EOL>|548,549
<EOL>|549,550
Of|550,552
note|553,557
,|557,558
patient|559,566
was|567,570
seen|571,575
in|576,578
the|579,582
Heart|583,588
Failure|589,596
Clinic|597,603
with|604,608
Dr|609,611
.|611,612
<EOL>|613,614
_|614,615
_|615,616
_|616,617
on|618,620
_|621,622
_|622,623
_|623,624
where|625,630
she|631,634
noted|635,640
that|641,645
she|646,649
has|650,653
had|654,657
<EOL>|658,659
persistent|659,669
dyspnea|670,677
on|678,680
exertion|681,689
and|690,693
PND|694,697
after|698,703
a|704,705
lengthy|706,713
prior|714,719
<EOL>|720,721
hospitalization|721,736
for|737,740
DVT|741,744
/|744,745
GIB|745,748
.|748,749
At|750,752
that|753,757
time|758,762
she|763,766
was|767,770
started|771,778
on|779,781
<EOL>|782,783
40mg|783,787
po|788,790
torsemide|791,800
which|801,806
initially|807,816
improved|817,825
her|826,829
symptoms|830,838
.|838,839
<EOL>|840,841
<EOL>|841,842
Over|842,846
the|847,850
holiday|851,858
she|859,862
indulged|863,871
in|872,874
a|875,876
high|877,881
salt|882,886
diet|887,891
and|892,895
developed|896,905
<EOL>|906,907
slow|907,911
-|911,912
onset|912,917
dyspnea|918,925
on|926,928
exertion|929,937
.|937,938
Denies|939,945
any|946,949
medication|950,960
<EOL>|961,962
noncompliance|962,975
,|975,976
chest|977,982
pain|983,987
,|987,988
palpitations|989,1001
,|1001,1002
palpitations|1003,1015
.|1015,1016
Describes|1017,1026
<EOL>|1027,1028
PND|1028,1031
,|1031,1032
worsening|1033,1042
exercise|1043,1051
tolerance|1052,1061
(|1062,1063
unable|1063,1069
to|1070,1072
walk|1073,1077
>|1078,1079
50|1079,1081
feet|1082,1086
)|1086,1087
and|1088,1091
<EOL>|1092,1093
orthopnea|1093,1102
.|1102,1103
<EOL>|1104,1105
<EOL>|1105,1106
In|1106,1108
the|1109,1112
ED|1113,1115
,|1115,1116
patient|1117,1124
was|1125,1128
found|1129,1134
to|1135,1137
have|1138,1142
1|1143,1144
+|1144,1145
bilateral|1146,1155
lower|1156,1161
<EOL>|1162,1163
extremity|1163,1172
edema|1173,1178
,|1178,1179
and|1180,1183
have|1184,1188
bibasilar|1189,1198
crackles|1199,1207
on|1208,1210
exam|1211,1215
.|1215,1216
Patient|1217,1224
<EOL>|1225,1226
underwent|1226,1235
CXR|1236,1239
,|1239,1240
BNP|1241,1244
,|1244,1245
and|1246,1249
was|1250,1253
given|1254,1259
one|1260,1263
dose|1264,1268
of|1269,1271
IV|1272,1274
40mg|1275,1279
Lasix|1280,1285
.|1285,1286
In|1287,1289
<EOL>|1290,1291
the|1291,1294
ED|1295,1297
initial|1298,1305
vitals|1306,1312
were|1313,1317
:|1317,1318
97.8|1319,1323
73|1324,1326
199|1327,1330
/|1330,1331
100|1331,1334
18|1335,1337
95|1338,1340
%|1340,1341
RA|1342,1344
.|1344,1345
Prior|1346,1351
to|1352,1354
<EOL>|1355,1356
transfer|1356,1364
,|1364,1365
vitals|1366,1372
were|1373,1377
74|1378,1380
188|1381,1384
/|1384,1385
95|1385,1387
18|1388,1390
100|1391,1394
%|1394,1395
RA.|1396,1399
Patient|1400,1407
's|1407,1409
labs|1410,1414
were|1415,1419
<EOL>|1420,1421
remarkable|1421,1431
for|1432,1435
sodium|1436,1442
146|1443,1446
,|1446,1447
Chloride|1448,1456
115|1457,1460
,|1460,1461
K|1462,1463
5.4|1464,1467
,|1467,1468
Bicarb|1469,1475
19|1476,1478
,|1478,1479
BUN|1480,1483
<EOL>|1484,1485
39|1485,1487
,|1487,1488
Creatinine|1489,1499
2.3|1500,1503
.|1503,1504
Patient|1505,1512
had|1513,1516
CK|1517,1519
229|1520,1523
,|1523,1524
with|1525,1529
MB|1530,1532
6|1533,1534
,|1534,1535
Trop|1536,1540
<|1541,1542
0.01|1543,1547
.|1547,1548
<EOL>|1549,1550
Patient|1550,1557
had|1558,1561
BNP|1562,1565
of|1566,1568
10,180|1569,1575
.|1575,1576
Patient|1577,1584
also|1585,1589
had|1590,1593
Hgb|1594,1597
8.1|1598,1601
,|1601,1602
Hct|1603,1606
26.8|1607,1611
,|1611,1612
<EOL>|1613,1614
Platelet|1614,1622
168|1623,1626
,|1626,1627
WBC|1628,1631
5.4|1632,1635
.|1635,1636
Urinalysis|1637,1647
still|1648,1653
pending|1654,1661
upon|1662,1666
discharge|1667,1676
.|1676,1677
<EOL>|1678,1679
<EOL>|1679,1680
EKG|1680,1683
:|1683,1684
notable|1685,1692
for|1693,1696
SR|1697,1699
76|1700,1702
,|1702,1703
with|1704,1708
LAD|1709,1712
,|1712,1713
TWI|1714,1717
in|1718,1720
the|1721,1724
inferior|1725,1733
leads|1734,1739
<EOL>|1740,1741
which|1741,1746
appears|1747,1754
unchanged|1755,1764
from|1765,1769
prior|1770,1775
on|1776,1778
_|1779,1780
_|1780,1781
_|1781,1782
<EOL>|1782,1783
<EOL>|1783,1784
On|1784,1786
the|1787,1790
floor|1791,1796
she|1797,1800
is|1801,1803
symptomatically|1804,1819
improved|1820,1828
since|1829,1834
coming|1835,1841
to|1842,1844
the|1845,1848
<EOL>|1849,1850
ED|1850,1852
.|1852,1853
<EOL>|1854,1855
<EOL>|1856,1857
-|1879,1880
hypertension|1881,1893
<EOL>|1895,1896
-|1896,1897
diabetes|1898,1906
<EOL>|1908,1909
-|1909,1910
hx|1911,1913
CVA|1914,1917
(|1918,1919
cerebellar|1919,1929
-|1929,1930
medullary|1930,1939
stroke|1940,1946
in|1947,1949
_|1950,1951
_|1951,1952
_|1952,1953
<EOL>|1955,1956
-|1956,1957
CAD|1958,1961
(|1962,1963
hx|1963,1965
of|1966,1968
MI|1969,1971
in|1972,1974
_|1975,1976
_|1976,1977
_|1977,1978
BMS|1979,1982
to|1983,1985
circumflex|1986,1996
and|1997,2000
POBA|2001,2005
_|2006,2007
_|2007,2008
_|2008,2009
<EOL>|2011,2012
-|2012,2013
peripheral|2014,2024
arterial|2025,2033
disease|2034,2041
-|2041,2042
claudication|2043,2055
,|2055,2056
followed|2057,2065
by|2066,2068
<EOL>|2069,2070
vascular|2070,2078
,|2078,2079
managed|2080,2087
conservatively|2088,2102
<EOL>|2102,2103
-|2103,2104
stage|2105,2110
IV|2111,2113
CKD|2114,2117
(|2118,2119
baseline|2119,2127
2.1|2128,2131
-|2131,2132
2.6|2132,2135
)|2135,2136
<EOL>|2138,2139
-|2139,2140
GERD|2141,2145
/|2145,2146
esophageal|2146,2156
rings|2157,2162
<EOL>|2162,2163
<EOL>|2164,2165
:|2179,2180
<EOL>|2180,2181
_|2181,2182
_|2182,2183
_|2183,2184
<EOL>|2184,2185
:|2199,2200
<EOL>|2200,2201
Father|2201,2207
died|2208,2212
in|2213,2215
his|2216,2219
_|2220,2221
_|2221,2222
_|2222,2223
due|2224,2227
to|2228,2230
lung|2231,2235
disease|2236,2243
.|2243,2244
Mother|2246,2252
died|2253,2257
in|2258,2260
her|2261,2264
<EOL>|2265,2266
_|2266,2267
_|2267,2268
_|2268,2269
due|2270,2273
to|2274,2276
an|2277,2279
unknown|2280,2287
cause|2288,2293
.|2293,2294
No|2296,2298
early|2299,2304
CAD|2305,2308
or|2309,2311
sudden|2312,2318
cardiac|2319,2326
<EOL>|2327,2328
death|2328,2333
.|2333,2334
No|2335,2337
other|2338,2343
known|2344,2349
history|2350,2357
of|2358,2360
cancer|2361,2367
.|2367,2368
<EOL>|2368,2369
<EOL>|2370,2371
ADMISSION|2386,2395
PHYSICAL|2396,2404
EXAMINATION|2405,2416
:|2416,2417
<EOL>|2419,2420
VS|2420,2422
:|2422,2423
T|2424,2425
=|2425,2426
98.0|2426,2430
BP|2431,2433
:|2433,2434
168|2435,2438
/|2438,2439
96|2439,2441
HR|2442,2444
=|2444,2445
67|2445,2447
RR|2448,2450
=|2450,2451
16|2451,2453
O2|2454,2456
sat|2457,2460
=|2460,2461
100|2461,2464
%|2464,2465
on|2466,2468
2L|2469,2471
NC|2472,2474
<EOL>|2476,2477
Admission|2477,2486
weight|2487,2493
178lbs|2494,2500
<EOL>|2500,2501
GENERAL|2501,2508
:|2508,2509
WDWN|2510,2514
,|2514,2515
obese|2516,2521
,|2521,2522
sitting|2523,2530
upright|2531,2538
in|2539,2541
bed|2542,2545
,|2545,2546
in|2547,2549
NAD|2550,2553
.|2553,2554
AOx3|2555,2559
.|2559,2560
<EOL>|2561,2562
Mood|2562,2566
,|2566,2567
affect|2568,2574
appropriate|2575,2586
.|2586,2587
<EOL>|2589,2590
HEENT|2590,2595
:|2595,2596
NCAT|2597,2601
.|2601,2602
Sclera|2603,2609
anicteric|2610,2619
.|2619,2620
PERRL|2621,2626
,|2626,2627
EOMI|2628,2632
.|2632,2633
Conjunctiva|2634,2645
were|2646,2650
<EOL>|2651,2652
pink|2652,2656
,|2656,2657
no|2658,2660
pallor|2661,2667
or|2668,2670
cyanosis|2671,2679
of|2680,2682
the|2683,2686
oral|2687,2691
mucosa|2692,2698
.|2698,2699
<EOL>|2699,2700
NECK|2700,2704
:|2704,2705
Supple|2706,2712
with|2713,2717
JVP|2718,2721
of|2722,2724
8cm|2725,2728
.|2728,2729
<EOL>|2731,2732
CARDIAC|2732,2739
:|2739,2740
PMI|2741,2744
located|2745,2752
in|2753,2755
_|2756,2757
_|2757,2758
_|2758,2759
intercostal|2760,2771
space|2772,2777
,|2777,2778
midclavicular|2779,2792
<EOL>|2793,2794
line|2794,2798
.|2798,2799
RR|2800,2802
,|2802,2803
normal|2804,2810
S1|2811,2813
,|2813,2814
S2|2815,2817
,|2817,2818
+|2819,2820
S3|2820,2822
.|2822,2823
No|2824,2826
murmurs|2827,2834
/|2834,2835
rubs|2835,2839
/|2839,2840
gallops|2840,2847
.|2847,2848
No|2849,2851
<EOL>|2852,2853
thrills|2853,2860
,|2860,2861
lifts|2862,2867
.|2867,2868
<EOL>|2869,2870
LUNGS|2870,2875
:|2875,2876
Resp|2877,2881
were|2882,2886
unlabored|2887,2896
,|2896,2897
no|2898,2900
accessory|2901,2910
muscle|2911,2917
use|2918,2921
,|2921,2922
dyspneic|2923,2931
at|2932,2934
<EOL>|2935,2936
the|2936,2939
end|2940,2943
of|2944,2946
a|2947,2948
long|2949,2953
sentence|2954,2962
.|2962,2963
Bibasilar|2964,2973
crackles|2974,2982
_|2983,2984
_|2984,2985
_|2985,2986
up|2987,2989
thorax|2990,2996
,|2996,2997
<EOL>|2998,2999
diffuse|2999,3006
wheezing|3007,3015
.|3015,3016
<EOL>|3018,3019
ABDOMEN|3019,3026
:|3026,3027
Soft|3028,3032
,|3032,3033
NTND|3034,3038
.|3038,3039
No|3040,3042
HSM|3043,3046
or|3047,3049
tenderness|3050,3060
.|3060,3061
<EOL>|3063,3064
EXTREMITIES|3064,3075
:|3075,3076
2|3077,3078
+|3078,3079
edema|3080,3085
to|3086,3088
shins|3089,3094
.|3094,3095
No|3096,3098
femoral|3099,3106
bruits|3107,3113
.|3113,3114
<EOL>|3116,3117
PULSES|3117,3123
:|3123,3124
Distal|3126,3132
pulses|3133,3139
palpable|3140,3148
and|3149,3152
symmetric|3153,3162
<EOL>|3162,3163
<EOL>|3163,3164
DISCHARGE|3164,3173
PHYSICAL|3174,3182
EXAMINATION|3183,3194
:|3194,3195
<EOL>|3197,3198
VS|3198,3200
:|3200,3201
T|3202,3203
=|3203,3204
98.0|3204,3208
BP|3209,3211
:|3211,3212
135|3213,3216
/|3216,3217
72|3217,3219
HR|3220,3222
=|3222,3223
67|3223,3225
RR|3226,3228
=|3228,3229
16|3229,3231
O2|3232,3234
sat|3235,3238
=|3238,3239
100|3239,3242
%|3242,3243
on|3244,3246
RA|3247,3249
<EOL>|3249,3250
weight|3250,3256
:|3256,3257
74kg|3258,3262
<EOL>|3262,3263
GENERAL|3263,3270
:|3270,3271
WDWN|3272,3276
,|3276,3277
obese|3278,3283
,|3283,3284
sitting|3285,3292
upright|3293,3300
in|3301,3303
bed|3304,3307
,|3307,3308
in|3309,3311
NAD|3312,3315
.|3315,3316
AOx3|3317,3321
.|3321,3322
<EOL>|3323,3324
Mood|3324,3328
,|3328,3329
affect|3330,3336
appropriate|3337,3348
.|3348,3349
<EOL>|3351,3352
HEENT|3352,3357
:|3357,3358
NCAT|3359,3363
.|3363,3364
Sclera|3365,3371
anicteric|3372,3381
.|3381,3382
PERRL|3383,3388
,|3388,3389
EOMI|3390,3394
.|3394,3395
Conjunctiva|3396,3407
were|3408,3412
<EOL>|3413,3414
pink|3414,3418
,|3418,3419
no|3420,3422
pallor|3423,3429
or|3430,3432
cyanosis|3433,3441
of|3442,3444
the|3445,3448
oral|3449,3453
mucosa|3454,3460
.|3460,3461
<EOL>|3461,3462
NECK|3462,3466
:|3466,3467
Supple|3468,3474
with|3475,3479
JVP|3480,3483
of|3484,3486
7cm|3487,3490
.|3490,3491
<EOL>|3493,3494
CARDIAC|3494,3501
:|3501,3502
PMI|3503,3506
located|3507,3514
in|3515,3517
_|3518,3519
_|3519,3520
_|3520,3521
intercostal|3522,3533
space|3534,3539
,|3539,3540
midclavicular|3541,3554
<EOL>|3555,3556
line|3556,3560
.|3560,3561
RR|3562,3564
,|3564,3565
normal|3566,3572
S1|3573,3575
,|3575,3576
S2|3577,3579
,|3579,3580
+|3581,3582
S3|3582,3584
.|3584,3585
No|3586,3588
murmurs|3589,3596
/|3596,3597
rubs|3597,3601
/|3601,3602
gallops|3602,3609
.|3609,3610
No|3611,3613
<EOL>|3614,3615
thrills|3615,3622
,|3622,3623
lifts|3624,3629
.|3629,3630
<EOL>|3631,3632
LUNGS|3632,3637
:|3637,3638
Resp|3639,3643
were|3644,3648
unlabored|3649,3658
,|3658,3659
no|3660,3662
accessory|3663,3672
muscle|3673,3679
use|3680,3683
.|3683,3684
Bibasilar|3685,3694
<EOL>|3695,3696
crackles|3696,3704
trace|3705,3710
,|3710,3711
diffuse|3712,3719
wheezing|3720,3728
.|3728,3729
<EOL>|3731,3732
ABDOMEN|3732,3739
:|3739,3740
Soft|3741,3745
,|3745,3746
NTND|3747,3751
.|3751,3752
No|3753,3755
HSM|3756,3759
or|3760,3762
tenderness|3763,3773
.|3773,3774
<EOL>|3776,3777
EXTREMITIES|3777,3788
:|3788,3789
dry|3790,3793
.|3793,3794
No|3795,3797
femoral|3798,3805
bruits|3806,3812
.|3812,3813
<EOL>|3815,3816
PULSES|3816,3822
:|3822,3823
Distal|3825,3831
pulses|3832,3838
palpable|3839,3847
and|3848,3851
symmetric|3852,3861
<EOL>|3861,3862
<EOL>|3863,3864
Pertinent|3864,3873
Results|3874,3881
:|3881,3882
<EOL>|3882,3883
ADMISSION|3883,3892
LABS|3893,3897
<EOL>|3897,3898
_|3898,3899
_|3899,3900
_|3900,3901
11|3902,3904
:|3904,3905
55AM|3905,3909
BLOOD|3910,3915
WBC|3916,3919
-|3919,3920
5.4|3920,3923
RBC|3924,3927
-|3927,3928
2|3928,3929
.|3929,3930
63|3930,3932
*|3932,3933
Hgb|3934,3937
-|3937,3938
8|3938,3939
.|3939,3940
1|3940,3941
*|3941,3942
Hct|3943,3946
-|3946,3947
26|3947,3949
.|3949,3950
8|3950,3951
*|3951,3952
<EOL>|3953,3954
MCV|3954,3957
-|3957,3958
102|3958,3961
*|3961,3962
#|3962,3963
MCH|3964,3967
-|3967,3968
30.8|3968,3972
MCHC|3973,3977
-|3977,3978
30|3978,3980
.|3980,3981
2|3981,3982
*|3982,3983
RDW|3984,3987
-|3987,3988
17|3988,3990
.|3990,3991
2|3991,3992
*|3992,3993
RDWSD|3994,3999
-|3999,4000
64|4000,4002
.|4002,4003
7|4003,4004
*|4004,4005
Plt|4006,4009
_|4010,4011
_|4011,4012
_|4012,4013
<EOL>|4013,4014
_|4014,4015
_|4015,4016
_|4016,4017
11|4018,4020
:|4020,4021
55AM|4021,4025
BLOOD|4026,4031
Neuts|4032,4037
-|4037,4038
80|4038,4040
.|4040,4041
6|4041,4042
*|4042,4043
Lymphs|4044,4050
-|4050,4051
11|4051,4053
.|4053,4054
2|4054,4055
*|4055,4056
Monos|4057,4062
-|4062,4063
5.0|4063,4066
<EOL>|4067,4068
Eos|4068,4071
-|4071,4072
2.4|4072,4075
Baso|4076,4080
-|4080,4081
0.2|4081,4084
Im|4085,4087
_|4088,4089
_|4089,4090
_|4090,4091
AbsNeut|4092,4099
-|4099,4100
4|4100,4101
.|4101,4102
38|4102,4104
AbsLymp|4105,4112
-|4112,4113
0|4113,4114
.|4114,4115
61|4115,4117
*|4117,4118
<EOL>|4119,4120
AbsMono|4120,4127
-|4127,4128
0|4128,4129
.|4129,4130
27|4130,4132
AbsEos|4133,4139
-|4139,4140
0|4140,4141
.|4141,4142
13|4142,4144
AbsBaso|4145,4152
-|4152,4153
0.01|4153,4157
<EOL>|4157,4158
_|4158,4159
_|4159,4160
_|4160,4161
12|4162,4164
:|4164,4165
45PM|4165,4169
BLOOD|4170,4175
_|4176,4177
_|4177,4178
_|4178,4179
PTT|4180,4183
-|4183,4184
32.9|4184,4188
_|4189,4190
_|4190,4191
_|4191,4192
<EOL>|4192,4193
_|4193,4194
_|4194,4195
_|4195,4196
07|4197,4199
:|4199,4200
30AM|4200,4204
BLOOD|4205,4210
Ret|4211,4214
Aut|4215,4218
-|4218,4219
2|4219,4220
.|4220,4221
4|4221,4222
*|4222,4223
Abs|4224,4227
Ret|4228,4231
-|4231,4232
0.06|4232,4236
<EOL>|4236,4237
_|4237,4238
_|4238,4239
_|4239,4240
11|4241,4243
:|4243,4244
55AM|4244,4248
BLOOD|4249,4254
Glucose|4255,4262
-|4262,4263
153|4263,4266
*|4266,4267
UreaN|4268,4273
-|4273,4274
39|4274,4276
*|4276,4277
Creat|4278,4283
-|4283,4284
2|4284,4285
.|4285,4286
3|4286,4287
*|4287,4288
Na|4289,4291
-|4291,4292
146|4292,4295
*|4295,4296
<EOL>|4297,4298
K|4298,4299
-|4299,4300
5|4300,4301
.|4301,4302
4|4302,4303
*|4303,4304
Cl|4305,4307
-|4307,4308
115|4308,4311
*|4311,4312
HCO3|4313,4317
-|4317,4318
19|4318,4320
*|4320,4321
AnGap|4322,4327
-|4327,4328
17|4328,4330
<EOL>|4330,4331
_|4331,4332
_|4332,4333
_|4333,4334
11|4335,4337
:|4337,4338
55AM|4338,4342
BLOOD|4343,4348
CK|4349,4351
-|4351,4352
MB|4352,4354
-|4354,4355
6|4355,4356
cTropnT|4357,4364
-|4364,4365
<|4365,4366
0|4366,4367
.|4367,4368
01|4368,4370
_|4371,4372
_|4372,4373
_|4373,4374
<EOL>|4374,4375
_|4375,4376
_|4376,4377
_|4377,4378
07|4379,4381
:|4381,4382
38PM|4382,4386
BLOOD|4387,4392
CK|4393,4395
-|4395,4396
MB|4396,4398
-|4398,4399
6|4399,4400
cTropnT|4401,4408
-|4408,4409
<|4409,4410
0|4410,4411
.|4411,4412
01|4412,4414
<EOL>|4414,4415
_|4415,4416
_|4416,4417
_|4417,4418
11|4419,4421
:|4421,4422
55AM|4422,4426
BLOOD|4427,4432
Calcium|4433,4440
-|4440,4441
9.0|4441,4444
Phos|4445,4449
-|4449,4450
3.9|4450,4453
Mg|4454,4456
-|4456,4457
1.8|4457,4460
<EOL>|4460,4461
<EOL>|4461,4462
DISCHARGE|4462,4471
LABS|4472,4476
<EOL>|4476,4477
=|4477,4478
=|4478,4479
=|4479,4480
=|4480,4481
=|4481,4482
<EOL>|4482,4483
_|4483,4484
_|4484,4485
_|4485,4486
07|4487,4489
:|4489,4490
10AM|4490,4494
BLOOD|4495,4500
WBC|4501,4504
-|4504,4505
3|4505,4506
.|4506,4507
9|4507,4508
*|4508,4509
RBC|4510,4513
-|4513,4514
2|4514,4515
.|4515,4516
81|4516,4518
*|4518,4519
Hgb|4520,4523
-|4523,4524
8|4524,4525
.|4525,4526
6|4526,4527
*|4527,4528
Hct|4529,4532
-|4532,4533
26|4533,4535
.|4535,4536
7|4536,4537
*|4537,4538
<EOL>|4539,4540
MCV|4540,4543
-|4543,4544
95|4544,4546
MCH|4547,4550
-|4550,4551
30.6|4551,4555
MCHC|4556,4560
-|4560,4561
32.2|4561,4565
RDW|4566,4569
-|4569,4570
16|4570,4572
.|4572,4573
0|4573,4574
*|4574,4575
RDWSD|4576,4581
-|4581,4582
56|4582,4584
.|4584,4585
4|4585,4586
*|4586,4587
Plt|4588,4591
_|4592,4593
_|4593,4594
_|4594,4595
<EOL>|4595,4596
_|4596,4597
_|4597,4598
_|4598,4599
07|4600,4602
:|4602,4603
10AM|4603,4607
BLOOD|4608,4613
_|4614,4615
_|4615,4616
_|4616,4617
<EOL>|4617,4618
_|4618,4619
_|4619,4620
_|4620,4621
07|4622,4624
:|4624,4625
10AM|4625,4629
BLOOD|4630,4635
Glucose|4636,4643
-|4643,4644
100|4644,4647
UreaN|4648,4653
-|4653,4654
37|4654,4656
*|4656,4657
Creat|4658,4663
-|4663,4664
1|4664,4665
.|4665,4666
9|4666,4667
*|4667,4668
Na|4669,4671
-|4671,4672
144|4672,4675
<EOL>|4676,4677
K|4677,4678
-|4678,4679
3.9|4679,4682
Cl|4683,4685
-|4685,4686
105|4686,4689
HCO3|4690,4694
-|4694,4695
29|4695,4697
AnGap|4698,4703
-|4703,4704
14|4704,4706
<EOL>|4706,4707
_|4707,4708
_|4708,4709
_|4709,4710
07|4711,4713
:|4713,4714
10AM|4714,4718
BLOOD|4719,4724
Calcium|4725,4732
-|4732,4733
9.5|4733,4736
Phos|4737,4741
-|4741,4742
4.4|4742,4745
Mg|4746,4748
-|4748,4749
1.8|4749,4752
<EOL>|4752,4753
<EOL>|4753,4754
IMAGING|4754,4761
<EOL>|4761,4762
=|4762,4763
=|4763,4764
=|4764,4765
=|4765,4766
=|4766,4767
<EOL>|4767,4768
_|4768,4769
_|4769,4770
_|4770,4771
CXR|4772,4775
<EOL>|4775,4776
:|4784,4785
<EOL>|4786,4787
There|4787,4792
is|4793,4795
mild|4796,4800
pulmonary|4801,4810
edema|4811,4816
with|4817,4821
superimposed|4822,4834
region|4835,4841
of|4842,4844
more|4845,4849
<EOL>|4850,4851
confluent|4851,4860
consolidation|4861,4874
in|4875,4877
the|4878,4881
left|4882,4886
upper|4887,4892
lung|4893,4897
.|4897,4898
There|4900,4905
are|4906,4909
<EOL>|4910,4911
possible|4911,4919
small|4920,4925
bilateral|4926,4935
pleural|4936,4943
effusions|4944,4953
.|4953,4954
Moderate|4956,4964
<EOL>|4965,4966
cardiomegaly|4966,4978
is|4979,4981
again|4982,4987
seen|4988,4992
as|4993,4995
well|4996,5000
as|5001,5003
tortuosity|5004,5014
of|5015,5017
the|5018,5021
<EOL>|5022,5023
descending|5023,5033
thoracic|5034,5042
aorta|5043,5048
.|5048,5049
No|5051,5053
acute|5054,5059
osseous|5060,5067
abnormalities|5068,5081
.|5081,5082
<EOL>|5082,5083
<EOL>|5084,5085
Mild|5098,5102
pulmonary|5103,5112
edema|5113,5118
with|5119,5123
superimposed|5124,5136
left|5137,5141
upper|5142,5147
lung|5148,5152
<EOL>|5153,5154
consolidation|5154,5167
,|5167,5168
potentially|5169,5180
more|5181,5185
confluent|5186,5195
edema|5196,5201
versus|5202,5208
<EOL>|5209,5210
superimposed|5210,5222
infection|5223,5232
.|5232,5233
<EOL>|5233,5234
<EOL>|5234,5235
<EOL>|5236,5237
_|5260,5261
_|5261,5262
_|5262,5263
year|5264,5268
-|5268,5269
old|5269,5272
female|5273,5279
with|5280,5284
history|5285,5292
of|5293,5295
hypertension|5296,5308
,|5308,5309
CAD|5310,5313
s|5314,5315
/|5315,5316
p|5316,5317
DES|5318,5321
<EOL>|5322,5323
with|5323,5327
ischemic|5328,5336
MR|5337,5339
and|5340,5343
systolic|5344,5352
dysfunction|5353,5364
,|5364,5365
_|5366,5367
_|5367,5368
_|5368,5369
,|5369,5370
hx|5371,5373
of|5374,5376
DVT|5377,5380
,|5380,5381
who|5382,5385
<EOL>|5386,5387
admitted|5387,5395
for|5396,5399
CHF|5400,5403
exacerbation|5404,5416
.|5416,5417
<EOL>|5417,5418
<EOL>|5418,5419
#|5419,5420
Acute|5421,5426
on|5427,5429
chronic|5430,5437
decompensated|5438,5451
heart|5452,5457
failure|5458,5465
:|5465,5466
presented|5467,5476
in|5477,5479
the|5480,5483
<EOL>|5484,5485
setting|5485,5492
of|5493,5495
high|5496,5500
salt|5501,5505
diet|5506,5510
with|5511,5515
dyspnea|5516,5523
on|5524,5526
exertion|5527,5535
,|5535,5536
decreased|5537,5546
<EOL>|5547,5548
exercise|5548,5556
tolerance|5557,5566
,|5566,5567
_|5568,5569
_|5569,5570
_|5570,5571
edema|5572,5577
,|5577,5578
crackles|5579,5587
on|5588,5590
exam|5591,5595
,|5595,5596
elevated|5597,5605
BNP|5606,5609
to|5610,5612
<EOL>|5613,5614
10K|5614,5617
,|5617,5618
8lbs|5619,5623
above|5624,5629
dry|5630,5633
weight|5634,5640
and|5641,5644
pulmonary|5645,5654
congestion|5655,5665
on|5666,5668
CXR|5669,5672
.|5672,5673
<EOL>|5674,5675
Later|5675,5680
discovered|5681,5691
on|5692,5694
pharmacy|5695,5703
review|5704,5710
that|5711,5715
patient|5716,5723
had|5724,5727
not|5728,5731
filled|5732,5738
<EOL>|5739,5740
torsemide|5740,5749
after|5750,5755
last|5756,5760
outpatient|5761,5771
Cardiology|5772,5782
appointment|5783,5794
where|5795,5800
she|5801,5804
<EOL>|5805,5806
was|5806,5809
instructed|5810,5820
to|5821,5823
start|5824,5829
taking|5830,5836
it|5837,5839
.|5839,5840
Troponins|5841,5850
cycled|5851,5857
and|5858,5861
<EOL>|5862,5863
negative|5863,5871
.|5871,5872
On|5873,5875
admission|5876,5885
,|5885,5886
she|5887,5890
was|5891,5894
placed|5895,5901
on|5902,5904
a|5905,5906
salt|5907,5911
and|5912,5915
fluid|5916,5921
<EOL>|5922,5923
restricted|5923,5933
diet|5934,5938
.|5938,5939
She|5940,5943
was|5944,5947
diuresed|5948,5956
with|5957,5961
IV|5962,5964
Lasix|5965,5970
80mg|5971,5975
for|5976,5979
2|5980,5981
days|5982,5986
<EOL>|5987,5988
and|5988,5991
then|5992,5996
transitioned|5997,6009
to|6010,6012
po|6013,6015
torsemide|6016,6025
40mg|6026,6030
with|6031,6035
steady|6036,6042
weight|6043,6049
<EOL>|6050,6051
decline|6051,6058
and|6059,6062
net|6063,6066
negative|6067,6075
fluid|6076,6081
balance|6082,6089
of|6090,6092
goal|6093,6097
-|6098,6099
_|6099,6100
_|6100,6101
_|6101,6102
and|6103,6106
<EOL>|6107,6108
stable|6108,6114
renal|6115,6120
function|6121,6129
.|6129,6130
Electrolytes|6131,6143
repleted|6144,6152
for|6153,6156
goal|6157,6161
Mg|6162,6164
>|6164,6165
2|6165,6166
and|6167,6170
<EOL>|6171,6172
K|6172,6173
>|6173,6174
4|6174,6175
.|6175,6176
She|6177,6180
was|6181,6184
continued|6185,6194
on|6195,6197
home|6198,6202
carvedilol|6203,6213
12.5|6214,6218
mg|6218,6220
BID|6221,6224
,|6224,6225
<EOL>|6226,6227
atorvastatin|6227,6239
80mg|6240,6244
daily|6245,6250
and|6251,6254
lisinopril|6255,6265
40mg|6266,6270
daily|6271,6276
for|6277,6280
blood|6281,6286
<EOL>|6287,6288
pressure|6288,6296
control|6297,6304
and|6305,6308
increased|6309,6318
home|6319,6323
nifedipine|6324,6334
CR|6335,6337
from|6338,6342
30|6343,6345
to|6346,6348
<EOL>|6349,6350
60mg|6350,6354
BID|6355,6358
to|6359,6361
achieve|6362,6369
goal|6370,6374
SBP|6375,6378
<|6379,6380
140|6380,6383
.|6383,6384
Discharged|6385,6395
with|6396,6400
close|6401,6406
PCP|6407,6410
and|6411,6414
<EOL>|6415,6416
_|6416,6417
_|6417,6418
_|6418,6419
to|6420,6422
monitor|6423,6430
weights|6431,6438
and|6439,6442
blood|6443,6448
pressure|6449,6457
<EOL>|6458,6459
control|6459,6466
.|6466,6467
<EOL>|6467,6468
<EOL>|6468,6469
#|6469,6470
Hypertension|6471,6483
:|6483,6484
She|6485,6488
was|6489,6492
continued|6493,6502
on|6503,6505
home|6506,6510
carvedilol|6511,6521
12.5|6522,6526
mg|6526,6528
BID|6529,6532
,|6532,6533
<EOL>|6534,6535
atorvastatin|6535,6547
80mg|6548,6552
daily|6553,6558
and|6559,6562
lisinopril|6563,6573
40mg|6574,6578
daily|6579,6584
for|6585,6588
blood|6589,6594
<EOL>|6595,6596
pressure|6596,6604
control|6605,6612
and|6613,6616
increased|6617,6626
home|6627,6631
nifedipine|6632,6642
CR|6643,6645
from|6646,6650
30|6651,6653
to|6654,6656
<EOL>|6657,6658
60mg|6658,6662
BID|6663,6666
to|6667,6669
achieve|6670,6677
goal|6678,6682
SBP|6683,6686
<|6687,6688
140|6688,6691
.|6691,6692
<EOL>|6693,6694
<EOL>|6694,6695
#|6695,6696
Positive|6697,6705
U|6706,6707
/|6707,6708
A|6708,6709
:|6709,6710
patient|6711,6718
asymptomatic|6719,6731
but|6732,6735
with|6736,6740
32WBCs|6741,6747
,|6747,6748
_|6749,6750
_|6750,6751
_|6751,6752
,|6752,6753
<EOL>|6754,6755
+|6755,6756
bacteria|6756,6764
(|6765,6766
although|6766,6774
3|6775,6776
epis|6777,6781
)|6781,6782
.|6782,6783
Asymptomatic|6784,6796
with|6797,6801
no|6802,6804
<EOL>|6805,6806
fevers|6806,6812
/|6812,6813
dysuria|6813,6820
/|6820,6821
malaise|6821,6828
.|6828,6829
Urine|6830,6835
culture|6836,6843
negative|6844,6852
.|6852,6853
<EOL>|6853,6854
<EOL>|6854,6855
#|6855,6856
Left|6857,6861
upper|6862,6867
lung|6868,6872
consolidation|6873,6886
:|6886,6887
infiltrate|6888,6898
per|6899,6902
Radiology|6903,6912
read|6913,6917
<EOL>|6918,6919
on|6919,6921
admission|6922,6931
CXR|6932,6935
.|6935,6936
No|6937,6939
cough|6940,6945
,|6945,6946
fevers|6947,6953
,|6953,6954
leukocytosis|6955,6967
.|6967,6968
Rereviewed|6969,6979
<EOL>|6980,6981
with|6981,6985
on|6986,6988
-|6988,6989
call|6989,6993
radiologist|6994,7005
who|7006,7009
favored|7010,7017
pulmonary|7018,7027
edema|7028,7033
with|7034,7038
no|7039,7041
<EOL>|7042,7043
need|7043,7047
for|7048,7051
repeat|7052,7058
imaging|7059,7066
or|7067,7069
PNA|7070,7073
treatment|7074,7083
unless|7084,7090
clinically|7091,7101
<EOL>|7102,7103
indicated|7103,7112
.|7112,7113
Monitored|7114,7123
without|7124,7131
any|7132,7135
significant|7136,7147
clinical|7148,7156
findings|7157,7165
.|7165,7166
<EOL>|7166,7167
<EOL>|7167,7168
#|7168,7169
DVT|7170,7173
:|7173,7174
anticoagulated|7175,7189
on|7190,7192
Coumadin|7193,7201
goal|7202,7206
2.0|7207,7210
-|7210,7211
3|7211,7212
.|7212,7213
0|7213,7214
,|7214,7215
no|7216,7218
signs|7219,7224
of|7225,7227
<EOL>|7228,7229
thrombus|7229,7237
on|7238,7240
exam|7241,7245
.|7245,7246
Daily|7247,7252
INR|7253,7256
trended|7257,7264
and|7265,7268
continued|7269,7278
on|7279,7281
home|7282,7286
<EOL>|7287,7288
Coumadin|7288,7296
5mg|7297,7300
daily|7301,7306
.|7306,7307
<EOL>|7308,7309
<EOL>|7309,7310
#|7310,7311
Anemia|7312,7318
:|7318,7319
no|7320,7322
signs|7323,7328
of|7329,7331
external|7332,7340
loss|7341,7345
,|7345,7346
specifically|7347,7359
denying|7360,7367
any|7368,7371
<EOL>|7372,7373
melena|7373,7379
.|7379,7380
Chronically|7381,7392
anemic|7393,7399
with|7400,7404
baseline|7405,7413
_|7414,7415
_|7415,7416
_|7416,7417
,|7417,7418
presented|7419,7428
with|7429,7433
Hgb|7434,7437
<EOL>|7438,7439
8.|7439,7441
Likely|7442,7448
_|7449,7450
_|7450,7451
_|7451,7452
renal|7453,7458
disease|7459,7466
and|7467,7470
ACD|7471,7474
however|7475,7482
elevated|7483,7491
MCV|7492,7495
<EOL>|7496,7497
indicates|7497,7506
possible|7507,7515
reticulocytosis|7516,7531
.|7531,7532
Altogether|7533,7543
low|7544,7547
suspicion|7548,7557
for|7558,7561
<EOL>|7562,7563
GIB|7563,7566
so|7567,7569
Coumadin|7570,7578
was|7579,7582
continued|7583,7592
.|7592,7593
Reticulocytes|7594,7607
2.4|7608,7611
which|7612,7617
is|7618,7620
<EOL>|7621,7622
inappropriate|7622,7635
arguing|7636,7643
against|7644,7651
acute|7652,7657
loss|7658,7662
.|7662,7663
Trended|7664,7671
daily|7672,7677
CBC|7678,7681
with|7682,7686
<EOL>|7687,7688
noted|7688,7693
uprising|7694,7702
by|7703,7705
discharge|7706,7715
.|7715,7716
<EOL>|7716,7717
<EOL>|7717,7718
#|7718,7719
Chronic|7720,7727
kidney|7728,7734
disease|7735,7742
,|7742,7743
stage|7744,7749
IV|7750,7752
-|7752,7753
baseline|7754,7762
_|7763,7764
_|7764,7765
_|7765,7766
,|7766,7767
likely|7768,7774
_|7775,7776
_|7776,7777
_|7777,7778
<EOL>|7779,7780
HTN|7780,7783
and|7784,7787
DM|7788,7790
.|7790,7791
Renally|7792,7799
dosed|7800,7805
medications|7806,7817
and|7818,7821
trended|7822,7829
Cr|7830,7832
with|7833,7837
no|7838,7840
<EOL>|7841,7842
significant|7842,7853
change|7854,7860
.|7860,7861
<EOL>|7862,7863
#|7863,7864
HLD|7865,7868
:|7868,7869
continued|7870,7879
home|7880,7884
atorvastatin|7885,7897
<EOL>|7897,7898
#|7898,7899
DM|7900,7902
:|7902,7903
held|7904,7908
home|7909,7913
25U|7914,7917
70|7918,7920
/|7920,7921
30|7921,7923
.|7923,7924
Patient|7926,7933
maintained|7934,7944
on|7945,7947
aspart|7948,7954
ISS|7955,7958
and|7959,7962
<EOL>|7963,7964
glargine|7964,7972
qHS|7973,7976
with|7977,7981
good|7982,7986
glycemic|7987,7995
control|7996,8003
.|8003,8004
<EOL>|8004,8005
<EOL>|8005,8006
TRANSITIONAL|8006,8018
ISSUES|8019,8025
<EOL>|8025,8026
=|8026,8027
=|8027,8028
=|8028,8029
=|8029,8030
=|8030,8031
=|8031,8032
=|8032,8033
=|8033,8034
=|8034,8035
=|8035,8036
=|8036,8037
=|8037,8038
=|8038,8039
=|8039,8040
=|8040,8041
=|8041,8042
=|8042,8043
=|8043,8044
<EOL>|8044,8045
CHF|8045,8048
:|8048,8049
diuresed|8050,8058
with|8059,8063
IV|8064,8066
lasix|8067,8072
,|8072,8073
transitioned|8074,8086
to|8087,8089
po|8090,8092
diuretics|8093,8102
,|8102,8103
<EOL>|8104,8105
discharged|8105,8115
home|8116,8120
on|8121,8123
40mg|8124,8128
po|8129,8131
torsemide|8132,8141
,|8141,8142
to|8143,8145
take|8146,8150
in|8151,8153
the|8154,8157
AM|8158,8160
and|8161,8164
take|8165,8169
<EOL>|8170,8171
a|8171,8172
banana|8173,8179
.|8179,8180
Pt|8181,8183
complained|8184,8194
of|8195,8197
unilateral|8198,8208
R|8209,8210
-|8210,8211
sided|8211,8216
incomplete|8217,8227
hearing|8228,8235
<EOL>|8236,8237
loss|8237,8241
on|8242,8244
day|8245,8248
of|8249,8251
discharge|8252,8261
-|8261,8262
was|8263,8266
not|8267,8270
felt|8271,8275
to|8276,8278
be|8279,8281
related|8282,8289
to|8290,8292
<EOL>|8293,8294
diuretics|8294,8303
but|8304,8307
would|8308,8313
_|8314,8315
_|8315,8316
_|8316,8317
.|8317,8318
<EOL>|8318,8319
HTN|8319,8322
:|8322,8323
increased|8324,8333
nifedipine|8334,8344
CR|8345,8347
to|8348,8350
60mg|8351,8355
BID|8356,8359
given|8360,8365
elevated|8366,8374
SBPs|8375,8379
.|8379,8380
<EOL>|8381,8382
Please|8382,8388
f|8389,8390
/|8390,8391
u|8391,8392
at|8393,8395
next|8396,8400
appointments|8401,8413
.|8413,8414
<EOL>|8414,8415
Anemia|8415,8421
:|8421,8422
multiple|8423,8431
prior|8432,8437
workups|8438,8445
showing|8446,8453
ACD|8454,8457
.|8457,8458
Hgb|8459,8462
8s|8463,8465
during|8466,8472
<EOL>|8473,8474
admission|8474,8483
<EOL>|8483,8484
Prior|8484,8489
DVT|8490,8493
/|8493,8494
PE|8494,8496
:|8496,8497
continued|8498,8507
on|8508,8510
warfarin|8511,8519
,|8519,8520
will|8521,8525
need|8526,8530
continued|8531,8540
<EOL>|8541,8542
monitoring|8542,8552
<EOL>|8552,8553
DM|8553,8555
:|8555,8556
stopped|8557,8564
home|8565,8569
70|8570,8572
/|8572,8573
30|8573,8575
while|8576,8581
in|8582,8584
-|8584,8585
house|8585,8590
and|8591,8594
put|8595,8598
on|8599,8601
<EOL>|8602,8603
aspart|8603,8609
/|8609,8610
glargine|8610,8618
,|8618,8619
discharged|8620,8630
on|8631,8633
home|8634,8638
regimen|8639,8646
<EOL>|8646,8647
<EOL>|8647,8648
Discharge|8648,8657
weight|8658,8664
:|8664,8665
74kg|8666,8670
<EOL>|8670,8671
Discharge|8671,8680
Cr|8681,8683
:|8683,8684
1.9|8685,8688
<EOL>|8688,8689
<EOL>|8690,8691
Medications|8691,8702
on|8703,8705
Admission|8706,8715
:|8715,8716
<EOL>|8716,8717
The|8717,8720
Preadmission|8721,8733
Medication|8734,8744
list|8745,8749
is|8750,8752
accurate|8753,8761
and|8762,8765
complete|8766,8774
.|8774,8775
<EOL>|8775,8776
1.|8776,8778
Acetaminophen|8779,8792
325|8793,8796
-|8796,8797
650|8797,8800
mg|8801,8803
PO|8804,8806
Q6H|8807,8810
:|8810,8811
PRN|8811,8814
pain|8815,8819
or|8820,8822
fever|8823,8828
<EOL>|8829,8830
2.|8830,8832
Aspirin|8833,8840
81|8841,8843
mg|8844,8846
PO|8847,8849
DAILY|8850,8855
<EOL>|8856,8857
3.|8857,8859
Atorvastatin|8860,8872
80|8873,8875
mg|8876,8878
PO|8879,8881
QPM|8882,8885
<EOL>|8886,8887
4.|8887,8889
Carvedilol|8890,8900
12.5|8901,8905
mg|8906,8908
PO|8909,8911
BID|8912,8915
<EOL>|8916,8917
5.|8917,8919
Docusate|8920,8928
Sodium|8929,8935
100|8936,8939
mg|8940,8942
PO|8943,8945
BID|8946,8949
<EOL>|8950,8951
6.|8951,8953
Gabapentin|8954,8964
100|8965,8968
mg|8969,8971
PO|8972,8974
QHS|8975,8978
neuropathic|8979,8990
pain|8991,8995
<EOL>|8996,8997
7.|8997,8999
Lisinopril|9000,9010
40|9011,9013
mg|9014,9016
PO|9017,9019
DAILY|9020,9025
<EOL>|9026,9027
8.|9027,9029
Multivitamins|9030,9043
1|9044,9045
TAB|9046,9049
PO|9050,9052
DAILY|9053,9058
<EOL>|9059,9060
9.|9060,9062
NIFEdipine|9063,9073
CR|9074,9076
30|9077,9079
mg|9080,9082
PO|9083,9085
BID|9086,9089
<EOL>|9090,9091
10.|9091,9094
Nitroglycerin|9095,9108
SL|9109,9111
0.3|9112,9115
mg|9116,9118
SL|9119,9121
Q5MIN|9122,9127
:|9127,9128
PRN|9128,9131
chest|9132,9137
pain|9138,9142
<EOL>|9143,9144
11|9144,9146
.|9146,9147
Pantoprazole|9148,9160
40|9161,9163
mg|9164,9166
PO|9167,9169
Q12H|9170,9174
<EOL>|9175,9176
12.|9176,9179
Polyethylene|9180,9192
Glycol|9193,9199
17|9200,9202
g|9203,9204
PO|9205,9207
DAILY|9208,9213
<EOL>|9214,9215
13.|9215,9218
Senna|9219,9224
8.6|9225,9228
mg|9229,9231
PO|9232,9234
BID|9235,9238
constipation|9239,9251
<EOL>|9252,9253
14.|9253,9256
Vitamin|9257,9264
D|9265,9266
_|9267,9268
_|9268,9269
_|9269,9270
UNIT|9271,9275
PO|9276,9278
DAILY|9279,9284
<EOL>|9285,9286
15.|9286,9289
Warfarin|9290,9298
5|9299,9300
mg|9301,9303
PO|9304,9306
DAILY16|9307,9314
<EOL>|9315,9316
16|9316,9318
.|9318,9319
Allopurinol|9320,9331
_|9332,9333
_|9333,9334
_|9334,9335
mg|9336,9338
PO|9339,9341
EVERY|9342,9347
OTHER|9348,9353
DAY|9354,9357
<EOL>|9358,9359
17.|9359,9362
Torsemide|9363,9372
40|9373,9375
mg|9376,9378
PO|9379,9381
DAILY|9382,9387
<EOL>|9388,9389
18.|9389,9392
HumuLIN|9393,9400
70|9401,9403
/|9403,9404
30|9404,9406
(|9407,9408
insulin|9408,9415
NPH|9416,9419
and|9420,9423
regular|9424,9431
human|9432,9437
)|9437,9438
100|9439,9442
unit|9443,9447
/|9447,9448
mL|9448,9450
<EOL>|9451,9452
(|9452,9453
70|9453,9455
-|9455,9456
30|9456,9458
)|9458,9459
subcutaneous|9460,9472
25|9473,9475
units|9476,9481
with|9482,9486
dinner|9487,9493
<EOL>|9494,9495
<EOL>|9495,9496
<EOL>|9497,9498
Discharge|9498,9507
Medications|9508,9519
:|9519,9520
<EOL>|9520,9521
1.|9521,9523
HumuLIN|9524,9531
70|9532,9534
/|9534,9535
30|9535,9537
(|9538,9539
insulin|9539,9546
NPH|9547,9550
and|9551,9554
regular|9555,9562
human|9563,9568
)|9568,9569
100|9570,9573
unit|9574,9578
/|9578,9579
mL|9579,9581
<EOL>|9582,9583
(|9583,9584
70|9584,9586
-|9586,9587
30|9587,9589
)|9589,9590
subcutaneous|9591,9603
25|9604,9606
units|9607,9612
with|9613,9617
dinner|9618,9624
<EOL>|9625,9626
2.|9626,9628
Warfarin|9629,9637
5|9638,9639
mg|9640,9642
PO|9643,9645
DAILY16|9646,9653
<EOL>|9654,9655
3.|9655,9657
Vitamin|9658,9665
D|9666,9667
_|9668,9669
_|9669,9670
_|9670,9671
UNIT|9672,9676
PO|9677,9679
DAILY|9680,9685
<EOL>|9686,9687
4.|9687,9689
Acetaminophen|9690,9703
325|9704,9707
-|9707,9708
650|9708,9711
mg|9712,9714
PO|9715,9717
Q6H|9718,9721
:|9721,9722
PRN|9722,9725
pain|9726,9730
or|9731,9733
fever|9734,9739
<EOL>|9740,9741
5.|9741,9743
Allopurinol|9744,9755
_|9756,9757
_|9757,9758
_|9758,9759
mg|9760,9762
PO|9763,9765
EVERY|9766,9771
OTHER|9772,9777
DAY|9778,9781
<EOL>|9782,9783
6.|9783,9785
Aspirin|9786,9793
81|9794,9796
mg|9797,9799
PO|9800,9802
DAILY|9803,9808
<EOL>|9809,9810
7.|9810,9812
Atorvastatin|9813,9825
80|9826,9828
mg|9829,9831
PO|9832,9834
QPM|9835,9838
<EOL>|9839,9840
8.|9840,9842
Docusate|9843,9851
Sodium|9852,9858
100|9859,9862
mg|9863,9865
PO|9866,9868
BID|9869,9872
<EOL>|9873,9874
9.|9874,9876
Gabapentin|9877,9887
100|9888,9891
mg|9892,9894
PO|9895,9897
QHS|9898,9901
neuropathic|9902,9913
pain|9914,9918
<EOL>|9919,9920
10|9920,9922
.|9922,9923
Lisinopril|9924,9934
40|9935,9937
mg|9938,9940
PO|9941,9943
DAILY|9944,9949
<EOL>|9950,9951
11.|9951,9954
Multivitamins|9955,9968
1|9969,9970
TAB|9971,9974
PO|9975,9977
DAILY|9978,9983
<EOL>|9984,9985
12.|9985,9988
Nitroglycerin|9989,10002
SL|10003,10005
0.3|10006,10009
mg|10010,10012
SL|10013,10015
Q5MIN|10016,10021
:|10021,10022
PRN|10022,10025
chest|10026,10031
pain|10032,10036
<EOL>|10037,10038
13|10038,10040
.|10040,10041
Polyethylene|10042,10054
Glycol|10055,10061
17|10062,10064
g|10065,10066
PO|10067,10069
DAILY|10070,10075
<EOL>|10076,10077
14.|10077,10080
Senna|10081,10086
8.6|10087,10090
mg|10091,10093
PO|10094,10096
BID|10097,10100
constipation|10101,10113
<EOL>|10114,10115
15.|10115,10118
Torsemide|10119,10128
40|10129,10131
mg|10132,10134
PO|10135,10137
DAILY|10138,10143
<EOL>|10144,10145
RX|10145,10147
*|10148,10149
torsemide|10149,10158
20|10159,10161
mg|10162,10164
2|10165,10166
tablet|10167,10173
(|10173,10174
s|10174,10175
)|10175,10176
by|10177,10179
mouth|10180,10185
once|10186,10190
daily|10191,10196
Disp|10197,10201
#|10202,10203
*|10203,10204
60|10204,10206
<EOL>|10207,10208
Tablet|10208,10214
Refills|10215,10222
:|10222,10223
*|10223,10224
0|10224,10225
<EOL>|10225,10226
16|10226,10228
.|10228,10229
Pantoprazole|10230,10242
20|10243,10245
mg|10246,10248
PO|10249,10251
Q12H|10252,10256
<EOL>|10257,10258
17.|10258,10261
Carvedilol|10262,10272
25|10273,10275
mg|10276,10278
PO|10279,10281
BID|10282,10285
<EOL>|10286,10287
18.|10287,10290
NIFEdipine|10291,10301
CR|10302,10304
60|10305,10307
mg|10308,10310
PO|10311,10313
BID|10314,10317
<EOL>|10318,10319
RX|10319,10321
*|10322,10323
nifedipine|10323,10333
20|10334,10336
mg|10337,10339
3|10340,10341
capsule|10342,10349
(|10349,10350
s|10350,10351
)|10351,10352
by|10353,10355
mouth|10356,10361
twice|10362,10367
daily|10368,10373
Disp|10374,10378
<EOL>|10379,10380
#|10380,10381
*|10381,10382
180|10382,10385
Capsule|10386,10393
Refills|10394,10401
:|10401,10402
*|10402,10403
0|10403,10404
<EOL>|10404,10405
<EOL>|10405,10406
<EOL>|10407,10408
Discharge|10408,10417
Disposition|10418,10429
:|10429,10430
<EOL>|10430,10431
Home|10431,10435
With|10436,10440
Service|10441,10448
<EOL>|10448,10449
<EOL>|10450,10451
Facility|10451,10459
:|10459,10460
<EOL>|10460,10461
_|10461,10462
_|10462,10463
_|10463,10464
<EOL>|10464,10465
<EOL>|10466,10467
Discharge|10467,10476
Diagnosis|10477,10486
:|10486,10487
<EOL>|10487,10488
Acute|10507,10512
on|10513,10515
chronic|10516,10523
decompensated|10524,10537
congestive|10538,10548
Heart|10549,10554
Failure|10555,10562
<EOL>|10562,10563
Hypertension|10563,10575
<EOL>|10575,10576
<EOL>|10576,10577
Secondary|10577,10586
Diagnoses|10587,10596
:|10596,10597
<EOL>|10597,10598
Anemia|10598,10604
<EOL>|10604,10605
Diabetes|10605,10613
mellitus|10614,10622
<EOL>|10622,10623
Prior|10623,10628
deep|10629,10633
vein|10634,10638
thrombosis|10639,10649
<EOL>|10649,10650
Chronic|10650,10657
Kidney|10658,10664
Disease|10665,10672
<EOL>|10672,10673
<EOL>|10673,10674
<EOL>|10675,10676
Mental|10697,10703
Status|10704,10710
:|10710,10711
Clear|10712,10717
and|10718,10721
coherent|10722,10730
.|10730,10731
<EOL>|10731,10732
Level|10732,10737
of|10738,10740
Consciousness|10741,10754
:|10754,10755
Alert|10756,10761
and|10762,10765
interactive|10766,10777
.|10777,10778
<EOL>|10778,10779
Activity|10779,10787
Status|10788,10794
:|10794,10795
Ambulatory|10796,10806
-|10807,10808
Independent|10809,10820
.|10820,10821
<EOL>|10821,10822
<EOL>|10822,10823
<EOL>|10824,10825
Mrs.|10849,10853
_|10854,10855
_|10855,10856
_|10856,10857
,|10857,10858
<EOL>|10859,10860
<EOL>|10860,10861
_|10861,10862
_|10862,10863
_|10863,10864
were|10865,10869
admitted|10870,10878
to|10879,10881
_|10882,10883
_|10883,10884
_|10884,10885
for|10886,10889
treatment|10890,10899
of|10900,10902
your|10903,10907
congestive|10908,10918
<EOL>|10919,10920
heart|10920,10925
failure|10926,10933
and|10934,10937
hypertension|10938,10950
.|10950,10951
_|10952,10953
_|10953,10954
_|10954,10955
were|10956,10960
given|10961,10966
IV|10967,10969
diuretics|10970,10979
with|10980,10984
<EOL>|10985,10986
improvement|10986,10997
in|10998,11000
your|11001,11005
symptoms|11006,11014
,|11014,11015
labs|11016,11020
and|11021,11024
exam|11025,11029
.|11029,11030
We|11031,11033
increased|11034,11043
one|11044,11047
of|11048,11050
<EOL>|11051,11052
your|11052,11056
blood|11057,11062
pressure|11063,11071
medications|11072,11083
and|11084,11087
continued|11088,11097
your|11098,11102
other|11103,11108
home|11109,11113
<EOL>|11114,11115
medicines|11115,11124
.|11124,11125
<EOL>|11126,11127
<EOL>|11127,11128
It|11128,11130
was|11131,11134
a|11135,11136
pleasure|11137,11145
taking|11146,11152
care|11153,11157
of|11158,11160
_|11161,11162
_|11162,11163
_|11163,11164
during|11165,11171
your|11172,11176
stay|11177,11181
-|11181,11182
we|11183,11185
wish|11186,11190
<EOL>|11191,11192
_|11192,11193
_|11193,11194
_|11194,11195
all|11196,11199
the|11200,11203
best|11204,11208
!|11208,11209
<EOL>|11209,11210
<EOL>|11210,11211
-|11211,11212
Your|11213,11217
_|11218,11219
_|11219,11220
_|11220,11221
Team|11222,11226
<EOL>|11226,11227
<EOL>|11228,11229
Followup|11229,11237
Instructions|11238,11250
:|11250,11251
<EOL>|11251,11252
_|11252,11253
_|11253,11254
_|11254,11255
<EOL>|11255,11256

