CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Orthopedics|Title|false|false||ORTHOPAEDICSnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|INJECTION, MEROPENEM, 100 MG ADMINISTERED|Drug|false|false||meropenem
null|meropenem|Drug|false|false||meropenem
null|meropenem|Drug|false|false||meropenemnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Chief complaint (finding)|Finding|false|false||Chief Complaintnull|Complaint (finding)|Finding|false|false||Complaintnull|null|Attribute|false|false||Complaintnull|Pain of left hip joint|Finding|false|false|C0524471;C0022122;C0228391;C0019552;C4299095|left hip painnull|Left hip region structure|Anatomy|false|false|C0019559;C4551516;C1552822;C1292890;C2141922;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1549543;C0030193|left hipnull|Table Cell Horizontal Align - left|Finding|false|false|C0524471|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Hip joint pain|Finding|false|false|C0524471;C0022122;C0228391;C0019552;C4299095|hip pain
null|Hip pain|Finding|false|false|C0524471;C0022122;C0228391;C0019552;C4299095|hip painnull|null|Attribute|false|false|C0022122;C0228391;C0019552;C4299095|hip painnull|heme iron polypeptide|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|ST13 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|ST13 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|RPL29 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|RPL29 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|HHIP protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|HHIP protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|heme iron polypeptide|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hipnull|RPL29 wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C0524471|hip
null|REG3A gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C0524471|hip
null|RPL29 gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C0524471|hip
null|ST13 wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C0524471|hip
null|ST13 gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C0524471|hip
null|HHIP gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C0524471|hip
null|HHIP wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C0524471|hip
null|REG3A wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C0524471|hipnull|Procedure on hip|Procedure|false|false|C0524471;C0022122;C0228391;C0019552;C4299095|hipnull|Lower extremity>Hip|Anatomy|false|false|C1549543;C0030193;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C0019559;C4551516;C1292890;C1430701;C0529134;C1505163;C1654726;C1716793;C2141922|hip
null|Hip structure|Anatomy|false|false|C1549543;C0030193;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C0019559;C4551516;C1292890;C1430701;C0529134;C1505163;C1654726;C1716793;C2141922|hip
null|Structure of habenulopeduncular tract|Anatomy|false|false|C1549543;C0030193;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C0019559;C4551516;C1292890;C1430701;C0529134;C1505163;C1654726;C1716793;C2141922|hip
null|Bone structure of ischium|Anatomy|false|false|C1549543;C0030193;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C0019559;C4551516;C1292890;C1430701;C0529134;C1505163;C1654726;C1716793;C2141922|hipnull|Administration Method - Pain|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C0524471|pain
null|Pain|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C0524471|painnull|null|Attribute|false|false||painnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Reduced|Finding|false|false||reductionnull|Reduction procedure|Procedure|false|false||reduction
null|Surgical reduction|Procedure|false|false||reductionnull|Reduction (chemical)|Phenomenon|false|false||reductionnull|Percutaneous Route of Drug Administration|Finding|false|false||percutaneousnull|Percutaneous|Modifier|false|false||percutaneousnull|Intramedullary Nailing|Procedure|false|false||pinningnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Femoral Neck Fractures|Disorder|false|false|C0027530;C3159206;C0015811;C0015815|femoral neck fracturenull|Structure of neck of femur|Anatomy|false|false|C0262414;C0016658;C0812434;C0684335;C0015806|femoral necknull|Femur|Anatomy|false|false|C0015806;C0262414;C0016658|femoralnull|Fracture of cervical spine|Disorder|false|false|C0015815;C0015811;C0027530;C3159206|neck fracturenull|Passive joint movement of neck (finding)|Finding|false|false|C0015815;C0027530;C3159206|neck
null|Neck problem|Finding|false|false|C0015815;C0027530;C3159206|necknull|dendritic spine neck|Anatomy|false|false|C0015806;C0016658;C0262414;C0812434;C0684335|neck
null|Neck|Anatomy|false|false|C0015806;C0016658;C0262414;C0812434;C0684335|necknull|Fracture|Disorder|false|false|C0015815;C0027530;C3159206;C0015811|fracturenull|History of present illness (finding)|Finding|false|false||History of Present Illnessnull|null|Attribute|false|false||History of Present Illnessnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Present illness|Finding|false|false||Present Illnessnull|Present|Finding|false|false||Present
null|Presentation|Finding|false|false||Presentnull|Illness (finding)|Finding|false|false||Illnessnull|Woman|Subject|false|false||woman
null|Human, Female adult|Subject|false|false||womannull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Presentation|Finding|false|false||presentationnull|mechanical method|Finding|false|false||mechanicalnull|Mechanical Treatments|Procedure|false|false||mechanicalnull|Falls|Finding|false|false||fallnull|Autumn|Time|false|false||fallnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Body Site Modifier - Lower|Anatomy|false|false|C2003888|lowernull|Lower (action)|Event|false|false|C1548802|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Limb structure|Anatomy|false|false|C2598155;C1548167;C1697779;C4036205;C1549543;C0030193;C5436357|extremitynull|Query Priority - Immediate|Finding|false|false|C0015385|immediate
null|immediate - ResponseCode|Finding|false|false|C0015385|immediatenull|Immediate|Time|false|false||immediate
null|Stat (do immediately)|Time|false|false||immediatenull|Administration Method - Pain|Finding|false|false|C0015385|pain
null|Pain|Finding|false|false|C0015385|painnull|null|Attribute|false|false|C0015385|painnull|Inability to ambulate|Finding|false|false|C0015385|inability to ambulatenull|Ambulate|Finding|false|false|C0015385|ambulatenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Location|Modifier|false|false||LOCnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Reactive Oxygen Species|Drug|false|false|C0262327|ROS
null|rosiglitazone|Drug|false|false|C0262327|ROS
null|rosiglitazone|Drug|false|false|C0262327|ROS
null|Reactive Oxygen Species|Drug|false|false|C0262327|ROSnull|ROS1 wt Allele|Finding|false|false|C0262327|ROS
null|ROS1 gene|Finding|false|false|C0262327|ROSnull|Review of systems (procedure)|Procedure|false|false|C0262327|ROSnull|rostral sulcus|Anatomy|false|false|C0812281;C1709820;C0289313;C0162772;C0489633|ROSnull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Anemia|Disorder|false|false||Anemianull|Anemia <Anemiaceae>|Entity|false|false||Anemianull|borderline cholesterol|Lab|false|false||Borderline cholesterolnull|Borderline|Modifier|false|false||Borderlinenull|cholesterol|Drug|false|false||cholesterol
null|cholesterol|Drug|false|false||cholesterolnull|Cholesterol measurement|Procedure|false|false||cholesterolnull|Recurrent|Time|false|false||Recurrent
null|Episodic|Time|false|false||Recurrentnull|Flatulence|Finding|false|false||Flatulencenull|Heart murmur|Finding|false|false|C4037974;C0018787|Heart Murmurnull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|Heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|Heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|Heartnull|Chest>Heart|Anatomy|false|false|C0018808;C0795691;C0153957;C0153500;C0018808|Heart
null|Heart|Anatomy|false|false|C0018808;C0795691;C0153957;C0153500;C0018808|Heartnull|Heart murmur|Finding|false|false|C4037974;C0018787|Murmurnull|Hypertensive disease|Disorder|false|false||Hypertensionnull|Hypothyroidism|Disorder|false|false||Hypothyroidismnull|Mitral Valve Insufficiency|Disorder|false|false||Mitral Regurgitationnull|mitral|Modifier|false|false||Mitralnull|Regurgitation|Finding|false|false||Regurgitation
null|Regurgitates after swallowing|Finding|false|false||Regurgitationnull|Regurgitation - mechanism|Phenomenon|false|false||Regurgitationnull|Osteoporosis|Disorder|false|false||Osteoporosisnull|Encounter due to family history of osteoporosis|Finding|false|false||Osteoporosisnull|Pneumonia|Disorder|false|false||Pneumonianull|Sinusitis|Disorder|false|false||Sinusitisnull|Social and personal history|Finding|false|false||Social History
null|Social History|Finding|false|false||Social Historynull|Social|Finding|false|false||Socialnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Family Medical History|Finding|false|false||Family Historynull|Entity Name Part Type - family|Finding|false|false||Family
null|Last Name|Finding|false|false||Family
null|Living Arrangement - Family|Finding|false|false||Family
null|Family (taxonomic)|Finding|false|false||Family
null|Family Collection|Finding|false|false||Familynull|Family|Subject|false|false||Familynull|History of present illness (finding)|Finding|false|true||History
null|History of previous events|Finding|false|true||History
null|Historical aspects qualifier|Finding|false|true||History
null|Medical History|Finding|false|true||History
null|Concept History|Finding|false|true||Historynull|History|Subject|false|false||Historynull|Long Variable|Modifier|false|false||Long
null|Long|Modifier|false|false||Longnull|null|Finding|false|false||history of hypertensionnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Hypertensive disease|Disorder|false|false||hypertensionnull|ErbB Receptors|Drug|false|false||her family
null|ErbB Receptors|Drug|false|false||her familynull|ErbB Receptors|Finding|false|false||her familynull|Entity Name Part Type - family|Finding|false|false||family
null|Last Name|Finding|false|false||family
null|Living Arrangement - Family|Finding|false|false||family
null|Family (taxonomic)|Finding|false|false||family
null|Family Collection|Finding|false|false||familynull|Family|Subject|false|false||familynull|Indirect exposure mechanism - Father|Finding|false|false||Father
null|Relationship - Father|Finding|false|false||Father
null|Father - courtesy title|Finding|false|false||Fathernull|Father (person)|Subject|false|false||Fathernull|Entity Name Part Type - family|Finding|false|false||family
null|Last Name|Finding|false|false||family
null|Living Arrangement - Family|Finding|false|false||family
null|Family (taxonomic)|Finding|false|false||family
null|Family Collection|Finding|false|false||familynull|Family|Subject|false|false||familynull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Numerous|LabModifier|false|false||multiplenull|Malignant Neoplasms|Disorder|false|false||cancersnull|Grandfather|Subject|false|false||grandfathernull|Medical History|Finding|false|false|C3714551;C0038351;C4266636|history ofnull|History of present illness (finding)|Finding|false|false|C3714551;C0038351;C4266636|history
null|History of previous events|Finding|false|false|C3714551;C0038351;C4266636|history
null|Historical aspects qualifier|Finding|false|false|C3714551;C0038351;C4266636|history
null|Medical History|Finding|false|false|C3714551;C0038351;C4266636|history
null|Concept History|Finding|false|false|C3714551;C0038351;C4266636|historynull|History|Subject|false|false||historynull|Malignant neoplasm of stomach|Disorder|false|false|C3714551;C0038351;C4266636|stomach cancer
null|Stomach Carcinoma|Disorder|false|false|C3714551;C0038351;C4266636|stomach cancernull|Neoplasm of uncertain or unknown behavior of stomach|Disorder|false|false|C3714551;C0038351;C4266636|stomach
null|Stomach Diseases|Disorder|false|false|C3714551;C0038351;C4266636|stomach
null|Benign neoplasm of stomach|Disorder|false|false|C3714551;C0038351;C4266636|stomach
null|Carcinoma in situ of stomach|Disorder|false|false|C3714551;C0038351;C4266636|stomachnull|Stomach problem|Finding|false|false|C3714551;C0038351;C4266636|stomachnull|Procedure on stomach|Procedure|false|false|C3714551;C0038351;C4266636|stomachnull|Stomach structure|Anatomy|false|false|C0038354;C0496905;C0153943;C0154060;C0577027;C0024623;C0699791;C0262926;C0006826;C0872393;C0262926;C1705255;C0019665;C0262512;C2004062|stomach
null|Abdomen>Stomach|Anatomy|false|false|C0038354;C0496905;C0153943;C0154060;C0577027;C0024623;C0699791;C0262926;C0006826;C0872393;C0262926;C1705255;C0019665;C0262512;C2004062|stomach
null|Stomach|Anatomy|false|false|C0038354;C0496905;C0153943;C0154060;C0577027;C0024623;C0699791;C0262926;C0006826;C0872393;C0262926;C1705255;C0019665;C0262512;C2004062|stomachnull|Malignant Neoplasms|Disorder|false|false|C3714551;C0038351;C4266636|cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Uncle|Subject|false|false||unclenull|Medical History|Finding|false|true|C0230069;C3665375;C0031354|history ofnull|History of present illness (finding)|Finding|false|false|C0230069;C3665375;C0031354|history
null|History of previous events|Finding|false|false|C0230069;C3665375;C0031354|history
null|Historical aspects qualifier|Finding|false|false|C0230069;C3665375;C0031354|history
null|Medical History|Finding|false|false|C0230069;C3665375;C0031354|history
null|Concept History|Finding|false|false|C0230069;C3665375;C0031354|historynull|History|Subject|false|false||historynull|Throat Homeopathic Medication|Drug|false|true|C0230069;C3665375;C0031354|throatnull|Specimen Type - Throat|Finding|false|true|C0230069;C3665375;C0031354|throat
null|null|Finding|false|true|C0230069;C3665375;C0031354|throatnull|Anterior portion of neck|Anatomy|false|false|C1550663;C1547926;C1950455;C0262926;C1705255;C0019665;C0262512;C2004062;C0262926|throat
null|Throat|Anatomy|false|false|C1550663;C1547926;C1950455;C0262926;C1705255;C0019665;C0262512;C2004062;C0262926|throat
null|Pharyngeal structure|Anatomy|false|false|C1550663;C1547926;C1950455;C0262926;C1705255;C0019665;C0262512;C2004062;C0262926|throatnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Medical History|Finding|true|false||history ofnull|History of present illness (finding)|Finding|true|false||history
null|History of previous events|Finding|true|false||history
null|Historical aspects qualifier|Finding|true|false||history
null|Medical History|Finding|true|false||history
null|Concept History|Finding|true|false||historynull|History|Subject|false|false||historynull|Malignant tumor of colon|Disorder|true|false|C0009368;C4071907|colon cancersnull|Neoplasm of uncertain or unknown behavior of colon|Disorder|true|false|C0009368;C4071907|colon
null|Colonic Diseases|Disorder|true|false|C0009368;C4071907|colon
null|Carcinoma in situ of colon|Disorder|true|false|C0009368;C4071907|colonnull|COLON PROBLEM|Finding|true|false|C0009368;C4071907|colonnull|Colon structure (body structure)|Anatomy|false|false|C0006826;C0007102;C0750873;C0009373;C0154061;C0496907|colon
null|Abdomen+Pelvis>Colon|Anatomy|false|false|C0006826;C0007102;C0750873;C0009373;C0154061;C0496907|colonnull|TUBE,COLON,22FR,RADIOPAQUE RUBBER B#7370|Device|true|false||colonnull|Colon <Coloninae>|Entity|true|false||colonnull|Malignant Neoplasms|Disorder|true|false|C0009368;C4071907|cancersnull|Indirect exposure mechanism - Father|Finding|false|false||Father
null|Relationship - Father|Finding|false|false||Father
null|Father - courtesy title|Finding|false|false||Fathernull|Father (person)|Subject|false|false||Fathernull|Cerebrovascular accident|Disorder|false|false||strokenull|Stroke (heart beat)|Finding|false|false||strokenull|Entity Name Part Type - family|Finding|false|false||family
null|Last Name|Finding|false|false||family
null|Living Arrangement - Family|Finding|false|false||family
null|Family (taxonomic)|Finding|false|false||family
null|Family Collection|Finding|false|false||familynull|Family|Subject|false|false||familynull|Relationship - Mother|Finding|false|false||Mothernull|Mother (person)|Subject|false|false||Mothernull|null|Anatomy|false|false|C0795691;C0153957;C0153500|heart valve
null|Heart Valves|Anatomy|false|false|C0795691;C0153957;C0153500|heart valvenull|Malignant neoplasm of heart|Disorder|false|false|C1186983;C4037974;C0018787;C0018826;C1305961|heart
null|benign neoplasm of heart|Disorder|false|false|C1186983;C4037974;C0018787;C0018826;C1305961|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787;C0018826;C1305961;C1186983|heartnull|Chest>Heart|Anatomy|false|false|C0795691;C0153957;C0153500|heart
null|Heart|Anatomy|false|false|C0795691;C0153957;C0153500|heartnull|Anatomical valve|Anatomy|false|false|C0153957;C0153500;C0795691|valvenull|Valve (physical object)|Device|false|false||valve
null|Valve Device|Device|false|false||valve
null|medical valve|Device|false|false||valvenull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|On admission|Time|false|false||On admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Malignant neoplasm of pelvis|Disorder|false|false|C4266535;C0030797;C0559769|Pelvisnull|Pelvis problem|Finding|false|false|C4266535;C0030797;C0559769|Pelvisnull|Pelvis+|Anatomy|false|false|C0332459;C4551657;C0812455;C0728907;C1547311;C0153663;C1257972;C0565514|Pelvis
null|Pelvic cavity structure|Anatomy|false|false|C0332459;C4551657;C0812455;C0728907;C1547311;C0153663;C1257972;C0565514|Pelvis
null|Pelvis|Anatomy|false|false|C0332459;C4551657;C0812455;C0728907;C1547311;C0153663;C1257972;C0565514|Pelvisnull|Patient Condition Code - Stable|Finding|false|false|C4266535;C0030797;C0559769|stablenull|Stable status|Modifier|false|false||stablenull|Lateral|Modifier|false|false||lateralnull|null|Finding|false|false|C4266535;C0030797;C0559769|compression
null|Compressed structure|Finding|false|false|C4266535;C0030797;C0559769|compressionnull|Compression Therapy|Procedure|false|false|C4266535;C0030797;C0559769|compression
null|Data Compression|Procedure|false|false|C4266535;C0030797;C0559769|compressionnull|Compression|Phenomenon|false|false|C4266535;C0030797;C0559769|compressionnull|Skin clean|Finding|false|false|C1123023;C4520765|skin cleannull|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765|skin
null|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765|skinnull|Skin Specimen Source Code|Finding|false|false|C1123023;C4520765|skin
null|Skin Specimen|Finding|false|false|C1123023;C4520765|skinnull|Skin, Human|Anatomy|false|false|C1947930;C0178298;C0496955;C1554187;C0574729;C1546781;C0444099|skin
null|Skin|Anatomy|false|false|C1947930;C0178298;C0496955;C1554187;C0574729;C1546781;C0444099|skinnull|Cleaning (activity)|Event|false|false|C1123023;C4520765|cleannull|Gender Status - Intact|Finding|false|false|C1123023;C4520765|intactnull|Intact|Modifier|false|false||intactnull|External|Modifier|false|false||externallynull|Rotated|Modifier|false|false||rotatednull|Pain|Finding|false|false||painfulnull|Code System Type - Internal|Modifier|false|false||internal
null|Internal Surface|Modifier|false|false||internal
null|Internal|Modifier|false|false||internalnull|External rotation|Finding|false|false|C1548801;C0022122;C0228391;C0019552;C4299095|external rotationnull|External route|Finding|false|false|C1548801;C0022122;C0228391;C0019552;C4299095|externalnull|Body Site Modifier - External|Anatomy|false|false|C0231462;C0521134;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725|externalnull|Code System Type - External|Modifier|false|false||external
null|External|Modifier|false|false||externalnull|Rotation (malposition) (morphologic abnormality)|Disorder|false|false|C0022122;C0228391;C0019552;C4299095|rotationnull|Musculoskeletal rotation|Finding|false|false|C0022122;C0228391;C0019552;C4299095|rotation
null|null|Finding|false|false|C0022122;C0228391;C0019552;C4299095|rotation
null|Rotation|Finding|false|false|C0022122;C0228391;C0019552;C4299095|rotationnull|heme iron polypeptide|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|ST13 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|ST13 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|RPL29 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|RPL29 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|HHIP protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|HHIP protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|heme iron polypeptide|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hipnull|RPL29 wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C1548801|hip
null|REG3A gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C1548801|hip
null|RPL29 gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C1548801|hip
null|ST13 wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C1548801|hip
null|ST13 gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C1548801|hip
null|HHIP gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C1548801|hip
null|HHIP wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C1548801|hip
null|REG3A wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C1548801|hipnull|Procedure on hip|Procedure|false|false|C0022122;C0228391;C0019552;C4299095|hipnull|Structure of habenulopeduncular tract|Anatomy|false|false|C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C2117331;C0677597;C0035868;C1292890;C1430701;C0529134;C1505163;C1654726;C3669037;C0521134;C0231462|hip
null|Hip structure|Anatomy|false|false|C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C2117331;C0677597;C0035868;C1292890;C1430701;C0529134;C1505163;C1654726;C3669037;C0521134;C0231462|hip
null|Lower extremity>Hip|Anatomy|false|false|C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C2117331;C0677597;C0035868;C1292890;C1430701;C0529134;C1505163;C1654726;C3669037;C0521134;C0231462|hip
null|Bone structure of ischium|Anatomy|false|false|C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C2117331;C0677597;C0035868;C1292890;C1430701;C0529134;C1505163;C1654726;C3669037;C0521134;C0231462|hipnull|Thigh structure|Anatomy|false|false|C3542022|Thighsnull|Leg|Anatomy|false|false||leg
null|Lower Extremity|Anatomy|false|false||legnull|Anatomical compartments|Finding|false|false||compartmentsnull|Compartments [PK]|Phenomenon|false|false||compartmentsnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false|C0039866|softnull|Soft|Modifier|false|false||softnull|sural|Drug|false|false||Suralnull|Deep Resection Margin|Attribute|false|false||Deepnull|Deep (qualifier value)|Modifier|false|false||Deepnull|Peroneal|Modifier|false|false||peronealnull|Superficial|Modifier|false|false||Superficialnull|Peroneal|Modifier|false|false||peronealnull|Feline hyperesthesia syndrome|Disorder|false|false||FHS
null|Fetal hydantoin syndrome|Disorder|false|false||FHSnull|Family Medical History|Finding|false|false||FHSnull|ADGRE4P gene|Finding|false|false||Firenull|Accident caused by unspecified fire|Phenomenon|false|false||Fire
null|Fire as a heat source|Phenomenon|false|false||Fire
null|Fire (physical force)|Phenomenon|false|false||Firenull|fire disaster|Event|false|false||Firenull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Examination of knee joint|Procedure|false|false|C1963703;C0022742;C4299094;C0022745|Kneenull|Knee region structure|Anatomy|false|false|C0042282;C0038435;C0562271;C1547311|Knee
null|Knee|Anatomy|false|false|C0042282;C0038435;C0562271;C1547311|Knee
null|Lower extremity>Knee|Anatomy|false|false|C0042282;C0038435;C0562271;C1547311|Knee
null|Knee joint|Anatomy|false|false|C0042282;C0038435;C0562271;C1547311|Kneenull|Patient Condition Code - Stable|Finding|false|false|C1963703;C0022742;C4299094;C0022745|stablenull|Stable status|Modifier|false|false||stablenull|Varus|Modifier|false|false||varusnull|Valgus deformity|Disorder|false|false|C1963703;C0022742;C4299094;C0022745|valgusnull|Valgus <Valginae>|Entity|false|false||valgusnull|Valgus position|Modifier|false|false||valgusnull|Stress bismuth subsalicylate|Drug|false|false||stress
null|Stress bismuth subsalicylate|Drug|false|false||stressnull|Stress|Finding|false|false|C1963703;C0022742;C4299094;C0022745|stressnull|W stress|Attribute|false|false||stressnull|Rh Negative Blood Group|Finding|false|false||Negative
null|Negative|Finding|false|false||Negative
null|Negative Finding|Finding|false|false||Negativenull|Expression Negative|Lab|false|false||Negativenull|Negative - qualifier|Modifier|false|false||Negative
null|Negative Charge|Modifier|false|false||Negativenull|Negative Number|LabModifier|false|false||Negativenull|Adenohypophyseal Diseases|Disorder|false|false||anteriornull|Anterior|Modifier|false|false||anteriornull|Posterior pituitary disease|Disorder|false|false||posteriornull|Dorsal|Modifier|false|false||posteriornull|Drawers|Device|false|false||drawernull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|On discharge|Time|false|false||On dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|Surgical wound|Disorder|false|false|C2338258|INcisionnull|Surgical incisions|Procedure|false|false|C2338258|INcisionnull|Cranial incision point|Anatomy|false|false|C0184898;C0332803|INcisionnull|Dressing Dosage Form|Drug|false|false||dressingnull|null|Finding|false|false||dressing
null|Ability to dress|Finding|false|false||dressingnull|Dressing patient (procedure)|Procedure|false|false||dressing
null|Dressing of skin or wound|Procedure|false|false||dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Spatial Distribution|Modifier|false|false||distributionsnull|Physiologic pulse|Finding|false|false||pulsenull|Pulse taking|Procedure|false|false||pulsenull|Pulse Rate|Attribute|false|false||pulsenull|Pulse phenomenon|Phenomenon|false|false||pulsenull|heme iron polypeptide|Drug|false|false|C0022122;C0228391;C0019552;C4299095|Hip
null|ST13 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|Hip
null|ST13 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|Hip
null|RPL29 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|Hip
null|RPL29 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|Hip
null|HHIP protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|Hip
null|HHIP protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|Hip
null|heme iron polypeptide|Drug|false|false|C0022122;C0228391;C0019552;C4299095|Hipnull|RPL29 wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095|Hip
null|REG3A gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095|Hip
null|RPL29 gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095|Hip
null|ST13 wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095|Hip
null|ST13 gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095|Hip
null|HHIP gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095|Hip
null|HHIP wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095|Hip
null|REG3A wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095|Hipnull|Procedure on hip|Procedure|false|false|C0022122;C0228391;C0019552;C4299095|Hipnull|Lower extremity>Hip|Anatomy|false|false|C1292890;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1430701;C0529134;C1505163;C1654726|Hip
null|Hip structure|Anatomy|false|false|C1292890;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1430701;C0529134;C1505163;C1654726|Hip
null|Structure of habenulopeduncular tract|Anatomy|false|false|C1292890;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1430701;C0529134;C1505163;C1654726|Hip
null|Bone structure of ischium|Anatomy|false|false|C1292890;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1430701;C0529134;C1505163;C1654726|Hipnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Impacted tooth|Disorder|false|false|C0015811;C0027530;C3159206;C0015815|Impactednull|Impacted|Finding|false|false|C0015815;C0027530;C3159206|Impactednull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Structure of neck of femur|Anatomy|false|false|C0333125;C0812434;C0684335;C0040456|femoral necknull|Femur|Anatomy|false|false|C0040456;C0812434;C0684335|femoralnull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206;C0015815;C0015811|neck
null|Neck problem|Finding|false|false|C0027530;C3159206;C0015815;C0015811|necknull|dendritic spine neck|Anatomy|false|false|C0812434;C0684335;C0040456;C0333125|neck
null|Neck|Anatomy|false|false|C0812434;C0684335;C0040456;C0333125|necknull|Fracture|Disorder|false|false||fracturenull|BRIEF Health Literacy Screening Tool|Finding|false|false||Brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||Briefnull|Brief|Time|false|false||Briefnull|Shortened|Modifier|false|false||Briefnull|Hospital course|Finding|false|false||Hospital Coursenull|null|Attribute|false|false||Hospital Coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||Coursenull|Ortho-|Finding|false|false||orthonull|Ortho Pharmaceutical Ltd|Entity|false|false||orthonull|Physical trauma|Disorder|false|false||trauma
null|Traumatic injury|Disorder|false|false||trauma
null|Trauma|Disorder|false|false||traumanull|Trauma assessment and care|Procedure|false|false||traumanull|Trauma, nursing specialty|Title|false|false||traumanull|trauma qualifier|Modifier|false|false||traumanull|ActInformationPrivacyReason - service|Finding|false|false||servicenull|Software Service|Device|false|false||servicenull|Services|Event|false|false||servicenull|Valgus deformity|Disorder|false|false|C0015815;C0015811;C0833290;C0027530;C3159206|valgusnull|Valgus <Valginae>|Entity|false|false||valgusnull|Valgus position|Modifier|false|false||valgusnull|Neck of left femur|Anatomy|false|false|C0019557;C0149531;C1292890;C0016658;C0042282;C0812434;C0684335;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1552822|left femoral necknull|Table Cell Horizontal Align - left|Finding|false|false|C0015815;C0833290|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Structure of neck of femur|Anatomy|false|false|C0019557;C0149531;C0042282;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1552822;C0016658;C1292890;C0812434;C0684335|femoral necknull|Femur|Anatomy|false|false|C0042282;C0812434;C0684335|femoralnull|Passive joint movement of neck (finding)|Finding|false|false|C0833290;C0027530;C3159206;C0015811;C0015815|neck
null|Neck problem|Finding|false|false|C0833290;C0027530;C3159206;C0015811;C0015815|necknull|dendritic spine neck|Anatomy|false|false|C0019557;C0149531;C0016658;C1292890;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C0812434;C0684335;C0042282|neck
null|Neck|Anatomy|false|false|C0019557;C0149531;C0016658;C1292890;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C0812434;C0684335;C0042282|necknull|Fracture of pelvis|Disorder|false|false|C0833290;C0015815;C0027530;C3159206;C0022122;C0228391;C0019552;C4299095|hip fracture
null|Hip Fractures|Disorder|false|false|C0833290;C0015815;C0027530;C3159206;C0022122;C0228391;C0019552;C4299095|hip fracturenull|heme iron polypeptide|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|ST13 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|ST13 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|RPL29 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|RPL29 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|HHIP protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|HHIP protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|heme iron polypeptide|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hipnull|RPL29 wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C0015815;C0833290;C0027530;C3159206|hip
null|REG3A gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C0015815;C0833290;C0027530;C3159206|hip
null|RPL29 gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C0015815;C0833290;C0027530;C3159206|hip
null|ST13 wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C0015815;C0833290;C0027530;C3159206|hip
null|ST13 gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C0015815;C0833290;C0027530;C3159206|hip
null|HHIP gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C0015815;C0833290;C0027530;C3159206|hip
null|HHIP wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C0015815;C0833290;C0027530;C3159206|hip
null|REG3A wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C0015815;C0833290;C0027530;C3159206|hipnull|Procedure on hip|Procedure|false|false|C0833290;C0022122;C0228391;C0019552;C4299095;C0027530;C3159206;C0015815|hipnull|Lower extremity>Hip|Anatomy|false|false|C1430701;C0529134;C1505163;C1654726;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1292890;C0019557;C0149531;C0016658|hip
null|Hip structure|Anatomy|false|false|C1430701;C0529134;C1505163;C1654726;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1292890;C0019557;C0149531;C0016658|hip
null|Structure of habenulopeduncular tract|Anatomy|false|false|C1430701;C0529134;C1505163;C1654726;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1292890;C0019557;C0149531;C0016658|hip
null|Bone structure of ischium|Anatomy|false|false|C1430701;C0529134;C1505163;C1654726;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1292890;C0019557;C0149531;C0016658|hipnull|Fracture|Disorder|false|false|C0027530;C3159206;C0015815;C0833290;C0022122;C0228391;C0019552;C4299095|fracturenull|Reduced|Finding|false|false||reductionnull|Reduction procedure|Procedure|false|false||reduction
null|Surgical reduction|Procedure|false|false||reductionnull|Reduction (chemical)|Phenomenon|false|false||reductionnull|Percutaneous Route of Drug Administration|Finding|false|false||percutaneousnull|Percutaneous|Modifier|false|false||percutaneousnull|Intramedullary Nailing|Procedure|false|false||pinningnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Femoral Neck Fractures|Disorder|false|false|C0015811;C0027530;C3159206;C0015815|femoral neck fracturenull|Structure of neck of femur|Anatomy|false|false|C0262414;C0812434;C0684335;C0016658;C0015806|femoral necknull|Femur|Anatomy|false|false|C0016658;C0015806;C0812434;C0684335;C0262414|femoralnull|Fracture of cervical spine|Disorder|false|false|C0027530;C3159206;C0015815;C0015811|neck fracturenull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206;C0015811;C0015815|neck
null|Neck problem|Finding|false|false|C0027530;C3159206;C0015811;C0015815|necknull|dendritic spine neck|Anatomy|false|false|C0262414;C0812434;C0684335;C0015806;C0016658|neck
null|Neck|Anatomy|false|false|C0262414;C0812434;C0684335;C0015806;C0016658|necknull|Fracture|Disorder|false|false|C0015811;C0015815;C0027530;C3159206|fracturenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Hypotensive|Finding|false|false||hypotensivenull|Diagnostic Service Section ID - Physical Therapy|Finding|false|false||physical therapynull|Physical therapy|Procedure|false|false||physical therapynull|Physical therapy (field)|Title|false|false||physical therapynull|physical examination (physical finding)|Finding|false|false||physical
null|Physical|Finding|false|false||physicalnull|Physical Examination|Procedure|false|false||physicalnull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|Exercise|Finding|false|false||exercisenull|Exercise Pain Management|Procedure|false|false||exercisenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Diagnostic Service Section ID - Physical Therapy|Finding|false|false||physical therapynull|Physical therapy|Procedure|false|false||physical therapynull|Physical therapy (field)|Title|false|false||physical therapynull|physical examination (physical finding)|Finding|false|false||physical
null|Physical|Finding|false|false||physicalnull|Physical Examination|Procedure|false|false||physicalnull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Rehab facility|Device|false|false||rehab facilitynull|Rehab facility|Entity|false|false||rehab facilitynull|Rehabilitation therapy|Procedure|false|false||rehabnull|ADMIN.FACILITY|Finding|false|false||facilitynull|Facility (object)|Device|false|false||facilitynull|Social Work (discipline)|Subject|false|false||SOcial worknull|Social|Finding|false|false||SOcialnull|Work|Event|false|false||worknull|Difficulty coping|Finding|false|false||difficulty copingnull|Has difficulty doing (qualifier value)|Finding|false|false||difficultynull|Child coping with hospitalization|Finding|false|false||coping
null|Coping Behavior|Finding|false|false||copingnull|COPING - Dental Restorative Procedure|Procedure|false|false||coping
null|COPING - Fixed Prosthodontics|Procedure|false|false||copingnull|Decreasing|Finding|false|false||decreased
null|Reduced|Finding|false|false||decreasednull|Decreased|LabModifier|false|false||decreasednull|Mobility finding|Finding|false|false||mobilitynull|Range of Motion, Articular|Attribute|false|false||mobilitynull|Mobility (attribute)|Modifier|false|false||mobilitynull|Laboratory test finding|Lab|false|false||labsnull|Sodium measurement|Procedure|false|false||sodium levelnull|Finding of sodium level|Lab|false|false||sodium levelnull|Sodium supplements|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|Sodium Drug Class|Drug|false|false||sodiumnull|Sodium metabolic function|Finding|false|false||sodiumnull|Sodium measurement|Procedure|false|false||sodiumnull|null|Finding|false|false||unchangednull|About The Same|Modifier|false|false||unchangednull|Similarity|Modifier|false|false||similarnull|On admission|Time|false|false||on admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Instructions|Finding|false|false||instructions
null|Instruction [Publication Type]|Finding|false|false||instructionsnull|null|Attribute|false|false||instructionsnull|Clinic|Device|false|false||clinic
null|Ambulatory Care Facilities|Device|false|false||clinicnull|Clinic|Entity|false|false||clinic
null|Ambulatory Care Facilities|Entity|false|false||clinicnull|Patient location type - Clinic|Modifier|false|false||clinic
null|Person location type - Clinic|Modifier|false|false||clinicnull|2 Weeks|Time|false|false||2 weeksnull|week|Time|false|false||weeksnull|Lovenox|Drug|false|false||lovenox
null|Lovenox|Drug|false|false||lovenoxnull|Daily|Time|false|false||dailynull|Interim|Time|false|false||interimnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Accurate (qualifier value)|Modifier|false|false||accuratenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|levothyroxine sodium|Drug|false|false||Levothyroxine Sodium
null|levothyroxine sodium|Drug|false|false||Levothyroxine Sodium
null|levothyroxine sodium|Drug|false|false||Levothyroxine Sodiumnull|Synthetic Levothyroxine|Drug|false|false||Levothyroxine
null|Synthetic Levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxinenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|microgram|LabModifier|false|false||mcgnull|Daily|Time|false|false||DAILYnull|lisinopril|Drug|false|false||Lisinopril
null|lisinopril|Drug|false|false||Lisinoprilnull|Daily|Time|false|false||DAILYnull|methylphenidate|Drug|false|false||MethylPHENIDATE
null|methylphenidate|Drug|false|false||MethylPHENIDATEnull|Poisoning by, adverse effect of and underdosing of methylphenidate|Disorder|false|false||MethylPHENIDATEnull|Methylphenidate measurement|Procedure|false|false||MethylPHENIDATEnull|Ritalin|Drug|false|false||Ritalin
null|Ritalin|Drug|false|false||Ritalinnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|mirtazapine|Drug|false|false||mirtazapine
null|mirtazapine|Drug|false|false||mirtazapinenull|Oral Dosage Form|Drug|false|false|C0226896|Oralnull|Oral Route of Administration|Finding|false|false|C0226896|Oral
null|Oral (intended site)|Finding|false|false|C0226896|Oralnull|Oral cavity|Anatomy|false|false|C1527415;C4521986;C1272919|Oralnull|Oral|Modifier|false|false||Oralnull|Once a day, at bedtime|Time|false|false||QHSnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|levothyroxine sodium|Drug|false|false||Levothyroxine Sodium
null|levothyroxine sodium|Drug|false|false||Levothyroxine Sodium
null|levothyroxine sodium|Drug|false|false||Levothyroxine Sodiumnull|Synthetic Levothyroxine|Drug|false|false||Levothyroxine
null|Synthetic Levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxinenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|microgram|LabModifier|false|false||mcgnull|Daily|Time|false|false||DAILYnull|lisinopril|Drug|false|false||Lisinopril
null|lisinopril|Drug|false|false||Lisinoprilnull|Daily|Time|false|false||DAILYnull|methylphenidate|Drug|false|false||MethylPHENIDATE
null|methylphenidate|Drug|false|false||MethylPHENIDATEnull|Poisoning by, adverse effect of and underdosing of methylphenidate|Disorder|false|false||MethylPHENIDATEnull|Methylphenidate measurement|Procedure|false|false||MethylPHENIDATEnull|Ritalin|Drug|false|false||Ritalin
null|Ritalin|Drug|false|false||Ritalinnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|mirtazapine|Drug|false|false||mirtazapine
null|mirtazapine|Drug|false|false||mirtazapinenull|Oral Dosage Form|Drug|false|false|C0226896|Oralnull|Oral Route of Administration|Finding|false|false|C0226896|Oral
null|Oral (intended site)|Finding|false|false|C0226896|Oralnull|Oral cavity|Anatomy|false|false|C1527415;C4521986;C1272919|Oralnull|Oral|Modifier|false|false||Oralnull|Once a day, at bedtime|Time|false|false||QHSnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|aluminum|Drug|false|false||Aluminum
null|aluminum|Drug|false|false||Aluminumnull|Aluminum measurement|Procedure|false|false||Aluminumnull|Magnesium supplements, alimentary tract and metabolism|Drug|false|false||Magnesium
null|magnesium|Drug|false|false||Magnesium
null|magnesium|Drug|false|false||Magnesium
null|Magnesium Drug Class|Drug|false|false||Magnesium
null|Magnesium supplements, alimentary tract and metabolism|Drug|false|false||Magnesiumnull|Magnesium measurement|Procedure|false|false||Magnesiumnull|simethicone|Drug|false|false||Simethicone
null|simethicone|Drug|false|false||Simethiconenull|Four times daily|Time|false|false||QIDnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Dyspepsia|Finding|false|false||Dyspepsianull|artificial tears (medication)|Drug|false|false||Artificial Tears
null|Lubricant Eye Drops|Drug|false|false||Artificial Tears
null|Artificial Tears|Drug|false|false||Artificial Tearsnull|Artificial (qualifier value)|Modifier|false|false||Artificialnull|Tears (substance)|Finding|false|false||Tears
null|null|Finding|false|false||Tears
null|Tears specimen|Finding|false|false||Tearsnull|Drops - Drug Form|Drug|false|false||DROPnull|Dropping|Event|false|false||DROPnull|Drop (unit of presentation)|LabModifier|false|false||DROP
null|Drop British|LabModifier|false|false||DROP
null|Drop Dosing Unit|LabModifier|false|false||DROP
null|Medical Drop|LabModifier|false|false||DROP
null|Drop Unit of Volume|LabModifier|false|false||DROPnull|Structure of both eyes|Anatomy|false|false|C1422467|BOTH EYESnull|Eye|Anatomy|false|false|C5848506;C1422467|EYESnull|null|Attribute|false|false|C0015392|EYESnull|CIAO3 gene|Finding|false|false|C0229118;C0015392|PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Dry Eyes brand of ocular lubricant|Drug|false|false|C0015392|dry eyesnull|Dry Eye Syndromes|Disorder|false|false|C0015392|dry eyes
null|Keratoconjunctivitis Sicca|Disorder|false|false|C0015392|dry eyesnull|Dryness of eye|Finding|false|false|C0015392|dry eyesnull|Eye|Anatomy|false|false|C5848506;C0720056;C0314719;C0022575;C0013238|eyesnull|null|Attribute|false|false|C0015392|eyesnull|Biotene Dry Mouth|Drug|false|false|C0230028;C0226896|Biotene Dry Mouthnull|Biotene|Drug|false|false||Biotene
null|Biotene|Drug|false|false||Biotene
null|Biotene|Drug|false|false||Biotenenull|Xerostomia|Disorder|false|false|C0230028;C0226896|Dry Mouthnull|Mouthwash|Drug|false|false|C0230028;C0226896|Mouth Rinsenull|Mouth Rinse Specimen|Finding|false|false|C0230028;C0226896|Mouth Rinsenull|Oral cavity|Anatomy|false|false|C5849077;C0026647;C0043352;C0036087;C0438730;C1546769;C5762022|Mouth
null|Oral region|Anatomy|false|false|C5849077;C0026647;C0043352;C0036087;C0438730;C1546769;C5762022|Mouthnull|Rinse Dosage Form|Finding|false|false||Rinsenull|Rinsing|Event|false|false||Rinsenull|Saliva specimen|Finding|false|false|C0230028;C0226896|saliva
null|null|Finding|false|false|C0230028;C0226896|saliva
null|saliva|Finding|false|false|C0230028;C0226896|salivanull|Substitution - ActClass|Finding|false|false||substitutionnull|Substitution - change|Event|false|false||substitutionnull|HL7 Version 2.5 - Application|Finding|false|false|C0026724|application
null|Application Document|Finding|false|false|C0026724|application
null|Computer Application|Finding|false|false|C0026724|application
null|Regulatory Application|Finding|false|false|C0026724|application
null|Apply|Finding|false|false|C0026724|applicationnull|Application procedure|Procedure|false|false|C0026724|applicationnull|Application - unit of product usage|LabModifier|false|false||applicationnull|Disease of mucous membrane|Disorder|false|false|C0026724;C0596901;C0025255|Mucous Membranenull|Route of Administration - Mucous Membrane|Finding|false|false|C0596901;C0025255;C0026724|Mucous Membranenull|Mucous Membrane|Anatomy|false|false|C0185125;C0151785;C0870325;C4048755;C2347934;C1947919;C1547755;C1549524;C2753459;C0026727|Mucous Membranenull|Mucus (substance)|Finding|false|false|C0026724|Mucous
null|mucus layer|Finding|false|false|C0026724|Mucousnull|Mucous appearance|Modifier|false|false||Mucousnull|Membrane Tissue|Anatomy|false|false|C1549524;C0151785|Membrane
null|Membrane|Anatomy|false|false|C1549524;C0151785|Membranenull|Membrane Device|Device|false|false||Membranenull|bisacodyl|Drug|false|false||Bisacodyl
null|bisacodyl|Drug|false|false||Bisacodylnull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Constipation|Finding|false|false||Constipationnull|calcium carbonate|Drug|false|false||Calcium Carbonate
null|calcium carbonate|Drug|false|false||Calcium Carbonatenull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|carbonate ion|Drug|false|false||Carbonate
null|Carbonates|Drug|false|false||Carbonate
null|Carbonates|Drug|false|false||Carbonatenull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|enoxaparin sodium|Drug|false|false||Enoxaparin Sodium
null|enoxaparin sodium|Drug|false|false||Enoxaparin Sodiumnull|enoxaparin|Drug|false|false||Enoxaparin
null|enoxaparin|Drug|false|false||Enoxaparinnull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false|C5239664|Sodiumnull|Daily|Time|false|false||DAILYnull|DVT prophylaxis|Procedure|false|false|C5239664|DVT prophylaxisnull|Deep thrombophlebitis|Disorder|false|false|C5239664|DVT
null|Deep Vein Thrombosis|Disorder|false|false|C5239664|DVTnull|area DVT|Anatomy|false|false|C2926618;C0149871;C0151950;C0337443;C0853245;C0199176|DVTnull|null|Attribute|false|false|C5239664|DVTnull|Prophylactic treatment|Procedure|false|false|C5239664|prophylaxisnull|prevention & control|Modifier|false|false||prophylaxisnull|Duration brand of oxymetazoline|Drug|false|false||Durationnull|Duration (temporal concept)|Time|false|false||Durationnull|14 days|Time|false|false||14 Daysnull|day|Time|false|false||Daysnull|Firstly|Modifier|false|false||Firstnull|First (number)|LabModifier|false|false||Firstnull|Unit dose|LabModifier|false|false||Dose
null|Dosage|LabModifier|false|false||Dosenull|next - HtmlLinkType|Finding|false|false||Nextnull|Following|Time|false|false||Next
null|Then|Time|false|false||Nextnull|Adjacent|Modifier|false|false||Nextnull|Extended Priority Codes - Routine|Finding|false|false||Routine
null|Report priority - Routine|Finding|false|false||Routine
null|Admission Type - Routine|Finding|false|false||Routine
null|Level of Care - Routine|Finding|false|false||Routine
null|Processing priority - Routine|Finding|false|false||Routine
null|Referral priority - Routine|Finding|false|false||Routinenull|Routine coag|Procedure|false|false||Routinenull|Priority - Routine|Time|false|false||Routinenull|Routine|Modifier|false|false||Routinenull|Administration (procedure)|Procedure|false|false||Administrationnull|Administration occupational activities|Event|false|false||Administrationnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||Time
null|Time (foundation metadata concept)|Finding|false|false||Time
null|Value type - Time|Finding|false|false||Time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||Time
null|Data types - Time|Finding|false|false||Time
null|null|Finding|false|false||Timenull|Time|Time|false|false||Timenull|enoxaparin|Drug|false|false||enoxaparin
null|enoxaparin|Drug|false|false||enoxaparinnull|Daily|Time|false|false||dailynull|Syringes|Device|false|false||Syringenull|Syringe (unit of presentation)|LabModifier|false|false||Syringe
null|Syringe Dosing Unit|LabModifier|false|false||Syringenull|refill|Finding|false|false||Refillsnull|Milk of Magnesia (Brand Name)|Drug|false|false||Milk of Magnesia
null|Milk of Magnesia (Brand Name)|Drug|false|false||Milk of Magnesia
null|magnesium hydroxide Oral Suspension|Drug|false|false||Milk of Magnesianull|cow milk allergenic extract|Drug|false|false||Milk
null|Milk antigen|Drug|false|false||Milk
null|Milk Beverage|Drug|false|false||Milk
null|Plant-Based Milk|Drug|false|false||Milk
null|cow milk allergenic extract|Drug|false|false||Milk
null|Milk Specimen|Drug|false|false||Milk
null|Cow's milk|Drug|false|false||Milk
null|null|Drug|false|false||Milknull|Milk (body substance)|Finding|false|false||Milk
null|Milk Specimen Code|Finding|false|false||Milknull|magnesium oxide|Drug|false|false||Magnesia
null|magnesium oxide|Drug|false|false||Magnesianull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Dyspepsia|Finding|false|false||Dyspepsianull|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitaminsnull|capsule (pharmacologic)|Drug|false|false||CAPnull|CATARACT, ANTERIOR POLAR|Disorder|false|false||CAPnull|BRD4 wt Allele|Finding|false|false||CAP
null|HACD1 gene|Finding|false|false||CAP
null|SERPINB6 gene|Finding|false|false||CAP
null|BRD4 gene|Finding|false|false||CAP
null|CAP1 gene|Finding|false|false||CAP
null|SORBS1 gene|Finding|false|false||CAP
null|LNPEP gene|Finding|false|false||CAPnull|CAP Regimen|Procedure|false|false||CAP
null|cisplatin/cyclophosphamide/doxorubicin protocol|Procedure|false|false||CAP
null|cyclophosphamide/doxorubicin/prednisone protocol|Procedure|false|false||CAPnull|Cap (physical object)|Device|false|false||CAP
null|Syringe Caps|Device|false|false||CAP
null|Cap device|Device|false|false||CAPnull|College of American Pathologists|Subject|false|false||CAPnull|Controlled Attenuation Parameter|Modifier|false|false||CAPnull|Capsule Dosing Unit|LabModifier|false|false||CAPnull|Daily|Time|false|false||DAILYnull|oxycodone|Drug|false|false||OxycoDONE
null|oxycodone|Drug|false|false||OxycoDONEnull|Oxycodone measurement|Procedure|false|false||OxycoDONEnull|Immediate Release Dosage Form|Drug|false|false||Immediate Releasenull|Query Priority - Immediate|Finding|false|false||Immediate
null|immediate - ResponseCode|Finding|false|false||Immediatenull|Immediate|Time|false|false||Immediate
null|Stat (do immediately)|Time|false|false||Immediatenull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|oxycodone|Drug|false|false||oxycodone
null|oxycodone|Drug|false|false||oxycodonenull|Oxycodone measurement|Procedure|false|false||oxycodonenull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1527415|mouth
null|Oral region|Anatomy|false|false|C1527415|mouthnull|Hour|Time|false|false||hoursnull|PRSS30P gene|Finding|false|false||Dispnull|Dispense (activity)|Event|false|false||Dispnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|pantoprazole|Drug|false|false||Pantoprazole
null|pantoprazole|Drug|false|false||Pantoprazolenull|Every twenty four hours|Time|false|false||Q24Hnull|sennosides, USP|Drug|false|false||Senna
null|sennosides, USP|Drug|false|false||Sennanull|Senna alexandrina|Entity|false|false||Senna
null|Senna Plant|Entity|false|false||Sennanull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|Storage Unit|Device|false|false||UNIT
null|Unit device|Device|false|false||UNITnull|Unit - NCI Thesaurus Property|LabModifier|false|false||UNIT
null|Unit of Measure|LabModifier|false|false||UNIT
null|Unit|LabModifier|false|false||UNIT
null|Enzyme Unit|LabModifier|false|false||UNITnull|Daily|Time|false|false||DAILYnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|long-term care|Procedure|false|false||Extended Carenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Neck of left femur|Anatomy|false|false|C0262414;C0812434;C0684335;C0016658;C1552822;C0015806|left femoral necknull|Table Cell Horizontal Align - left|Finding|false|false|C0015815;C0833290|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Femoral Neck Fractures|Disorder|false|false|C0015811;C0027530;C3159206;C0015815;C0833290|femoral neck fracturenull|Structure of neck of femur|Anatomy|false|false|C1552822;C0015806;C0262414;C0016658;C0812434;C0684335|femoral necknull|Femur|Anatomy|false|false|C0015806;C0812434;C0684335;C0262414|femoralnull|Fracture of cervical spine|Disorder|false|false|C0833290;C0027530;C3159206;C0015811;C0015815|neck fracturenull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206;C0833290;C0015811;C0015815|neck
null|Neck problem|Finding|false|false|C0027530;C3159206;C0833290;C0015811;C0015815|necknull|dendritic spine neck|Anatomy|false|false|C0015806;C0016658;C0262414;C0812434;C0684335|neck
null|Neck|Anatomy|false|false|C0015806;C0016658;C0262414;C0812434;C0684335|necknull|Fracture|Disorder|false|false|C0027530;C3159206;C0833290;C0015815|fracturenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Disease|Disorder|false|false||Conditionnull|Logical Condition|Finding|false|false||Conditionnull|null|Attribute|false|false||Conditionnull|Condition|Modifier|false|false||Conditionnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|BORNHOLM EYE DISEASE|Disorder|false|false||Bednull|Bachelor of Education|Finding|false|false||Bednull|Beds|Device|false|false||Bednull|Patient Location - Bed|Modifier|false|false||Bednull|Helping Behavior|Finding|false|false||assistancenull|Assisted (qualifier value)|Modifier|false|false||assistancenull|Chairs|Device|false|false||chairnull|Chairperson|Subject|false|false||chairnull|has wheelchair at home (history)|Finding|false|false||wheelchair
null|Wheelchair Usually Used|Finding|false|false||wheelchairnull|wheelchair|Device|false|false||wheelchairnull|Discharge instructions|Finding|false|false||Discharge Instructionsnull|hospital discharge instructions (treatment)|Procedure|false|false||Discharge Instructionsnull|null|Attribute|false|false||Discharge Instructionsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|Pharmaceutical Preparations|Drug|false|false||MEDICATIONSnull|Medications|Finding|false|false||MEDICATIONSnull|null|Attribute|false|false||MEDICATIONS
null|null|Attribute|false|false||MEDICATIONSnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Physicians|Subject|false|false||physiciansnull|At discharge|Time|false|false||at dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|null|Attribute|false|false||surgeonnull|Surgeon|Subject|false|false||surgeonnull|Alcohols|Drug|false|false||alcohol
null|Alcohols|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcoholnull|Alcohol - Recreational Drug Use Code|Finding|false|false||alcoholnull|Motor Vehicles|Device|false|false||motor vehiclenull|motor movement|Finding|false|false||motornull|Motor Device|Device|false|false||motornull|Drug vehicle|Drug|false|false||vehiclenull|Vehicle (transportation)|Device|false|false||vehiclenull|operate|Finding|false|false||operatenull|Contact with machinery|Disorder|false|false||machinerynull|Industrial machine|Device|false|false||machinerynull|Narcotics|Drug|false|false||narcotic
null|Narcotics|Drug|false|false||narcoticnull|Pain Relieve brand of acetaminophen|Drug|false|false||pain relievers
null|Pain Relieve brand of acetaminophen|Drug|false|false||pain relievers
null|Analgesics|Drug|false|false||pain relievers
null|Analgesics|Drug|false|false||pain relievers
null|Analgesics|Drug|false|false||pain relieversnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Narcotics|Drug|false|false||Narcotic
null|Narcotics|Drug|false|false||Narcoticnull|Pain Relieve brand of acetaminophen|Drug|false|false||pain relievers
null|Pain Relieve brand of acetaminophen|Drug|false|false||pain relievers
null|Analgesics|Drug|false|false||pain relievers
null|Analgesics|Drug|false|false||pain relievers
null|Analgesics|Drug|false|false||pain relieversnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Constipation|Finding|false|false||constipationnull|Drink (dietary substance)|Drug|false|false||drinknull|Eyeglasses|Device|false|false||glassesnull|Water Specimen|Drug|false|false||water
null|water|Drug|false|false||water
null|water|Drug|false|false||waternull|Water - Specimen Source Codes|Finding|false|false||waternull|Hydrotherapy|Procedure|false|false||waternull|Daily|Time|false|false||dailynull|Stool Softener brand of docusate sodium|Drug|false|false||stool softener
null|Stool Softener brand of docusate sodium|Drug|false|false||stool softener
null|Stool Softener|Drug|false|false||stool softenernull|Feces|Finding|false|false||stoolnull|Stool seat|Device|false|false||stoolnull|Colace|Drug|false|false||colace
null|Colace|Drug|false|false||colacenull|Adverse effects|Finding|false|false||side effectnull|Side|Modifier|false|false||sidenull|Effect, Appearance|Modifier|false|false||effect
null|Effect|Modifier|false|false||effectnull|ANTICOAGULATION (finding)|Finding|false|false||ANTICOAGULATION
null|Anticoagulation function|Finding|false|false||ANTICOAGULATION
null|Decreased Coagulation Activity [PE]|Finding|false|false||ANTICOAGULATIONnull|Anticoagulation Therapy|Procedure|false|false||ANTICOAGULATIONnull|Lovenox|Drug|false|false||lovenox
null|Lovenox|Drug|false|false||lovenoxnull|Daily|Time|false|false||dailynull|2 Weeks|Time|false|false||2 weeksnull|week|Time|false|false||weeksnull|Wound care management|Procedure|false|false||WOUND CARE
null|wound care|Procedure|false|false||WOUND CAREnull|Wound Care kit|Device|false|false||WOUND CAREnull|Traumatic Wound|Disorder|false|false||WOUND
null|Wounds and Injuries|Disorder|false|false||WOUND
null|Traumatic injury|Disorder|false|false||WOUNDnull|Route of Administration - Wound|Finding|false|false||WOUND
null|null|Finding|false|false||WOUND
null|Specimen Type - Wound|Finding|false|false||WOUNDnull|In care (finding)|Finding|false|false||CARE
null|Continuity Assessment Record and Evaluation|Finding|false|false||CAREnull|care activity|Event|false|false||CAREnull|Traumatic Wound|Disorder|false|false||wound
null|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|Moist|Modifier|false|false||wetnull|take a shower|Finding|false|false||take a showernull|Shower (physical object)|Device|false|false||showernull|3 Days|Time|false|false||3 daysnull|day|Time|false|false||daysnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Gently|Modifier|false|false||gentlynull|Soap Dosage Form|Drug|false|false||soapnull|Soap|Device|false|false||soapnull|Water Specimen|Drug|false|false||water
null|water|Drug|false|false||water
null|water|Drug|false|false||waternull|Water - Specimen Source Codes|Finding|false|false||waternull|Hydrotherapy|Procedure|false|false||waternull|Fenamole|Drug|false|false||pat
null|Fenamole|Drug|false|false||patnull|Paroxysmal atrial tachycardia|Disorder|false|false||patnull|glutamate-prephenate aminotransferase activity|Finding|false|false||pat
null|aspartate-prephenate aminotransferase activity|Finding|false|false||pat
null|protein acetyltransferase activity|Finding|false|false||patnull|Thermoacoustic Computed Tomography|Procedure|false|false||patnull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0184898;C0332803|incisionnull|Bathing|Procedure|true|false||bathsnull|Baths (medical device)|Device|true|false||bathsnull|swimming (history)|Finding|true|false||swimming
null|Swimming|Finding|true|false||swimmingnull|4 Weeks|Time|false|false||4 weeksnull|week|Time|false|false||weeksnull|Staple, Surgical|Device|false|false||staplesnull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Appointments|Event|false|false||appointmentnull|Dressing Dosage Form|Drug|true|false||dressingnull|Ability to dress|Finding|true|false||dressing
null|null|Finding|true|false||dressingnull|Dressing of skin or wound|Procedure|true|false||dressing
null|Dressing patient (procedure)|Procedure|true|false||dressingnull|Wound Dressings (device)|Device|true|false||dressing
null|Dress (garment)|Device|true|false||dressing
null|Medical dressing|Device|true|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Traumatic Wound|Disorder|false|false||wound
null|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|Activity (animal life circumstance)|Finding|false|false||ACTIVITY
null|Physical activity|Finding|false|false||ACTIVITYnull|Activities|Event|false|false||ACTIVITYnull|null|Modifier|false|false||ACTIVITYnull|Weight-Bearing state|Subject|false|false||WEIGHT BEARINGnull|infant weight for previous delivery (history)|Finding|false|false||WEIGHT
null|Weight symptom (finding)|Finding|false|false||WEIGHTnull|Weighing patient|Procedure|false|false||WEIGHTnull|null|Attribute|false|false||WEIGHTnull|Body Weight|Subject|false|false||WEIGHTnull|Importance Weight|Modifier|false|false||WEIGHTnull|Weight|LabModifier|false|false||WEIGHTnull|Bearing Device|Device|false|false||BEARINGnull|Touch Perception|Finding|false|false||touch
null|Touch sensation|Finding|false|false||touchnull|Therapeutic Touch|Procedure|false|false||touchnull|Tactile|Modifier|false|false||touchnull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|Diagnostic Service Section ID - Physical Therapy|Finding|false|false||Physical Therapynull|Physical therapy|Procedure|false|false||Physical Therapynull|Physical therapy (field)|Title|false|false||Physical Therapynull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Therapy Object (animal model)|Finding|false|false||Therapy
null|therapeutic aspects|Finding|false|false||Therapynull|Therapeutic procedure|Procedure|false|false||Therapynull|Touch Perception|Finding|false|false||Touch
null|Touch sensation|Finding|false|false||Touchnull|Therapeutic Touch|Procedure|false|false||Touchnull|Tactile|Modifier|false|false||Touchnull|Weight-Bearing state|Subject|false|false||weight bearingnull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|Bearing Device|Device|false|false||bearingnull|Therapeutic procedure|Procedure|false|false||Treatmentsnull|Frequency|Finding|false|false||Frequency
null|How Often|Finding|false|false||Frequencynull|With frequency|Time|false|false||Frequency
null|Frequencies (time pattern)|Time|false|false||Frequencynull|Kind of quantity - Frequency|LabModifier|false|false||Frequency
null|Statistical Frequency|LabModifier|false|false||Frequency
null|Spatial Frequency|LabModifier|false|false||Frequencynull|Wound care management|Procedure|false|false||WOUND CARE
null|wound care|Procedure|false|false||WOUND CAREnull|Wound Care kit|Device|false|false||WOUND CAREnull|Traumatic Wound|Disorder|false|false||WOUND
null|Wounds and Injuries|Disorder|false|false||WOUND
null|Traumatic injury|Disorder|false|false||WOUNDnull|Route of Administration - Wound|Finding|false|false||WOUND
null|null|Finding|false|false||WOUND
null|Specimen Type - Wound|Finding|false|false||WOUNDnull|In care (finding)|Finding|false|false||CARE
null|Continuity Assessment Record and Evaluation|Finding|false|false||CAREnull|care activity|Event|false|false||CAREnull|Traumatic Wound|Disorder|false|false||wound
null|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|Moist|Modifier|false|false||wetnull|take a shower|Finding|false|false||take a showernull|Shower (physical object)|Device|false|false||showernull|3 Days|Time|false|false||3 daysnull|day|Time|false|false||daysnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Gently|Modifier|false|false||gentlynull|Soap Dosage Form|Drug|false|false||soapnull|Soap|Device|false|false||soapnull|Water Specimen|Drug|false|false||water
null|water|Drug|false|false||water
null|water|Drug|false|false||waternull|Water - Specimen Source Codes|Finding|false|false||waternull|Hydrotherapy|Procedure|false|false||waternull|Fenamole|Drug|false|false||pat
null|Fenamole|Drug|false|false||patnull|Paroxysmal atrial tachycardia|Disorder|false|false||patnull|glutamate-prephenate aminotransferase activity|Finding|false|false||pat
null|aspartate-prephenate aminotransferase activity|Finding|false|false||pat
null|protein acetyltransferase activity|Finding|false|false||patnull|Thermoacoustic Computed Tomography|Procedure|false|false||patnull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0332803;C0184898|incisionnull|Bathing|Procedure|true|false||bathsnull|Baths (medical device)|Device|true|false||bathsnull|swimming (history)|Finding|true|false||swimming
null|Swimming|Finding|true|false||swimmingnull|4 Weeks|Time|false|false||4 weeksnull|week|Time|false|false||weeksnull|Staple, Surgical|Device|false|false||staplesnull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Appointments|Event|false|false||appointmentnull|Dressing Dosage Form|Drug|true|false||dressingnull|Ability to dress|Finding|true|false||dressing
null|null|Finding|true|false||dressingnull|Dressing of skin or wound|Procedure|true|false||dressing
null|Dressing patient (procedure)|Procedure|true|false||dressingnull|Wound Dressings (device)|Device|true|false||dressing
null|Dress (garment)|Device|true|false||dressing
null|Medical dressing|Device|true|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Traumatic Wound|Disorder|false|false||wound
null|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions