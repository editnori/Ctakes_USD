 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|49,58|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|49,58|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|49,63|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|83,92|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|83,92|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|83,92|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|83,92|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|83,92|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|83,97|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|115,120|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|115,120|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|115,120|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|139,142|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|139,142|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|139,142|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|139,142|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|139,142|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|150,157|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|150,157|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|159,167|true|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|Allergies|191,200|true|false|false|C1717415||Allergies
Event|Event|Allergies|191,200|true|false|false|||Allergies
Finding|Pathologic Function|Allergies|191,200|true|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|Allergies|203,225|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|Allergies|211,215|true|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|Allergies|211,215|true|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|Allergies|211,225|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Event|Event|Allergies|216,225|true|false|false|||Reactions
Event|Event|Allergies|228,237|false|false|false|||Attending
Finding|Functional Concept|Allergies|228,237|false|false|false|C1999232|Attending (action)|Attending
Finding|Functional Concept|Chief Complaint|263,269|false|false|false|C0234621|Visual|Visual
Finding|Sign or Symptom|Chief Complaint|263,284|false|false|false|C0233763|Hallucinations, Visual|Visual hallucinations
Disorder|Mental or Behavioral Dysfunction|Chief Complaint|270,284|false|false|false|C0018524|Hallucinations|hallucinations
Event|Event|Chief Complaint|270,284|false|false|false|||hallucinations
Finding|Classification|Chief Complaint|287,292|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|293,301|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|293,301|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|305,323|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|314,323|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|314,323|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|314,323|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|314,323|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|314,323|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|Chief Complaint|325,326|false|false|false|||N
Finding|Finding|History of Present Illness|364,368|false|false|false|C1706180|Male Gender|male
Disorder|Disease or Syndrome|History of Present Illness|378,385|false|false|false|C0012634|Disease|disease
Event|Event|History of Present Illness|378,385|false|false|false|||disease
Disorder|Disease or Syndrome|History of Present Illness|387,399|false|false|false|C0242339|Dyslipidemias|dyslipidemia
Event|Event|History of Present Illness|387,399|false|false|false|||dyslipidemia
Event|Event|History of Present Illness|407,414|false|false|false|||history
Finding|Conceptual Entity|History of Present Illness|407,414|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|407,414|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|407,414|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|407,417|false|false|false|C0262926|Medical History|history of
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|418,426|false|false|false|C0033572;C4266527|Prostate;Structure of prostate (body structure)|prostate
Disorder|Disease or Syndrome|History of Present Illness|418,426|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|prostate
Disorder|Neoplastic Process|History of Present Illness|418,426|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|prostate
Disorder|Neoplastic Process|History of Present Illness|418,433|false|false|false|C0376358;C0600139|Malignant neoplasm of prostate;Prostate carcinoma|prostate cancer
Disorder|Neoplastic Process|History of Present Illness|427,433|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|History of Present Illness|427,433|false|false|false|||cancer
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|439,452|false|false|false|C0033573|Prostatectomy|prostatectomy
Event|Event|History of Present Illness|462,470|false|false|false|||referred
Event|Event|History of Present Illness|514,518|false|false|false|||gait
Finding|Finding|History of Present Illness|514,518|false|false|false|C0016928|Gait|gait
Disorder|Injury or Poisoning|History of Present Illness|520,525|false|false|false|C0000921|Accidental Falls|falls
Event|Event|History of Present Illness|520,525|false|false|false|||falls
Finding|Finding|History of Present Illness|520,525|false|false|false|C0085639|Falls|falls
Finding|Functional Concept|History of Present Illness|531,537|false|false|false|C0234621|Visual|visual
Finding|Sign or Symptom|History of Present Illness|531,552|false|false|false|C0233763|Hallucinations, Visual|visual hallucinations
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|538,552|false|false|false|C0018524|Hallucinations|hallucinations
Event|Event|History of Present Illness|538,552|false|false|false|||hallucinations
Event|Event|History of Present Illness|570,577|false|false|false|||history
Finding|Conceptual Entity|History of Present Illness|570,577|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|570,577|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|570,577|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Event|Event|History of Present Illness|581,586|false|false|false|||taken
Finding|Intellectual Product|History of Present Illness|592,597|false|false|false|C0684240|Charts (publication)|chart
Procedure|Health Care Activity|History of Present Illness|592,604|false|false|false|C0541653|Chart evaluation by healthcare professional|chart review
Event|Event|History of Present Illness|598,604|false|false|false|||review
Finding|Idea or Concept|History of Present Illness|598,604|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Intellectual Product|History of Present Illness|598,604|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Body Substance|History of Present Illness|612,619|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|612,619|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|612,619|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|624,628|false|false|false|||seen
Finding|Finding|History of Present Illness|664,668|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|History of Present Illness|664,668|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|History of Present Illness|664,668|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|History of Present Illness|676,681|false|false|false|||noted
Finding|Functional Concept|History of Present Illness|690,696|false|false|false|C0234621|Visual|visual
Finding|Sign or Symptom|History of Present Illness|690,711|false|false|false|C0233763|Hallucinations, Visual|visual hallucinations
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|697,711|false|false|false|C0018524|Hallucinations|hallucinations
Event|Event|History of Present Illness|697,711|false|false|false|||hallucinations
Finding|Idea or Concept|History of Present Illness|716,725|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Event|Event|History of Present Illness|726,730|false|false|false|||gait
Finding|Finding|History of Present Illness|726,730|false|false|false|C0016928|Gait|gait
Event|Event|History of Present Illness|731,739|false|false|false|||freezing
Finding|Functional Concept|History of Present Illness|731,739|false|false|false|C0677542|Frozen behavior|freezing
Phenomenon|Natural Phenomenon or Process|History of Present Illness|731,739|false|false|false|C0016701|Freezing|freezing
Finding|Finding|History of Present Illness|749,753|false|false|false|C0016928|Gait|gait
Event|Event|History of Present Illness|754,762|false|false|false|||freezing
Finding|Functional Concept|History of Present Illness|754,762|false|false|false|C0677542|Frozen behavior|freezing
Phenomenon|Natural Phenomenon or Process|History of Present Illness|754,762|false|false|false|C0016701|Freezing|freezing
Drug|Organic Chemical|History of Present Illness|768,775|false|false|false|C0721754|Mirapex|mirapex
Drug|Pharmacologic Substance|History of Present Illness|768,775|false|false|false|C0721754|Mirapex|mirapex
Event|Event|History of Present Illness|768,775|false|false|false|||mirapex
Event|Event|History of Present Illness|780,789|false|false|false|||increased
Finding|Intellectual Product|History of Present Illness|808,812|false|false|false|C1561540|Transaction counts and value totals - week|week
Finding|Idea or Concept|History of Present Illness|818,822|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Finding|Intellectual Product|History of Present Illness|818,822|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Event|Event|History of Present Illness|823,827|false|false|false|||dose
Event|Event|History of Present Illness|865,873|false|false|false|||titrated
Drug|Pharmacologic Substance|History of Present Illness|878,886|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Event|Event|History of Present Illness|878,886|false|false|false|||medicine
Event|Event|History of Present Illness|911,916|false|false|false|||began
Finding|Functional Concept|History of Present Illness|925,931|false|false|false|C0234621|Visual|visual
Finding|Sign or Symptom|History of Present Illness|925,946|false|false|false|C0233763|Hallucinations, Visual|visual hallucinations
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|932,946|false|false|false|C0018524|Hallucinations|hallucinations
Event|Event|History of Present Illness|932,946|false|false|false|||hallucinations
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|951,960|false|false|false|C0009676|Confusion|confusion
Event|Event|History of Present Illness|951,960|false|false|false|||confusion
Finding|Finding|History of Present Illness|951,960|false|false|false|C0683369|Clouded consciousness|confusion
Event|Event|History of Present Illness|987,998|false|false|false|||recommended
Event|Event|History of Present Illness|999,1009|false|false|false|||decreasing
Event|Event|History of Present Illness|1014,1018|false|false|false|||dose
Event|Event|History of Present Illness|1028,1031|false|false|false|||TID
Event|Event|History of Present Illness|1046,1053|false|false|false|||changes
Finding|Functional Concept|History of Present Illness|1046,1053|false|false|false|C0392747|Changing|changes
Drug|Organic Chemical|History of Present Illness|1061,1068|false|false|false|C0721754|Mirapex|Mirapex
Drug|Pharmacologic Substance|History of Present Illness|1061,1068|false|false|false|C0721754|Mirapex|Mirapex
Finding|Body Substance|History of Present Illness|1074,1081|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1074,1081|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1074,1081|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|1097,1102|false|false|false|||noted
Finding|Functional Concept|History of Present Illness|1103,1114|false|false|false|C0205329|Progressive|progressive
Finding|Finding|History of Present Illness|1115,1119|false|false|false|C0016928|Gait|gait
Event|Event|History of Present Illness|1120,1129|false|false|false|||stiffness
Finding|Sign or Symptom|History of Present Illness|1120,1129|false|false|false|C0427008|Stiffness|stiffness
Event|Event|History of Present Illness|1134,1143|false|false|false|||increased
Event|Event|History of Present Illness|1144,1154|false|false|false|||difficulty
Finding|Finding|History of Present Illness|1144,1154|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Event|Event|History of Present Illness|1174,1182|false|false|false|||resulted
Event|Event|History of Present Illness|1186,1196|false|false|false|||difficulty
Finding|Finding|History of Present Illness|1186,1196|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Finding|Finding|History of Present Illness|1186,1201|false|false|false|C0332218|Difficult (qualifier value)|difficulty with
Event|Event|History of Present Illness|1209,1216|false|false|false|||getting
Event|Event|History of Present Illness|1233,1240|false|false|false|||leading
Event|Event|History of Present Illness|1244,1252|false|false|false|||episodes
Disorder|Disease or Syndrome|History of Present Illness|1256,1268|false|false|false|C0021167|Incontinence|incontinence
Event|Event|History of Present Illness|1256,1268|false|false|false|||incontinence
Event|Event|History of Present Illness|1296,1306|false|false|false|||reassuring
Procedure|Health Care Activity|History of Present Illness|1296,1306|false|false|false|C0557055|Reassuring (procedure)|reassuring
Finding|Idea or Concept|History of Present Illness|1317,1320|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|History of Present Illness|1317,1320|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|History of Present Illness|1324,1336|false|false|false|||presentation
Finding|Idea or Concept|History of Present Illness|1324,1336|false|false|false|C0449450|Presentation|presentation
Finding|Idea or Concept|History of Present Illness|1344,1352|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Body Substance|History of Present Illness|1358,1365|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1358,1365|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1358,1365|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|1366,1371|false|false|false|||began
Event|Event|History of Present Illness|1375,1385|false|false|false|||experience
Finding|Mental Process|History of Present Illness|1375,1385|false|false|false|C0237607;C0596545|Experience;Experience (Practice)|experience
Finding|Functional Concept|History of Present Illness|1386,1392|false|false|false|C0234621|Visual|visual
Finding|Sign or Symptom|History of Present Illness|1386,1407|false|false|false|C0233763|Hallucinations, Visual|visual hallucinations
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|1393,1407|false|false|false|C0018524|Hallucinations|hallucinations
Event|Event|History of Present Illness|1393,1407|false|false|false|||hallucinations
Finding|Functional Concept|History of Present Illness|1413,1418|false|false|false|C1513492|motor movement|motor
Disorder|Disease or Syndrome|History of Present Illness|1419,1424|false|false|false|C2936910|Cross syndrome|cross
Finding|Conceptual Entity|History of Present Illness|1419,1424|false|false|false|C2828360|Traverse|cross
Attribute|Clinical Attribute|History of Present Illness|1425,1429|false|false|false|C1315098||race
Event|Event|History of Present Illness|1425,1429|false|false|false|||race
Finding|Gene or Genome|History of Present Illness|1425,1429|false|false|false|C1412374;C1706779|AMACR gene;AMACR wt Allele|race
Procedure|Molecular Biology Research Technique|History of Present Illness|1425,1429|false|false|false|C5551096|Rapid Amplification of cDNA Ends|race
Event|Event|History of Present Illness|1437,1445|false|false|false|||backyard
Finding|Finding|History of Present Illness|1467,1473|false|false|false|C1561668|History of fall|a fall
Event|Event|History of Present Illness|1469,1473|false|false|false|||fall
Finding|Finding|History of Present Illness|1469,1473|false|false|false|C0085639|Falls|fall
Event|Event|History of Present Illness|1480,1492|false|false|false|||transferring
Event|Event|History of Present Illness|1502,1507|false|false|false|||couch
Event|Event|History of Present Illness|1533,1539|false|false|false|||unable
Finding|Finding|History of Present Illness|1533,1539|false|false|false|C1299582|Unable|unable
Anatomy|Anatomical Structure|History of Present Illness|1559,1564|false|false|false|C3714591|Floor (anatomic)|floor
Finding|Finding|History of Present Illness|1570,1574|true|false|false|C0085639|Falls|fall
Event|Event|History of Present Illness|1579,1588|true|false|false|||witnessed
Anatomy|Body Location or Region|History of Present Illness|1606,1610|true|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1606,1610|true|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|History of Present Illness|1606,1610|true|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1606,1610|true|false|false|C0876917|Procedure on head|head
Event|Event|History of Present Illness|1611,1617|true|false|false|||strike
Event|Occupational Activity|History of Present Illness|1611,1617|true|false|false|C0038452|Strikes, Employee|strike
Finding|Body Substance|History of Present Illness|1627,1634|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1627,1634|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1627,1634|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|1647,1651|false|false|false|||gait
Finding|Finding|History of Present Illness|1647,1651|false|false|false|C0016928|Gait|gait
Event|Event|History of Present Illness|1664,1672|false|false|false|||worsened
Event|Event|History of Present Illness|1690,1695|false|false|false|||hours
Event|Event|History of Present Illness|1727,1733|false|false|false|||unable
Finding|Finding|History of Present Illness|1727,1733|false|false|false|C1299582|Unable|unable
Event|Event|History of Present Illness|1737,1745|false|false|false|||ambulate
Finding|Finding|History of Present Illness|1737,1745|false|false|false|C4036205|Ambulate|ambulate
Event|Event|History of Present Illness|1753,1756|false|false|false|||own
Finding|Finding|History of Present Illness|1753,1756|false|false|false|C5939094|Own|own
Finding|Body Substance|History of Present Illness|1762,1769|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1762,1769|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1762,1769|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|1781,1787|false|false|false|||called
Event|Event|History of Present Illness|1808,1819|false|false|false|||recommended
Event|Event|History of Present Illness|1820,1832|false|false|false|||presentation
Finding|Idea or Concept|History of Present Illness|1820,1832|false|false|false|C0449450|Presentation|presentation
Finding|Body Substance|History of Present Illness|1861,1868|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1861,1868|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1861,1868|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|1873,1881|false|false|false|||afebrile
Finding|Finding|History of Present Illness|1873,1881|false|false|false|C0277797|Apyrexial|afebrile
Disorder|Disease or Syndrome|History of Present Illness|1883,1886|false|false|false|C0751781|Dentatorubral-Pallidoluysian Atrophy|HRs
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1883,1886|false|false|false|C1568891|HGS protein, human|HRs
Drug|Biologically Active Substance|History of Present Illness|1883,1886|false|false|false|C1568891|HGS protein, human|HRs
Event|Event|History of Present Illness|1883,1886|false|false|false|||HRs
Finding|Gene or Genome|History of Present Illness|1883,1886|false|false|false|C1366514;C1415473;C1419996;C1708271;C5575450;C5780798|ATN1 wt Allele;HARS1 gene;HARS1 wt Allele;HGS gene;HGS wt Allele;SRSF5 gene|HRs
Attribute|Clinical Attribute|History of Present Illness|1910,1914|false|false|false|C2317096|Saturation of Peripheral Oxygen|SpO2
Event|Event|History of Present Illness|1927,1931|false|false|false|||exam
Finding|Functional Concept|History of Present Illness|1927,1931|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|History of Present Illness|1927,1931|false|false|false|C0582103|Medical Examination|exam
Event|Event|History of Present Illness|1939,1944|false|false|false|||noted
Event|Event|History of Present Illness|1953,1964|false|false|false|||cogwheeling
Finding|Sign or Symptom|History of Present Illness|1953,1964|false|false|false|C0151564|Cogwheel Rigidity|cogwheeling
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1974,1985|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Event|Event|History of Present Illness|1990,1998|false|false|false|||decrease
Finding|Finding|History of Present Illness|1990,1998|false|false|false|C0392756|Reduced|decrease
Event|Event|History of Present Illness|2003,2011|false|false|false|||strength
Finding|Idea or Concept|History of Present Illness|2003,2011|false|false|false|C0808080|Strength (attribute)|strength
Event|Event|History of Present Illness|2013,2017|false|false|false|||Labs
Lab|Laboratory or Test Result|History of Present Illness|2013,2017|false|false|false|C0587081|Laboratory test finding|Labs
Event|Event|History of Present Illness|2023,2033|false|false|false|||remarkable
Event|Event|History of Present Illness|2040,2048|false|false|false|||negative
Finding|Classification|History of Present Illness|2040,2048|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|History of Present Illness|2040,2048|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|History of Present Illness|2040,2048|false|false|false|C5237010|Expression Negative|negative
Event|Event|History of Present Illness|2049,2054|false|false|false|||urine
Finding|Body Substance|History of Present Illness|2049,2054|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|History of Present Illness|2049,2054|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|History of Present Illness|2049,2054|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Drug|Indicator, Reagent, or Diagnostic Aid|History of Present Illness|2059,2064|false|false|false|C5575602|Cell Culture Serum|serum
Finding|Body Substance|History of Present Illness|2059,2064|false|false|false|C0229671;C1546774;C1550100|Serum;Serum specimen|serum
Finding|Intellectual Product|History of Present Illness|2059,2064|false|false|false|C0229671;C1546774;C1550100|Serum;Serum specimen|serum
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|2065,2068|false|false|false|C3177193|TOX protein, human|tox
Drug|Biologically Active Substance|History of Present Illness|2065,2068|false|false|false|C3177193|TOX protein, human|tox
Event|Event|History of Present Illness|2065,2068|false|false|false|||tox
Finding|Gene or Genome|History of Present Illness|2065,2068|false|false|false|C1847320|TOX gene|tox
Event|Event|History of Present Illness|2085,2094|true|false|false|||hemolyzed
Event|Event|History of Present Illness|2103,2106|true|false|false|||EKG
Finding|Intellectual Product|History of Present Illness|2103,2106|true|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|History of Present Illness|2103,2106|true|false|false|C1623258|Electrocardiography|EKG
Event|Event|History of Present Illness|2107,2114|true|false|false|||changes
Finding|Functional Concept|History of Present Illness|2107,2114|true|false|false|C0392747|Changing|changes
Finding|Classification|History of Present Illness|2117,2125|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|History of Present Illness|2117,2125|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|History of Present Illness|2117,2125|false|false|false|C5237010|Expression Negative|negative
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|2126,2134|false|false|false|C0041199|Troponin|troponin
Drug|Biologically Active Substance|History of Present Illness|2126,2134|false|false|false|C0041199|Troponin|troponin
Event|Event|History of Present Illness|2126,2134|false|false|false|||troponin
Procedure|Laboratory Procedure|History of Present Illness|2126,2134|false|false|false|C0523952|Troponin measurement|troponin
Event|Event|History of Present Illness|2143,2147|false|false|false|||LFTs
Anatomy|Cell Component|History of Present Illness|2162,2165|false|false|false|C2263086|Nuclear cap binding complex location|CBC
Event|Event|History of Present Illness|2162,2165|false|false|false|||CBC
Procedure|Laboratory Procedure|History of Present Illness|2162,2165|false|false|false|C0009555|Complete Blood Count|CBC
Anatomy|Body Location or Region|History of Present Illness|2168,2173|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|History of Present Illness|2168,2173|true|false|false|C0741025|Chest problem|Chest
Event|Event|History of Present Illness|2174,2178|true|false|false|||Xray
Phenomenon|Natural Phenomenon or Process|History of Present Illness|2174,2178|true|false|false|C0043309|Roentgen Rays|Xray
Procedure|Diagnostic Procedure|History of Present Illness|2174,2178|true|false|false|C0043299|Diagnostic radiologic examination|Xray
Event|Event|History of Present Illness|2179,2185|true|false|false|||showed
Finding|Intellectual Product|History of Present Illness|2189,2194|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2195,2202|true|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|History of Present Illness|2195,2202|true|false|false|C1951340|Process Pharmacologic Substance|process
Event|Event|History of Present Illness|2195,2202|true|false|false|||process
Finding|Functional Concept|History of Present Illness|2195,2202|true|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|History of Present Illness|2195,2202|true|false|false|C1522240|Process|process
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|2207,2210|true|false|false|C5849006|CTH protein, human|CTH
Drug|Enzyme|History of Present Illness|2207,2210|true|false|false|C5849006|CTH protein, human|CTH
Event|Event|History of Present Illness|2207,2210|true|false|false|||CTH
Finding|Gene or Genome|History of Present Illness|2207,2210|true|false|false|C1413792;C1538070|CTH gene;VSIG2 gene|CTH
Event|Event|History of Present Illness|2215,2225|true|false|false|||reassuring
Procedure|Health Care Activity|History of Present Illness|2215,2225|true|false|false|C0557055|Reassuring (procedure)|reassuring
Event|Event|History of Present Illness|2234,2243|false|false|false|||evaluated
Event|Event|History of Present Illness|2261,2272|false|false|false|||recommended
Event|Event|History of Present Illness|2273,2282|false|false|false|||admission
Procedure|Health Care Activity|History of Present Illness|2273,2282|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Drug|Pharmacologic Substance|History of Present Illness|2286,2294|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Event|Event|History of Present Illness|2286,2294|false|false|false|||medicine
Event|Event|History of Present Illness|2299,2306|false|false|false|||failure
Finding|Functional Concept|History of Present Illness|2299,2306|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|History of Present Illness|2299,2306|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|History of Present Illness|2299,2306|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|History of Present Illness|2310,2316|false|false|false|||thrive
Event|Event|History of Present Illness|2321,2329|false|false|false|||continue
Finding|Body Substance|History of Present Illness|2334,2341|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|2334,2341|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|2334,2341|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|2344,2348|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|History of Present Illness|2344,2348|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|History of Present Illness|2344,2348|false|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|History of Present Illness|2349,2360|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|History of Present Illness|2349,2360|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|History of Present Illness|2349,2360|false|false|false|||medications
Finding|Intellectual Product|History of Present Illness|2349,2360|false|false|false|C4284232|Medications|medications
Event|Event|History of Present Illness|2366,2374|false|false|false|||complete
Finding|Cell Function|History of Present Illness|2382,2391|false|false|false|C0311400;C1524026|Metabolic;Metabolic Process, Cellular|metabolic
Finding|Functional Concept|History of Present Illness|2382,2391|false|false|false|C0311400;C1524026|Metabolic;Metabolic Process, Cellular|metabolic
Procedure|Diagnostic Procedure|History of Present Illness|2382,2391|false|false|false|C4263342|Multisection metabolic|metabolic
Event|Event|History of Present Illness|2392,2398|false|false|false|||workup
Finding|Body Substance|History of Present Illness|2404,2411|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|2404,2411|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|2404,2411|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|2426,2430|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|History of Present Illness|2426,2430|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|History of Present Illness|2426,2430|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|History of Present Illness|2431,2442|false|false|false|C0074710|pramipexole|pramipexole
Drug|Pharmacologic Substance|History of Present Illness|2431,2442|false|false|false|C0074710|pramipexole|pramipexole
Event|Event|History of Present Illness|2431,2442|false|false|false|||pramipexole
Drug|Organic Chemical|History of Present Illness|2447,2458|false|false|false|C0085542|pravastatin|pravastatin
Drug|Pharmacologic Substance|History of Present Illness|2447,2458|false|false|false|C0085542|pravastatin|pravastatin
Event|Event|History of Present Illness|2447,2458|false|false|false|||pravastatin
Event|Event|History of Present Illness|2473,2481|false|false|false|||admitted
Event|Activity|History of Present Illness|2489,2496|false|false|false|C1706079||arrival
Event|Event|History of Present Illness|2489,2496|false|false|false|||arrival
Finding|Functional Concept|History of Present Illness|2489,2496|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Anatomy|Anatomical Structure|History of Present Illness|2504,2509|false|false|false|C3714591|Floor (anatomic)|floor
Finding|Body Substance|History of Present Illness|2515,2522|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|2515,2522|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|2515,2522|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|2526,2537|false|false|false|||comfortable
Finding|Finding|History of Present Illness|2526,2537|false|false|false|C5546696|Feeling comfortable|comfortable
Disorder|Disease or Syndrome|History of Present Illness|2541,2544|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Event|Event|History of Present Illness|2541,2544|false|false|false|||bed
Finding|Intellectual Product|History of Present Illness|2541,2544|false|false|false|C2346952|Bachelor of Education|bed
Event|Event|History of Present Illness|2557,2568|true|false|false|||accompanied
Finding|Classification|History of Present Illness|2572,2578|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|History of Present Illness|2572,2578|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|History of Present Illness|2572,2578|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|History of Present Illness|2572,2578|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Event|Activity|History of Present Illness|2585,2594|true|false|false|C0021822|Interview|interview
Event|Event|History of Present Illness|2585,2594|true|false|false|||interview
Finding|Intellectual Product|History of Present Illness|2585,2594|true|false|false|C0935630|Published Interview|interview
Event|Event|History of Present Illness|2599,2604|false|false|false|||knows
Finding|Idea or Concept|History of Present Illness|2624,2632|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|History of Present Illness|2663,2667|true|false|false|||sure
Finding|Intellectual Product|History of Present Illness|2663,2667|true|false|false|C4724437|SURE Test|sure
Event|Event|History of Present Illness|2687,2693|false|false|false|||begins
Event|Event|History of Present Illness|2697,2701|false|false|false|||tell
Event|Event|History of Present Illness|2713,2718|false|false|false|||party
Finding|Conceptual Entity|History of Present Illness|2713,2718|false|false|true|C1518904|Party|party
Event|Event|History of Present Illness|2739,2744|false|false|false|||motor
Finding|Functional Concept|History of Present Illness|2739,2744|false|false|true|C1513492|motor movement|motor
Disorder|Disease or Syndrome|History of Present Illness|2745,2750|false|false|false|C2936910|Cross syndrome|cross
Event|Event|History of Present Illness|2745,2750|false|false|false|||cross
Finding|Conceptual Entity|History of Present Illness|2745,2750|false|false|false|C2828360|Traverse|cross
Attribute|Clinical Attribute|History of Present Illness|2751,2755|false|false|false|C1315098||race
Event|Event|History of Present Illness|2751,2755|false|false|false|||race
Finding|Gene or Genome|History of Present Illness|2751,2755|false|false|false|C1412374;C1706779|AMACR gene;AMACR wt Allele|race
Procedure|Molecular Biology Research Technique|History of Present Illness|2751,2755|false|false|false|C5551096|Rapid Amplification of cDNA Ends|race
Event|Event|History of Present Illness|2780,2785|false|false|false|||asked
Event|Event|History of Present Illness|2800,2804|false|false|false|||fall
Finding|Finding|History of Present Illness|2800,2804|false|false|true|C0085639|Falls|fall
Event|Event|History of Present Illness|2809,2817|false|false|false|||mentions
Finding|Finding|History of Present Illness|2838,2844|true|false|true|C1561668|History of fall|a fall
Event|Event|History of Present Illness|2840,2844|true|false|false|||fall
Finding|Finding|History of Present Illness|2840,2844|true|false|true|C0085639|Falls|fall
Event|Event|History of Present Illness|2863,2869|true|false|false|||denies
Event|Event|History of Present Illness|2874,2880|true|false|false|||fevers
Finding|Sign or Symptom|History of Present Illness|2874,2880|true|false|false|C0015967|Fever|fevers
Event|Event|History of Present Illness|2882,2888|true|false|false|||chills
Finding|Sign or Symptom|History of Present Illness|2882,2888|true|false|false|C0085593|Chills|chills
Drug|Organic Chemical|History of Present Illness|2890,2895|true|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|2890,2895|true|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|History of Present Illness|2890,2895|true|false|false|||cough
Finding|Sign or Symptom|History of Present Illness|2890,2895|true|false|false|C0010200|Coughing|cough
Anatomy|Body Location or Region|History of Present Illness|2897,2902|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|2897,2902|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|2897,2907|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|2897,2907|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|2903,2907|false|false|false|C2598155||pain
Event|Event|History of Present Illness|2903,2907|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|2903,2907|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|2903,2907|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|2903,2918|false|false|false|C0000737|Abdominal Pain|pain, abdominal
Anatomy|Body Location or Region|History of Present Illness|2909,2918|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|History of Present Illness|2909,2923|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|History of Present Illness|2919,2923|false|false|false|C2598155||pain
Event|Event|History of Present Illness|2919,2923|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|2919,2923|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|2919,2923|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|History of Present Illness|2925,2931|false|false|false|C4255480||nausea
Event|Event|History of Present Illness|2925,2931|false|false|false|||nausea
Finding|Sign or Symptom|History of Present Illness|2925,2931|false|false|false|C0027497|Nausea|nausea
Event|Event|History of Present Illness|2933,2941|false|false|false|||diarrhea
Finding|Finding|History of Present Illness|2933,2941|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|History of Present Illness|2933,2941|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Event|Event|History of Present Illness|2946,2953|false|false|false|||dysuria
Finding|Sign or Symptom|History of Present Illness|2946,2953|false|false|false|C0013428|Dysuria|dysuria
Event|Event|History of Present Illness|2957,2963|false|false|false|||REVIEW
Finding|Idea or Concept|History of Present Illness|2957,2963|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|REVIEW
Finding|Intellectual Product|History of Present Illness|2957,2963|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|REVIEW
Finding|Functional Concept|History of Present Illness|2957,2966|false|false|false|C0699752|Review of|REVIEW OF
Attribute|Clinical Attribute|History of Present Illness|2957,2974|false|false|false|C0488564;C0488565||REVIEW OF SYSTEMS
Procedure|Health Care Activity|History of Present Illness|2957,2974|false|false|false|C0489633|Review of systems (procedure)|REVIEW OF SYSTEMS
Event|Event|History of Present Illness|2967,2974|false|false|false|||SYSTEMS
Finding|Functional Concept|History of Present Illness|2967,2974|false|false|false|C0449913|System|SYSTEMS
Disorder|Disease or Syndrome|History of Present Illness|2999,3002|false|false|false|C0268529|Proline dehydrogenase deficiency|HPI
Event|Event|History of Present Illness|2999,3002|false|false|false|||HPI
Finding|Finding|History of Present Illness|2999,3002|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Finding|Molecular Function|History of Present Illness|2999,3002|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Event|Event|History of Present Illness|3024,3030|false|false|false|||review
Finding|Idea or Concept|History of Present Illness|3024,3030|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Intellectual Product|History of Present Illness|3024,3030|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Functional Concept|History of Present Illness|3024,3033|false|false|false|C0699752|Review of|review of
Attribute|Clinical Attribute|History of Present Illness|3024,3041|false|false|false|C0488564;C0488565||review of systems
Procedure|Health Care Activity|History of Present Illness|3024,3041|false|false|false|C0489633|Review of systems (procedure)|review of systems
Event|Event|History of Present Illness|3034,3041|false|false|false|||systems
Finding|Functional Concept|History of Present Illness|3034,3041|false|false|false|C0449913|System|systems
Event|Event|History of Present Illness|3053,3059|false|false|false|||normal
Event|Event|History of Present Illness|3060,3066|false|false|false|||limits
Finding|Functional Concept|History of Present Illness|3060,3066|false|false|false|C0439801|Limited (extensiveness)|limits
Disorder|Disease or Syndrome|Past Medical History|3097,3104|false|false|false|C0012634|Disease|disease
Event|Event|Past Medical History|3097,3104|false|false|false|||disease
Anatomy|Anatomical Structure|Past Medical History|3109,3113|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|Body
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|3109,3113|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|Body
Finding|Intellectual Product|Past Medical History|3109,3113|false|false|false|C1551342|Document Body|Body
Disorder|Mental or Behavioral Dysfunction|Past Medical History|3114,3122|false|false|false|C0011265;C0497327|Dementia;Presenile dementia|Dementia
Event|Event|Past Medical History|3114,3122|false|false|false|||Dementia
Disorder|Disease or Syndrome|Past Medical History|3124,3136|false|false|false|C0242339|Dyslipidemias|dyslipidemia
Event|Event|Past Medical History|3124,3136|false|false|false|||dyslipidemia
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|3138,3146|false|false|false|C0033572;C4266527|Prostate;Structure of prostate (body structure)|prostate
Disorder|Disease or Syndrome|Past Medical History|3138,3146|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|prostate
Disorder|Neoplastic Process|Past Medical History|3138,3146|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|prostate
Disorder|Neoplastic Process|Past Medical History|3138,3153|false|false|false|C0376358;C0600139|Malignant neoplasm of prostate;Prostate carcinoma|prostate cancer
Disorder|Neoplastic Process|Past Medical History|3147,3153|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Past Medical History|3147,3153|false|false|false|||cancer
Procedure|Therapeutic or Preventive Procedure|Past Medical History|3159,3172|false|false|false|C0033573|Prostatectomy|prostatectomy
Event|Event|Family Medical History|3216,3222|false|false|false|||mother
Finding|Idea or Concept|Family Medical History|3216,3222|false|false|false|C1546508|Relationship - Mother|mother
Event|Event|Family Medical History|3223,3227|false|false|false|||died
Attribute|Clinical Attribute|Family Medical History|3231,3234|false|false|false|C1114365||age
Drug|Biologically Active Substance|Family Medical History|3231,3234|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|Family Medical History|3231,3234|false|false|false|C0162574|Glycation End Products, Advanced|age
Finding|Finding|Family Medical History|3243,3250|false|false|false|C0231337|Senility|old age
Attribute|Clinical Attribute|Family Medical History|3247,3250|false|false|false|C1114365||age
Drug|Biologically Active Substance|Family Medical History|3247,3250|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|Family Medical History|3247,3250|false|false|false|C0162574|Glycation End Products, Advanced|age
Event|Event|Family Medical History|3247,3250|false|false|false|||age
Event|Event|Family Medical History|3257,3263|false|false|false|||father
Finding|Conceptual Entity|Family Medical History|3257,3263|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Finding|Idea or Concept|Family Medical History|3257,3263|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Event|Event|Family Medical History|3264,3268|false|false|false|||died
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3272,3280|false|false|false|C0033572;C4266527|Prostate;Structure of prostate (body structure)|prostate
Disorder|Disease or Syndrome|Family Medical History|3272,3280|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|prostate
Disorder|Neoplastic Process|Family Medical History|3272,3280|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|prostate
Disorder|Neoplastic Process|Family Medical History|3272,3287|false|false|false|C0376358;C0600139|Malignant neoplasm of prostate;Prostate carcinoma|prostate cancer
Disorder|Neoplastic Process|Family Medical History|3281,3287|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Family Medical History|3281,3287|false|false|false|||cancer
Event|Event|Family Medical History|3307,3312|false|false|false|||older
Finding|Conceptual Entity|Family Medical History|3314,3320|false|false|false|C1546515;C1704647|Relationship - Sister;Sister - courtesy title|sister
Attribute|Clinical Attribute|Family Medical History|3322,3325|false|false|false|C1114365||age
Drug|Biologically Active Substance|Family Medical History|3322,3325|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|Family Medical History|3322,3325|false|false|false|C0162574|Glycation End Products, Advanced|age
Event|Event|Family Medical History|3322,3325|false|false|false|||age
Event|Event|Family Medical History|3344,3350|false|false|false|||sister
Finding|Conceptual Entity|Family Medical History|3344,3350|false|false|false|C1546515;C1704647|Relationship - Sister;Sister - courtesy title|sister
Attribute|Clinical Attribute|Family Medical History|3352,3355|false|false|false|C1114365||age
Drug|Biologically Active Substance|Family Medical History|3352,3355|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|Family Medical History|3352,3355|false|false|false|C0162574|Glycation End Products, Advanced|age
Finding|Conceptual Entity|Family Medical History|3380,3387|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|brother
Finding|Idea or Concept|Family Medical History|3380,3387|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|brother
Attribute|Clinical Attribute|Family Medical History|3389,3392|false|false|false|C1114365||age
Drug|Biologically Active Substance|Family Medical History|3389,3392|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|Family Medical History|3389,3392|false|false|false|C0162574|Glycation End Products, Advanced|age
Event|Event|Family Medical History|3389,3392|false|false|false|||age
Event|Event|Family Medical History|3402,3407|false|false|false|||noted
Event|Event|Family Medical History|3418,3427|false|false|false|||daughters
Finding|Classification|Family Medical History|3442,3448|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Family Medical History|3442,3448|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Family Medical History|3442,3448|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Family Medical History|3442,3448|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Event|Event|Family Medical History|3449,3456|true|false|false|||history
Finding|Conceptual Entity|Family Medical History|3449,3456|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|3449,3456|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Family Medical History|3449,3456|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|3449,3459|true|false|false|C0262926|Medical History|history of
Event|Event|Family Medical History|3471,3478|true|false|false|||illness
Finding|Sign or Symptom|Family Medical History|3471,3478|true|false|false|C0221423|Illness (finding)|illness
Disorder|Mental or Behavioral Dysfunction|Family Medical History|3482,3490|false|false|false|C0011265;C0497327|Dementia;Presenile dementia|dementia
Event|Event|Family Medical History|3482,3490|false|false|false|||dementia
Finding|Classification|Family Medical History|3505,3511|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Family Medical History|3505,3511|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Family Medical History|3505,3511|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Family Medical History|3505,3511|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Event|Event|Family Medical History|3512,3519|true|false|false|||history
Finding|Conceptual Entity|Family Medical History|3512,3519|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|3512,3519|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Family Medical History|3512,3519|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|3512,3522|true|false|false|C0262926|Medical History|history of
Finding|Mental Process|Family Medical History|3542,3548|true|false|false|C0229992|Psyche structure|mental
Disorder|Mental or Behavioral Dysfunction|Family Medical History|3542,3558|true|false|false|C0004936|Mental disorders|mental disorders
Disorder|Disease or Syndrome|Family Medical History|3549,3558|true|false|false|C0012634|Disease|disorders
Event|Event|Family Medical History|3549,3558|true|false|false|||disorders
Event|Event|Family Medical History|3567,3575|false|false|false|||learning
Finding|Mental Process|Family Medical History|3567,3575|false|false|false|C0023185|Learning|learning
Procedure|Educational Activity|Family Medical History|3567,3575|false|false|false|C0013621|Knowledge acquisition|learning
Attribute|Clinical Attribute|Family Medical History|3576,3586|false|false|false|C5240435||disability
Event|Event|Family Medical History|3576,3586|false|false|false|||disability
Finding|Finding|Family Medical History|3576,3586|false|false|false|C0231170|Disability|disability
Disorder|Mental or Behavioral Dysfunction|Family Medical History|3590,3594|false|false|false|C1263846|Attention deficit hyperactivity disorder|ADHD
Event|Event|Family Medical History|3590,3594|false|false|false|||ADHD
Finding|Classification|Family Medical History|3609,3615|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Family Medical History|3609,3615|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Family Medical History|3609,3615|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Family Medical History|3609,3615|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Finding|Family Medical History|3609,3623|true|false|false|C0241889|Family Medical History|family history
Finding|Finding|Family Medical History|3609,3626|true|false|false|C0241889|Family Medical History|family history of
Event|Event|Family Medical History|3616,3623|true|false|false|||history
Finding|Conceptual Entity|Family Medical History|3616,3623|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|3616,3623|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Family Medical History|3616,3623|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|3616,3626|true|false|false|C0262926|Medical History|history of
Event|Event|Family Medical History|3627,3638|true|false|false|||psychiatric
Finding|Finding|Family Medical History|3627,3638|true|false|false|C0205487;C1548428|Psychiatric;Referral type - Psychiatric|psychiatric
Finding|Functional Concept|Family Medical History|3627,3638|true|false|false|C0205487;C1548428|Psychiatric;Referral type - Psychiatric|psychiatric
Procedure|Therapeutic or Preventive Procedure|Family Medical History|3627,3638|true|false|false|C3526598|Psychiatric service|psychiatric
Event|Event|Family Medical History|3639,3647|true|false|false|||problems
Finding|Idea or Concept|Family Medical History|3639,3647|true|false|false|C1546466|Problems - What subject filter|problems
Procedure|Health Care Activity|General Exam|3666,3675|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|General Exam|3676,3684|false|false|false|||PHYSICAL
Finding|Finding|General Exam|3676,3684|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|General Exam|3676,3684|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|General Exam|3676,3684|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|General Exam|3676,3689|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|General Exam|3676,3689|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Event|Event|General Exam|3685,3689|false|false|false|||EXAM
Finding|Functional Concept|General Exam|3685,3689|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|3685,3689|false|false|false|C0582103|Medical Examination|EXAM
Event|Event|General Exam|3716,3722|false|false|false|||VITALS
Event|Event|General Exam|3724,3732|false|false|false|||reviewed
Event|Event|General Exam|3736,3739|false|false|false|||OMR
Finding|Gene or Genome|General Exam|3736,3739|false|false|false|C1412647|ATP5F1A gene|OMR
Event|Event|General Exam|3741,3748|false|false|false|||GENERAL
Finding|Classification|General Exam|3741,3748|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|General Exam|3741,3748|false|false|false|C3812897|General medical service|GENERAL
Attribute|Clinical Attribute|General Exam|3750,3755|false|false|false|C5890168||Alert
Drug|Organic Chemical|General Exam|3750,3755|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|General Exam|3750,3755|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|General Exam|3750,3755|false|false|false|||Alert
Finding|Finding|General Exam|3750,3755|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|General Exam|3750,3755|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|General Exam|3750,3755|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|General Exam|3760,3771|false|false|false|||interactive
Finding|Functional Concept|General Exam|3760,3771|false|false|false|C1704675|Interaction|interactive
Finding|Finding|General Exam|3773,3793|false|false|false|C2051415|patient appears in no acute distress (physical finding)|In no acute distress
Finding|Intellectual Product|General Exam|3779,3784|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|General Exam|3785,3793|true|false|false|||distress
Finding|Finding|General Exam|3785,3793|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|General Exam|3785,3793|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|General Exam|3795,3800|false|false|false|C1512338|HEENT|HEENT
Event|Event|General Exam|3802,3807|false|false|false|||PERRL
Finding|Finding|General Exam|3802,3807|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Event|Event|General Exam|3809,3813|false|false|false|||EOMI
Anatomy|Body Part, Organ, or Organ Component|General Exam|3815,3821|true|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|General Exam|3815,3821|true|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|General Exam|3815,3821|true|false|false|||Sclera
Procedure|Health Care Activity|General Exam|3815,3821|true|false|false|C2228481|examination of sclera|Sclera
Event|Event|General Exam|3822,3831|true|false|false|||anicteric
Finding|Finding|General Exam|3822,3831|true|false|false|C0205180|Anicteric|anicteric
Drug|Biomedical or Dental Material|General Exam|3844,3853|true|false|false|C1272883|Injection|injection
Event|Event|General Exam|3844,3853|true|false|false|||injection
Finding|Functional Concept|General Exam|3844,3853|true|false|false|C1828121|Injection Route of Administration|injection
Procedure|Therapeutic or Preventive Procedure|General Exam|3844,3853|true|false|false|C0021485;C1533685|Injection of therapeutic agent;Injection procedure|injection
Anatomy|Body Part, Organ, or Organ Component|General Exam|3855,3858|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|General Exam|3855,3858|false|false|false|C0026987|Myelofibrosis|MMM
Event|Event|General Exam|3855,3858|false|false|false|||MMM
Anatomy|Body Location or Region|General Exam|3860,3864|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|General Exam|3860,3864|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|General Exam|3860,3864|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Anatomy|Body Location or Region|General Exam|3869,3877|true|false|false|C0027530|Neck|cervical
Disorder|Disease or Syndrome|General Exam|3869,3893|true|false|false|C0235592|Cervical lymphadenopathy|cervical lymphadenopathy
Finding|Finding|General Exam|3869,3893|true|false|false|C4551446|Swollen lymph nodes in the neck|cervical lymphadenopathy
Disorder|Disease or Syndrome|General Exam|3878,3893|true|false|false|C0497156|Lymphadenopathy|lymphadenopathy
Event|Event|General Exam|3878,3893|true|false|false|||lymphadenopathy
Finding|Sign or Symptom|General Exam|3878,3893|true|false|false|C4282165|Swollen Lymph Node|lymphadenopathy
Event|Event|General Exam|3898,3901|true|false|false|||JVD
Finding|Finding|General Exam|3898,3901|true|false|false|C0425687|Jugular venous engorgement|JVD
Anatomy|Body Part, Organ, or Organ Component|General Exam|3903,3910|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|General Exam|3903,3910|false|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Event|General Exam|3920,3926|false|false|false|||rhythm
Finding|Finding|General Exam|3920,3926|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|General Exam|3920,3926|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Event|Activity|General Exam|3935,3939|false|false|false|C0871208|Rating (action)|rate
Event|Event|General Exam|3935,3939|false|false|false|||rate
Finding|Idea or Concept|General Exam|3935,3939|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|General Exam|3963,3970|true|false|false|||murmurs
Finding|Finding|General Exam|3963,3970|true|false|false|C0018808|Heart murmur|murmurs
Event|Event|General Exam|3971,3975|true|false|false|||rubs
Finding|Finding|General Exam|3971,3975|true|false|false|C0232267|Pericardial friction rub|rubs
Event|Event|General Exam|3976,3983|true|false|false|||gallops
Anatomy|Body Part, Organ, or Organ Component|General Exam|3985,3990|false|false|false|C0024109|Lung|LUNGS
Event|Event|General Exam|3992,3997|false|false|false|||Clear
Finding|Idea or Concept|General Exam|3992,3997|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|General Exam|4001,4013|false|false|false|||auscultation
Procedure|Diagnostic Procedure|General Exam|4001,4013|false|false|false|C0004339|Auscultation|auscultation
Event|Event|General Exam|4030,4037|true|false|false|||wheezes
Finding|Sign or Symptom|General Exam|4030,4037|true|false|false|C0043144|Wheezing|wheezes
Event|Event|General Exam|4039,4046|true|false|false|||rhonchi
Finding|Finding|General Exam|4039,4046|true|false|false|C0035508|Rhonchi|rhonchi
Event|Event|General Exam|4050,4055|true|false|false|||rales
Finding|Finding|General Exam|4050,4055|true|false|false|C0034642;C0240859|Basilar Rales;Rales|rales
Event|Event|General Exam|4060,4069|true|false|false|||increased
Finding|Finding|General Exam|4060,4069|true|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Functional Concept|General Exam|4060,4069|true|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Sign or Symptom|General Exam|4060,4087|true|false|false|C0859927|Increased work of breathing|increased work of breathing
Event|Event|General Exam|4070,4074|true|false|false|||work
Event|Occupational Activity|General Exam|4070,4074|true|false|false|C0043227|Work|work
Finding|Organ or Tissue Function|General Exam|4070,4087|true|false|false|C0043229|Work of Breathing|work of breathing
Attribute|Clinical Attribute|General Exam|4078,4087|true|false|false|C5885990||breathing
Event|Event|General Exam|4078,4087|true|false|false|||breathing
Finding|Finding|General Exam|4078,4087|true|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|General Exam|4078,4087|true|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|General Exam|4078,4087|true|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|General Exam|4078,4087|true|false|false|C1160636|respiratory system process|breathing
Event|Event|General Exam|4089,4093|false|false|false|||BACK
Disorder|Disease or Syndrome|General Exam|4098,4101|true|false|false|C0001365;C0038454|Acute ill-defined cerebrovascular disease;Cerebrovascular accident|CVA
Drug|Pharmacologic Substance|General Exam|4098,4101|true|false|false|C5779650|Cyclophosphamide/Doxorubicin/Vincristine|CVA
Event|Event|General Exam|4098,4101|true|false|false|||CVA
Finding|Sign or Symptom|General Exam|4098,4112|true|false|false|C0235634|Renal angle tenderness|CVA tenderness
Event|Event|General Exam|4102,4112|true|false|false|||tenderness
Finding|Mental Process|General Exam|4102,4112|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|General Exam|4102,4112|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Anatomy|Body Location or Region|General Exam|4114,4121|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|General Exam|4114,4121|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|General Exam|4114,4121|false|false|false|||ABDOMEN
Finding|Finding|General Exam|4114,4121|false|false|false|C0941288|Abdomen problem|ABDOMEN
Anatomy|Body Part, Organ, or Organ Component|General Exam|4130,4136|false|false|false|C0021853|Intestines|bowels
Event|Event|General Exam|4137,4143|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|General Exam|4137,4143|false|false|false|C0037709||sounds
Event|Event|General Exam|4149,4158|false|false|false|||distended
Finding|Finding|General Exam|4149,4158|false|false|false|C0700124|Dilated|distended
Attribute|Clinical Attribute|General Exam|4174,4178|false|false|false|C4318566|Deep Resection Margin|deep
Event|Event|General Exam|4179,4188|false|false|false|||palpation
Procedure|Diagnostic Procedure|General Exam|4179,4188|false|false|false|C0030247|Palpation|palpation
Event|Event|General Exam|4215,4227|true|false|false|||organomegaly
Finding|Finding|General Exam|4215,4227|true|false|false|C4054315|Organomegaly|organomegaly
Anatomy|Body Part, Organ, or Organ Component|General Exam|4229,4240|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Disorder|Anatomical Abnormality|General Exam|4245,4253|true|false|false|C0149651|Clubbing|clubbing
Event|Event|General Exam|4245,4253|true|false|false|||clubbing
Event|Event|General Exam|4255,4263|true|false|false|||cyanosis
Finding|Sign or Symptom|General Exam|4255,4263|true|false|false|C0010520|Cyanosis|cyanosis
Attribute|Clinical Attribute|General Exam|4268,4273|true|false|false|C1717255||edema
Event|Event|General Exam|4268,4273|true|false|false|||edema
Finding|Pathologic Function|General Exam|4268,4273|true|false|false|C0013604|Edema|edema
Drug|Food|General Exam|4275,4281|false|false|false|C5890763||Pulses
Event|Event|General Exam|4275,4281|false|false|false|||Pulses
Finding|Physiologic Function|General Exam|4275,4281|false|false|false|C0391850|Physiologic pulse|Pulses
Procedure|Health Care Activity|General Exam|4275,4281|false|false|false|C0034107|Pulse taking|Pulses
Event|Event|General Exam|4282,4284|false|false|false|||DP
Finding|Conceptual Entity|General Exam|4285,4291|false|false|false|C0442038;C0920847|Circumpennate;Radial|Radial
Anatomy|Body System|General Exam|4309,4313|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|General Exam|4309,4313|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|General Exam|4309,4313|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|General Exam|4309,4313|false|false|false|||SKIN
Finding|Body Substance|General Exam|4309,4313|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|General Exam|4309,4313|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Event|Event|General Exam|4315,4319|false|false|false|||Warm
Finding|Finding|General Exam|4315,4319|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|4315,4319|false|false|false|C0687712|warming process|Warm
Disorder|Congenital Abnormality|General Exam|4321,4324|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|Cap
Drug|Biomedical or Dental Material|General Exam|4321,4324|false|false|false|C0006935|capsule (pharmacologic)|Cap
Event|Event|General Exam|4321,4324|false|false|false|||Cap
Finding|Gene or Genome|General Exam|4321,4324|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|Cap
Procedure|Therapeutic or Preventive Procedure|General Exam|4321,4324|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|Cap
Event|Event|General Exam|4325,4331|false|false|false|||refill
Finding|Idea or Concept|General Exam|4325,4331|false|false|false|C0807726|refill|refill
Event|Event|General Exam|4340,4346|true|false|false|||rashes
Finding|Sign or Symptom|General Exam|4340,4346|true|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Event|Event|General Exam|4348,4358|false|false|false|||NEUROLOGIC
Event|Event|General Exam|4360,4364|false|false|false|||AOx3
Finding|Gene or Genome|General Exam|4366,4369|false|false|false|C1539110|CNDP2 gene|CN2
Event|Event|General Exam|4373,4379|false|false|false|||intact
Finding|Finding|General Exam|4373,4379|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Finding|General Exam|4398,4412|false|false|false|C0026826|Muscle Hypertonia|Increased tone
Event|Event|General Exam|4408,4412|false|false|false|||tone
Anatomy|Body Part, Organ, or Organ Component|General Exam|4416,4419|false|false|false|C0227192|Inferior esophageal sphincter structure|LEs
Finding|Classification|General Exam|4416,4419|false|false|false|C0023595|Lewis Blood-Group System|LEs
Finding|Idea or Concept|General Exam|4425,4433|false|false|false|C0808080|Strength (attribute)|strength
Event|Event|General Exam|4450,4459|false|false|false|||sensation
Finding|Finding|General Exam|4450,4459|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|General Exam|4450,4459|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|General Exam|4450,4459|false|false|false|C2229507|sensory exam|sensation
Finding|Body Substance|General Exam|4462,4471|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|4462,4471|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|4462,4471|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|4462,4471|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|General Exam|4472,4480|false|false|false|||PHYSICAL
Finding|Finding|General Exam|4472,4480|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|General Exam|4472,4480|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|General Exam|4472,4480|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|General Exam|4472,4485|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|General Exam|4472,4485|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Event|Event|General Exam|4481,4485|false|false|false|||EXAM
Finding|Functional Concept|General Exam|4481,4485|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|4481,4485|false|false|false|C0582103|Medical Examination|EXAM
Event|Event|General Exam|4515,4519|false|false|false|||Data
Finding|Idea or Concept|General Exam|4515,4519|false|false|false|C1511726|Data|Data
Event|Event|General Exam|4526,4533|false|false|false|||updated
Event|Event|General Exam|4550,4554|false|false|false|||Temp
Finding|Gene or Genome|General Exam|4550,4554|false|false|false|C1823816|C1orf210 gene|Temp
Procedure|Therapeutic or Preventive Procedure|General Exam|4550,4554|false|false|false|C0279848|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Temp
Event|Event|General Exam|4600,4602|false|false|false|||HR
Event|Event|General Exam|4657,4665|false|false|false|||delivery
Finding|Finding|General Exam|4657,4665|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Finding|Functional Concept|General Exam|4657,4665|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Finding|Organism Function|General Exam|4657,4665|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Procedure|Therapeutic or Preventive Procedure|General Exam|4657,4665|false|false|false|C0011209|Obstetric Delivery|delivery
Event|Event|General Exam|4673,4680|false|false|false|||GENERAL
Finding|Classification|General Exam|4673,4680|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|General Exam|4673,4680|false|false|false|C3812897|General medical service|GENERAL
Finding|Finding|General Exam|4682,4702|false|false|false|C2051415|patient appears in no acute distress (physical finding)|In no acute distress
Finding|Intellectual Product|General Exam|4688,4693|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|General Exam|4694,4702|true|false|false|||distress
Finding|Finding|General Exam|4694,4702|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|General Exam|4694,4702|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Part, Organ, or Organ Component|General Exam|4726,4733|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|General Exam|4726,4733|false|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Event|General Exam|4743,4749|false|false|false|||rhythm
Finding|Finding|General Exam|4743,4749|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|General Exam|4743,4749|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Event|Activity|General Exam|4758,4762|false|false|false|C0871208|Rating (action)|rate
Event|Event|General Exam|4758,4762|false|false|false|||rate
Finding|Idea or Concept|General Exam|4758,4762|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|General Exam|4786,4793|true|false|false|||murmurs
Finding|Finding|General Exam|4786,4793|true|false|false|C0018808|Heart murmur|murmurs
Event|Event|General Exam|4794,4798|true|false|false|||rubs
Finding|Finding|General Exam|4794,4798|true|false|false|C0232267|Pericardial friction rub|rubs
Event|Event|General Exam|4799,4806|true|false|false|||gallops
Anatomy|Body Part, Organ, or Organ Component|General Exam|4808,4813|false|false|false|C0024109|Lung|LUNGS
Event|Event|General Exam|4815,4820|false|false|false|||Clear
Finding|Idea or Concept|General Exam|4815,4820|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|General Exam|4824,4836|false|false|false|||auscultation
Procedure|Diagnostic Procedure|General Exam|4824,4836|false|false|false|C0004339|Auscultation|auscultation
Event|Event|General Exam|4853,4860|true|false|false|||wheezes
Finding|Sign or Symptom|General Exam|4853,4860|true|false|false|C0043144|Wheezing|wheezes
Event|Event|General Exam|4862,4869|true|false|false|||rhonchi
Finding|Finding|General Exam|4862,4869|true|false|false|C0035508|Rhonchi|rhonchi
Event|Event|General Exam|4873,4878|true|false|false|||rales
Finding|Finding|General Exam|4873,4878|true|false|false|C0034642;C0240859|Basilar Rales;Rales|rales
Event|Event|General Exam|4883,4892|true|false|false|||increased
Finding|Finding|General Exam|4883,4892|true|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Functional Concept|General Exam|4883,4892|true|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Sign or Symptom|General Exam|4883,4910|true|false|false|C0859927|Increased work of breathing|increased work of breathing
Event|Event|General Exam|4893,4897|true|false|false|||work
Event|Occupational Activity|General Exam|4893,4897|true|false|false|C0043227|Work|work
Finding|Organ or Tissue Function|General Exam|4893,4910|true|false|false|C0043229|Work of Breathing|work of breathing
Attribute|Clinical Attribute|General Exam|4901,4910|true|false|false|C5885990||breathing
Event|Event|General Exam|4901,4910|true|false|false|||breathing
Finding|Finding|General Exam|4901,4910|true|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|General Exam|4901,4910|true|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|General Exam|4901,4910|true|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|General Exam|4901,4910|true|false|false|C1160636|respiratory system process|breathing
Anatomy|Body Location or Region|General Exam|4912,4919|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|General Exam|4912,4919|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|General Exam|4912,4919|false|false|false|||ABDOMEN
Finding|Finding|General Exam|4912,4919|false|false|false|C0941288|Abdomen problem|ABDOMEN
Anatomy|Body Part, Organ, or Organ Component|General Exam|4928,4934|false|false|false|C0021853|Intestines|bowels
Event|Event|General Exam|4935,4941|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|General Exam|4935,4941|false|false|false|C0037709||sounds
Event|Event|General Exam|4947,4956|false|false|false|||distended
Finding|Finding|General Exam|4947,4956|false|false|false|C0700124|Dilated|distended
Attribute|Clinical Attribute|General Exam|4972,4976|false|false|false|C4318566|Deep Resection Margin|deep
Event|Event|General Exam|4977,4986|false|false|false|||palpation
Procedure|Diagnostic Procedure|General Exam|4977,4986|false|false|false|C0030247|Palpation|palpation
Anatomy|Body Part, Organ, or Organ Component|General Exam|5010,5021|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Disorder|Anatomical Abnormality|General Exam|5026,5034|true|false|false|C0149651|Clubbing|clubbing
Event|Event|General Exam|5026,5034|true|false|false|||clubbing
Event|Event|General Exam|5036,5044|true|false|false|||cyanosis
Finding|Sign or Symptom|General Exam|5036,5044|true|false|false|C0010520|Cyanosis|cyanosis
Attribute|Clinical Attribute|General Exam|5049,5054|true|false|false|C1717255||edema
Event|Event|General Exam|5049,5054|true|false|false|||edema
Finding|Pathologic Function|General Exam|5049,5054|true|false|false|C0013604|Edema|edema
Drug|Food|General Exam|5056,5062|false|false|false|C5890763||Pulses
Event|Event|General Exam|5056,5062|false|false|false|||Pulses
Finding|Physiologic Function|General Exam|5056,5062|false|false|false|C0391850|Physiologic pulse|Pulses
Procedure|Health Care Activity|General Exam|5056,5062|false|false|false|C0034107|Pulse taking|Pulses
Event|Event|General Exam|5063,5065|false|false|false|||DP
Finding|Conceptual Entity|General Exam|5066,5072|false|false|false|C0442038;C0920847|Circumpennate;Radial|Radial
Anatomy|Body System|General Exam|5090,5094|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|General Exam|5090,5094|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|General Exam|5090,5094|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|General Exam|5090,5094|false|false|false|||SKIN
Finding|Body Substance|General Exam|5090,5094|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|General Exam|5090,5094|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Event|Event|General Exam|5096,5100|false|false|false|||Warm
Finding|Finding|General Exam|5096,5100|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|5096,5100|false|false|false|C0687712|warming process|Warm
Event|Event|General Exam|5102,5112|false|false|false|||NEUROLOGIC
Event|Event|General Exam|5114,5118|false|false|false|||AOx3
Finding|Gene or Genome|General Exam|5120,5123|false|false|false|C1539110|CNDP2 gene|CN2
Event|Event|General Exam|5127,5133|false|false|false|||intact
Finding|Finding|General Exam|5127,5133|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Finding|General Exam|5152,5166|false|false|false|C0026826|Muscle Hypertonia|Increased tone
Event|Event|General Exam|5162,5166|false|false|false|||tone
Anatomy|Body Part, Organ, or Organ Component|General Exam|5170,5173|false|false|false|C0227192|Inferior esophageal sphincter structure|LEs
Finding|Classification|General Exam|5170,5173|false|false|false|C0023595|Lewis Blood-Group System|LEs
Finding|Idea or Concept|General Exam|5179,5187|false|false|false|C0808080|Strength (attribute)|strength
Event|Event|General Exam|5204,5213|false|false|false|||sensation
Finding|Finding|General Exam|5204,5213|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|General Exam|5204,5213|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|General Exam|5204,5213|false|false|false|C2229507|sensory exam|sensation
Procedure|Health Care Activity|General Exam|5237,5246|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|General Exam|5247,5251|false|false|false|||LABS
Lab|Laboratory or Test Result|General Exam|5247,5251|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|General Exam|5281,5286|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|5281,5286|false|false|false|||BLOOD
Finding|Body Substance|General Exam|5281,5286|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|5287,5290|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|5295,5298|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|5295,5298|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|5295,5298|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|5305,5308|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|5305,5308|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|5305,5308|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|5305,5308|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|5315,5318|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|5315,5318|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|5326,5329|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|5326,5329|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|5326,5329|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|5326,5329|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|5326,5329|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|5333,5336|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|5333,5336|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|5333,5336|false|false|false|||MCH
Finding|Gene or Genome|General Exam|5333,5336|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|5333,5336|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|5333,5336|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|5342,5346|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|5342,5346|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|5372,5375|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|5392,5397|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|5392,5397|false|false|false|||BLOOD
Finding|Body Substance|General Exam|5392,5397|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Antibiotic|General Exam|5413,5418|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|General Exam|5413,5418|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|General Exam|5413,5418|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|General Exam|5426,5429|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Event|Event|General Exam|5426,5429|false|false|false|||Eos
Finding|Gene or Genome|General Exam|5426,5429|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|General Exam|5528,5533|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|5528,5533|false|false|false|||BLOOD
Finding|Body Substance|General Exam|5528,5533|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|5538,5541|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|General Exam|5538,5541|false|false|false|||PTT
Procedure|Laboratory Procedure|General Exam|5538,5541|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|General Exam|5564,5569|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|5564,5569|false|false|false|||BLOOD
Finding|Body Substance|General Exam|5564,5569|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|5564,5577|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|5564,5577|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|5564,5577|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|5570,5577|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|5570,5577|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|5570,5577|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|5570,5577|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|5570,5577|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|5570,5577|false|false|false|C0337438|Glucose measurement|Glucose
Event|Event|General Exam|5612,5613|false|false|false|||5
Drug|Inorganic Chemical|General Exam|5623,5627|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|5623,5627|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|5623,5627|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|5653,5658|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|5653,5658|false|false|false|||BLOOD
Finding|Body Substance|General Exam|5653,5658|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|5659,5662|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|5659,5662|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|General Exam|5659,5662|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|General Exam|5659,5662|false|false|false|||ALT
Finding|Gene or Genome|General Exam|5659,5662|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|General Exam|5659,5662|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|General Exam|5659,5662|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|General Exam|5659,5662|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|General Exam|5666,5669|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|General Exam|5666,5669|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|5666,5669|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|General Exam|5666,5669|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|General Exam|5666,5669|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|General Exam|5666,5669|false|false|false|||AST
Finding|Gene or Genome|General Exam|5666,5669|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|5673,5680|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|General Exam|5673,5680|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|General Exam|5709,5714|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|5709,5714|false|false|false|||BLOOD
Finding|Body Substance|General Exam|5709,5714|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|5715,5721|false|false|false|C0023764|lipase|Lipase
Drug|Enzyme|General Exam|5715,5721|false|false|false|C0023764|lipase|Lipase
Drug|Pharmacologic Substance|General Exam|5715,5721|false|false|false|C0023764|lipase|Lipase
Event|Event|General Exam|5715,5721|false|false|false|||Lipase
Procedure|Laboratory Procedure|General Exam|5715,5721|false|false|false|C0373670|Lipase measurement|Lipase
Disorder|Disease or Syndrome|General Exam|5737,5742|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|5737,5742|false|false|false|||BLOOD
Finding|Body Substance|General Exam|5737,5742|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|General Exam|5769,5774|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|5769,5774|false|false|false|||BLOOD
Finding|Body Substance|General Exam|5769,5774|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|5769,5782|false|false|false|C0853248|Blood albumin|BLOOD Albumin
Drug|Amino Acid, Peptide, or Protein|General Exam|5775,5782|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Biologically Active Substance|General Exam|5775,5782|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Pharmacologic Substance|General Exam|5775,5782|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Event|Event|General Exam|5775,5782|false|false|false|||Albumin
Finding|Gene or Genome|General Exam|5775,5782|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Finding|Physiologic Function|General Exam|5775,5782|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Procedure|Laboratory Procedure|General Exam|5775,5782|false|false|false|C0201838|Albumin measurement|Albumin
Drug|Biologically Active Substance|General Exam|5787,5794|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|5787,5794|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|5787,5794|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|5787,5794|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|5787,5794|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|General Exam|5787,5794|false|false|false|||Calcium
Finding|Physiologic Function|General Exam|5787,5794|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|5787,5794|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|General Exam|5827,5832|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|5827,5832|false|false|false|||BLOOD
Finding|Body Substance|General Exam|5827,5832|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|General Exam|5856,5861|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|5856,5861|false|false|false|||BLOOD
Finding|Body Substance|General Exam|5856,5861|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Attribute|Clinical Attribute|General Exam|5862,5865|false|false|false|C2708739||TSH
Drug|Amino Acid, Peptide, or Protein|General Exam|5862,5865|false|false|false|C0040160|thyrotropin|TSH
Drug|Hormone|General Exam|5862,5865|false|false|false|C0040160|thyrotropin|TSH
Drug|Pharmacologic Substance|General Exam|5862,5865|false|false|false|C0040160|thyrotropin|TSH
Event|Event|General Exam|5862,5865|false|false|false|||TSH
Procedure|Laboratory Procedure|General Exam|5862,5865|false|false|false|C0202230|Thyroid stimulating hormone measurement|TSH
Disorder|Disease or Syndrome|General Exam|5882,5887|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|5882,5887|false|false|false|||BLOOD
Finding|Body Substance|General Exam|5882,5887|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Event|General Exam|5896,5899|false|false|false|||NEG
Finding|Finding|General Exam|5896,5899|false|false|false|C5848551|Neg - answer|NEG
Disorder|Disease or Syndrome|General Exam|5912,5917|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|5912,5917|false|false|false|||BLOOD
Finding|Body Substance|General Exam|5912,5917|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|5918,5921|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Enzyme|General Exam|5918,5921|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Organic Chemical|General Exam|5918,5921|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Pharmacologic Substance|General Exam|5918,5921|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Event|Event|General Exam|5918,5921|false|false|false|||ASA
Finding|Gene or Genome|General Exam|5918,5921|false|false|false|C1412553|ARSA gene|ASA
Event|Event|General Exam|5922,5925|false|false|false|||NEG
Finding|Finding|General Exam|5922,5925|false|false|false|C5848551|Neg - answer|NEG
Disorder|Injury or Poisoning|General Exam|5926,5933|false|false|false|C0161679|Toxic effect of ethyl alcohol|Ethanol
Drug|Organic Chemical|General Exam|5926,5933|false|false|false|C0001962;C3854029;C3854030|CNS depressants ethanol;antiseptics ethanol;ethanol|Ethanol
Drug|Pharmacologic Substance|General Exam|5926,5933|false|false|false|C0001962;C3854029;C3854030|CNS depressants ethanol;antiseptics ethanol;ethanol|Ethanol
Event|Event|General Exam|5926,5933|false|false|false|||Ethanol
Procedure|Laboratory Procedure|General Exam|5926,5933|false|false|false|C0202304|Ethanol measurement|Ethanol
Event|Event|General Exam|5934,5937|false|false|false|||NEG
Finding|Finding|General Exam|5934,5937|false|false|false|C5848551|Neg - answer|NEG
Event|Event|General Exam|5946,5949|false|false|false|||NEG
Finding|Finding|General Exam|5946,5949|false|false|false|C5848551|Neg - answer|NEG
Event|Event|General Exam|5959,5962|false|false|false|||NEG
Finding|Finding|General Exam|5959,5962|false|false|false|C5848551|Neg - answer|NEG
Event|Event|General Exam|5964,5971|false|false|false|||IMAGING
Finding|Finding|General Exam|5964,5971|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|General Exam|5964,5971|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Finding|Finding|General Exam|5986,5993|false|false|false|C0740845|Imaging problem|Imaging
Procedure|Diagnostic Procedure|General Exam|5986,5993|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|Imaging
Attribute|Clinical Attribute|General Exam|5994,6001|false|false|false|C0881943||CT HEAD
Procedure|Diagnostic Procedure|General Exam|5994,6001|false|false|false|C0202691|CAT scan of head|CT HEAD
Anatomy|Body Location or Region|General Exam|5997,6001|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|HEAD
Anatomy|Body Part, Organ, or Organ Component|General Exam|5997,6001|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|HEAD
Disorder|Disease or Syndrome|General Exam|5997,6001|false|false|false|C0362076|Problems with head|HEAD
Event|Event|General Exam|5997,6001|false|false|false|||HEAD
Procedure|Therapeutic or Preventive Procedure|General Exam|5997,6001|false|false|false|C0876917|Procedure on head|HEAD
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|6006,6014|false|false|false|C0009924|Contrast Media|CONTRAST
Event|Event|Findings|6041,6049|true|false|false|||evidence
Finding|Idea or Concept|Findings|6041,6049|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Findings|6041,6052|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Event|Event|Findings|6053,6063|true|false|false|||infarction
Finding|Pathologic Function|Findings|6053,6063|true|false|false|C0021308|Infarction|infarction
Event|Event|Findings|6065,6075|true|false|false|||hemorrhage
Finding|Pathologic Function|Findings|6065,6075|true|false|false|C0019080|Hemorrhage|hemorrhage
Attribute|Clinical Attribute|Findings|6077,6082|true|false|false|C1717255||edema
Event|Event|Findings|6077,6082|true|false|false|||edema
Finding|Pathologic Function|Findings|6077,6082|true|false|false|C0013604|Edema|edema
Event|Event|Findings|6087,6091|false|false|false|||mass
Finding|Finding|Findings|6087,6091|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|Findings|6087,6091|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Findings|6087,6091|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Event|Event|Findings|6105,6115|false|false|false|||prominence
Anatomy|Body Part, Organ, or Organ Component|Findings|6123,6133|false|false|false|C0018827|Heart Ventricle|ventricles
Event|Event|Findings|6144,6154|false|false|false|||suggestive
Finding|Functional Concept|Findings|6144,6154|false|false|false|C0332299|Suggestive of|suggestive
Finding|Functional Concept|Findings|6144,6157|false|false|false|C0332299|Suggestive of|suggestive of
Event|Event|Findings|6172,6179|false|false|false|||changes
Finding|Functional Concept|Findings|6172,6179|false|false|false|C0392747|Changing|changes
Event|Event|Findings|6194,6202|true|false|false|||evidence
Finding|Idea or Concept|Findings|6194,6202|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Findings|6194,6205|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Injury or Poisoning|Findings|6206,6214|true|false|false|C0016658|Fracture|fracture
Event|Event|Findings|6206,6214|true|false|false|||fracture
Anatomy|Body Space or Junction|Findings|6259,6276|false|false|false|C0030471|Nasal sinus|paranasal sinuses
Anatomy|Body Space or Junction|Findings|6269,6276|false|false|false|C0030471;C4071871|Head>Sinuses;Nasal sinus|sinuses
Disorder|Anatomical Abnormality|Findings|6269,6276|false|false|false|C0016169|pathologic fistula|sinuses
Event|Event|Findings|6269,6276|false|false|false|||sinuses
Finding|Intellectual Product|Findings|6281,6287|false|false|false|C1552826|Table Cell Vertical Align - middle|middle
Anatomy|Body Space or Junction|Findings|6281,6291|false|false|false|C0013455|middle ear|middle ear
Disorder|Disease or Syndrome|Findings|6281,6291|false|false|false|C0271428;C0496788|Disorder of middle ear;Malignant neoplasm of middle ear|middle ear
Disorder|Neoplastic Process|Findings|6281,6291|false|false|false|C0271428;C0496788|Disorder of middle ear;Malignant neoplasm of middle ear|middle ear
Procedure|Health Care Activity|Findings|6281,6291|false|false|false|C2228461|examination of middle ear|middle ear
Anatomy|Body Part, Organ, or Organ Component|Findings|6288,6291|false|false|false|C0013443;C0521421|Ear structure|ear
Disorder|Disease or Syndrome|Findings|6288,6291|false|false|false|C0851354|Ear and labyrinth disorders|ear
Finding|Body Substance|Findings|6288,6291|false|false|false|C1546608;C1550629|SpecimenType - Ear|ear
Finding|Intellectual Product|Findings|6288,6291|false|false|false|C1546608;C1550629|SpecimenType - Ear|ear
Anatomy|Body Space or Junction|Findings|6292,6300|false|false|false|C0333343|Body cavities|cavities
Disorder|Anatomical Abnormality|Findings|6292,6300|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavities
Disorder|Disease or Syndrome|Findings|6292,6300|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavities
Event|Event|Findings|6292,6300|false|false|false|||cavities
Event|Event|Findings|6305,6310|false|false|false|||clear
Finding|Idea or Concept|Findings|6305,6310|false|false|false|C1550016|Remote control command - Clear|clear
Event|Event|Findings|6318,6328|false|false|false|||visualized
Anatomy|Body Space or Junction|Findings|6344,6350|false|false|false|C0029180|Ocular orbit|orbits
Event|Event|Findings|6355,6367|false|false|false|||unremarkable
Anatomy|Body Part, Organ, or Organ Component|Findings|6390,6394|false|false|false|C0023317|Lens, Crystalline|lens
Disorder|Disease or Syndrome|Findings|6390,6394|false|false|false|C0023308|Lens Diseases|lens
Event|Event|Findings|6390,6394|false|false|false|||lens
Procedure|Health Care Activity|Findings|6390,6394|false|false|false|C2239142|examination of lens|lens
Event|Event|Findings|6395,6407|false|false|false|||replacements
Procedure|Therapeutic or Preventive Procedure|Findings|6395,6407|false|false|false|C0035139|Surgical Replantation|replacements
Finding|Intellectual Product|Impression|6429,6434|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Location or Region|Impression|6435,6447|true|false|false|C0524466|Intracranial|intracranial
Finding|Functional Concept|Impression|6435,6447|true|false|false|C1522213|Intracranial Route of Administration|intracranial
Disorder|Congenital Abnormality|Impression|6448,6459|true|false|false|C0000768|Congenital Abnormality|abnormality
Event|Event|Impression|6448,6459|true|false|false|||abnormality
Finding|Finding|Impression|6448,6459|true|false|false|C1704258|Abnormality|abnormality
Disorder|Disease or Syndrome|Impression|6465,6478|true|false|false|C0020255|Hydrocephalus|hydrocephalus
Event|Event|Impression|6465,6478|true|false|false|||hydrocephalus
Event|Event|Impression|6486,6493|false|false|false|||Imaging
Finding|Finding|Impression|6486,6493|false|false|false|C0740845|Imaging problem|Imaging
Procedure|Diagnostic Procedure|Impression|6486,6493|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|Imaging
Anatomy|Body Location or Region|Impression|6494,6499|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|CHEST
Finding|Finding|Impression|6494,6499|false|false|false|C0741025|Chest problem|CHEST
Drug|Amino Acid, Peptide, or Protein|Impression|6506,6509|false|false|false|C1366678;C1433371;C4049852|L-Type Amino Acid Transporter;LAT protein, human;ORC3 protein, human|LAT
Drug|Biologically Active Substance|Impression|6506,6509|false|false|false|C1366678;C1433371;C4049852|L-Type Amino Acid Transporter;LAT protein, human;ORC3 protein, human|LAT
Drug|Immunologic Factor|Impression|6506,6509|false|false|false|C1366678;C1433371;C4049852|L-Type Amino Acid Transporter;LAT protein, human;ORC3 protein, human|LAT
Event|Event|Impression|6506,6509|false|false|false|||LAT
Finding|Gene or Genome|Impression|6506,6509|false|false|false|C1335085;C1425844;C1705279;C2240043|LAT gene;ORC3 gene;ORC3 wt Allele;SPNS1 gene|LAT
Finding|Intellectual Product|Impression|6526,6530|true|false|false|C1547225|Mild Severity of Illness Code|Mild
Event|Event|Impression|6531,6542|true|false|false|||atelectasis
Finding|Pathologic Function|Impression|6531,6542|true|false|false|C0004144|Atelectasis|atelectasis
Anatomy|Body Location or Region|Impression|6550,6554|true|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Impression|6550,6554|true|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Impression|6550,6554|true|false|false|C0024115|Lung diseases|lung
Finding|Finding|Impression|6550,6554|true|false|false|C0740941|Lung Problem|lung
Drug|Chemical Viewed Functionally|Impression|6555,6560|true|false|false|C0178499|Base|bases
Event|Event|Impression|6555,6560|true|false|false|||bases
Disorder|Disease or Syndrome|Impression|6575,6588|true|false|false|C0521530|Lung consolidation|consolidation
Event|Event|Impression|6575,6588|true|false|false|||consolidation
Attribute|Clinical Attribute|Impression|6593,6596|false|false|false|C1114365||Age
Drug|Biologically Active Substance|Impression|6593,6596|false|false|false|C0162574|Glycation End Products, Advanced|Age
Drug|Organic Chemical|Impression|6593,6596|false|false|false|C0162574|Glycation End Products, Advanced|Age
Event|Event|Impression|6611,6619|false|false|false|||moderate
Finding|Finding|Impression|6611,6619|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|Impression|6611,6619|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Finding|Impression|6623,6629|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Impression|6623,6629|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Event|Event|Impression|6630,6641|false|false|false|||compression
Finding|Functional Concept|Impression|6630,6641|false|false|false|C0332459;C4551657|Compressed structure|compression
Phenomenon|Natural Phenomenon or Process|Impression|6630,6641|false|false|false|C0728907|Compression|compression
Procedure|Machine Activity|Impression|6630,6641|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Procedure|Therapeutic or Preventive Procedure|Impression|6630,6641|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Disorder|Anatomical Abnormality|Impression|6642,6651|false|false|false|C0000768;C0302142|Congenital Abnormality;Deformity|deformity
Disorder|Congenital Abnormality|Impression|6642,6651|false|false|false|C0000768;C0302142|Congenital Abnormality;Deformity|deformity
Event|Event|Impression|6642,6651|false|false|false|||deformity
Finding|Finding|Impression|6642,6651|false|false|false|C2117111||deformity
Finding|Finding|Impression|6658,6661|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Impression|6658,6661|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Anatomy|Body Location or Region|Impression|6662,6670|false|false|false|C0817096|Chest|thoracic
Disorder|Disease or Syndrome|Impression|6662,6670|false|false|false|C5779551|Dissecting Thoracic Aortic Aneurysm|thoracic
Anatomy|Body Part, Organ, or Organ Component|Impression|6662,6685|false|false|false|C0223199;C1305451|Structure of body of thoracic vertebra|thoracic vertebral body
Anatomy|Body Part, Organ, or Organ Component|Impression|6671,6680|false|false|false|C0549207|Bone structure of spine|vertebral
Anatomy|Body Part, Organ, or Organ Component|Impression|6671,6685|false|false|false|C0223084|Body of vertebra|vertebral body
Anatomy|Anatomical Structure|Impression|6681,6685|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Anatomy|Body Part, Organ, or Organ Component|Impression|6681,6685|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Finding|Intellectual Product|Impression|6681,6685|false|false|false|C1551342|Document Body|body
Finding|Body Substance|Impression|6689,6698|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|Impression|6689,6698|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|Impression|6689,6698|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|Impression|6689,6698|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|Impression|6699,6703|false|false|false|||LABS
Lab|Laboratory or Test Result|Impression|6699,6703|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|Impression|6733,6738|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Impression|6733,6738|false|false|false|||BLOOD
Finding|Body Substance|Impression|6733,6738|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|Impression|6739,6742|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|Impression|6747,6750|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|Impression|6747,6750|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|Impression|6747,6750|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|Impression|6757,6760|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Impression|6757,6760|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|Impression|6757,6760|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Impression|6757,6760|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|Impression|6767,6770|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|Impression|6767,6770|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|Impression|6778,6781|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|Impression|6778,6781|false|false|false|||MCV
Lab|Laboratory or Test Result|Impression|6778,6781|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|Impression|6778,6781|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|Impression|6778,6781|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|Impression|6785,6788|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|Impression|6785,6788|false|false|false|C0600370|methacholine|MCH
Event|Event|Impression|6785,6788|false|false|false|||MCH
Finding|Gene or Genome|Impression|6785,6788|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|Impression|6785,6788|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|Impression|6785,6788|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|Impression|6795,6799|false|false|false|||MCHC
Procedure|Laboratory Procedure|Impression|6795,6799|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|Impression|6825,6828|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|Impression|6845,6850|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Impression|6845,6850|false|false|false|||BLOOD
Finding|Body Substance|Impression|6845,6850|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|Impression|6845,6858|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|Impression|6845,6858|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|Impression|6845,6858|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|Impression|6851,6858|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|Impression|6851,6858|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|Impression|6851,6858|false|false|false|C0017725|glucose|Glucose
Event|Event|Impression|6851,6858|false|false|false|||Glucose
Lab|Laboratory or Test Result|Impression|6851,6858|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|Impression|6851,6858|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|Impression|6902,6906|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|Impression|6902,6906|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|Impression|6902,6906|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|Impression|6931,6936|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Impression|6931,6936|false|false|false|||BLOOD
Finding|Body Substance|Impression|6931,6936|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|Impression|6931,6944|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|Impression|6937,6944|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|Impression|6937,6944|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|Impression|6937,6944|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|Impression|6937,6944|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|Impression|6937,6944|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|Impression|6937,6944|false|false|false|||Calcium
Finding|Physiologic Function|Impression|6937,6944|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|Impression|6937,6944|false|false|false|C0201925|Calcium measurement|Calcium
Finding|Finding|Impression|6967,6971|false|false|false|C1706180|Male Gender|male
Disorder|Disease or Syndrome|Impression|6981,6988|false|false|false|C0012634|Disease|disease
Event|Event|Impression|6981,6988|false|false|false|||disease
Disorder|Disease or Syndrome|Impression|6990,7002|false|false|false|C0242339|Dyslipidemias|dyslipidemia
Event|Event|Impression|6990,7002|false|false|false|||dyslipidemia
Event|Event|Impression|7010,7017|false|false|false|||history
Finding|Conceptual Entity|Impression|7010,7017|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Impression|7010,7017|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Impression|7010,7017|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Impression|7010,7020|false|false|false|C0262926|Medical History|history of
Anatomy|Body Part, Organ, or Organ Component|Impression|7021,7029|false|false|false|C0033572;C4266527|Prostate;Structure of prostate (body structure)|prostate
Disorder|Disease or Syndrome|Impression|7021,7029|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|prostate
Disorder|Neoplastic Process|Impression|7021,7029|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|prostate
Disorder|Neoplastic Process|Impression|7021,7036|false|false|false|C0376358;C0600139|Malignant neoplasm of prostate;Prostate carcinoma|prostate cancer
Disorder|Neoplastic Process|Impression|7030,7036|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Impression|7030,7036|false|false|false|||cancer
Procedure|Therapeutic or Preventive Procedure|Impression|7042,7055|false|false|false|C0033573|Prostatectomy|prostatectomy
Event|Event|Impression|7065,7073|false|false|false|||referred
Event|Event|Impression|7117,7121|false|false|false|||gait
Finding|Finding|Impression|7117,7121|false|false|false|C0016928|Gait|gait
Disorder|Injury or Poisoning|Impression|7123,7128|false|false|false|C0000921|Accidental Falls|falls
Event|Event|Impression|7123,7128|false|false|false|||falls
Finding|Finding|Impression|7123,7128|false|false|false|C0085639|Falls|falls
Finding|Functional Concept|Impression|7134,7140|false|false|false|C0234621|Visual|visual
Finding|Sign or Symptom|Impression|7134,7155|false|false|false|C0233763|Hallucinations, Visual|visual hallucinations
Disorder|Mental or Behavioral Dysfunction|Impression|7141,7155|false|false|false|C0018524|Hallucinations|hallucinations
Event|Event|Impression|7141,7155|false|false|false|||hallucinations
Event|Event|Impression|7156,7166|false|false|false|||concerning
Event|Event|Impression|7171,7182|false|false|false|||progression
Finding|Functional Concept|Impression|7171,7182|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Finding|Pathologic Function|Impression|7171,7182|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Disorder|Disease or Syndrome|Impression|7190,7209|false|false|false|C0027765|nervous system disorder|neurologic disorder
Disorder|Disease or Syndrome|Impression|7201,7209|false|false|false|C0012634|Disease|disorder
Event|Event|Impression|7201,7209|false|false|false|||disorder
Finding|Intellectual Product|Impression|7213,7218|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|ACUTE
Disorder|Disease or Syndrome|Impression|7259,7266|false|false|false|C0012634|Disease|disease
Event|Event|Impression|7259,7266|false|false|false|||disease
Anatomy|Anatomical Structure|Impression|7271,7275|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|Body
Anatomy|Body Part, Organ, or Organ Component|Impression|7271,7275|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|Body
Finding|Intellectual Product|Impression|7271,7275|false|false|false|C1551342|Document Body|Body
Disorder|Mental or Behavioral Dysfunction|Impression|7276,7284|false|false|false|C0011265;C0497327|Dementia;Presenile dementia|Dementia
Event|Event|Impression|7276,7284|false|false|false|||Dementia
Finding|Functional Concept|Impression|7287,7293|false|false|false|C0234621|Visual|Visual
Finding|Sign or Symptom|Impression|7287,7308|false|false|false|C0233763|Hallucinations, Visual|Visual Hallucinations
Disorder|Mental or Behavioral Dysfunction|Impression|7294,7308|false|false|false|C0018524|Hallucinations|Hallucinations
Event|Event|Impression|7294,7308|false|false|false|||Hallucinations
Finding|Body Substance|Impression|7314,7321|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Impression|7314,7321|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Impression|7314,7321|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Impression|7338,7343|false|false|false|||acute
Finding|Intellectual Product|Impression|7338,7343|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Intellectual Product|Impression|7347,7354|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Impression|7347,7354|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Event|Event|Impression|7355,7366|false|false|false|||progression
Finding|Functional Concept|Impression|7355,7366|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Finding|Pathologic Function|Impression|7355,7366|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Disorder|Disease or Syndrome|Impression|7378,7385|false|false|false|C0012634|Disease|disease
Event|Event|Impression|7378,7385|false|false|false|||disease
Disorder|Disease or Syndrome|Impression|7406,7413|false|false|false|C0012634|Disease|disease
Event|Event|Impression|7406,7413|false|false|false|||disease
Finding|Pathologic Function|Impression|7406,7425|false|false|false|C0242656|Disease Progression|disease progression
Event|Event|Impression|7414,7425|false|false|false|||progression
Finding|Functional Concept|Impression|7414,7425|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Finding|Pathologic Function|Impression|7414,7425|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Event|Event|Impression|7429,7439|false|false|false|||underlying
Finding|Functional Concept|Impression|7440,7447|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|Impression|7440,7447|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|Impression|7440,7447|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|Impression|7440,7447|false|false|false|C0199168|Medical service|medical
Event|Event|Impression|7448,7453|false|false|false|||cause
Finding|Conceptual Entity|Impression|7448,7453|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Finding|Functional Concept|Impression|7448,7453|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Drug|Organic Chemical|Impression|7465,7472|false|false|false|C0721754|Mirapex|mirapex
Drug|Pharmacologic Substance|Impression|7465,7472|false|false|false|C0721754|Mirapex|mirapex
Event|Event|Impression|7465,7472|false|false|false|||mirapex
Drug|Organic Chemical|Impression|7474,7484|false|false|false|C0525678|rasagiline|rasagiline
Drug|Pharmacologic Substance|Impression|7474,7484|false|false|false|C0525678|rasagiline|rasagiline
Event|Event|Impression|7474,7484|false|false|false|||rasagiline
Drug|Organic Chemical|Impression|7491,7503|false|false|false|C0649350|rivastigmine|rivastigmine
Drug|Pharmacologic Substance|Impression|7491,7503|false|false|false|C0649350|rivastigmine|rivastigmine
Event|Event|Impression|7491,7503|false|false|false|||rivastigmine
Event|Event|Impression|7515,7526|false|false|false|||recommended
Event|Event|Impression|7527,7534|false|false|false|||started
Drug|Organic Chemical|Impression|7535,7543|false|false|false|C0287163|Seroquel|Seroquel
Drug|Pharmacologic Substance|Impression|7535,7543|false|false|false|C0287163|Seroquel|Seroquel
Event|Event|Impression|7535,7543|false|false|false|||Seroquel
Disorder|Mental or Behavioral Dysfunction|Impression|7553,7567|false|false|false|C0018524|Hallucinations|hallucinations
Event|Event|Impression|7553,7567|false|false|false|||hallucinations
Event|Event|Impression|7577,7586|false|false|false|||evaluated
Finding|Finding|Impression|7590,7598|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Finding|Functional Concept|Impression|7590,7598|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Procedure|Health Care Activity|Impression|7590,7598|false|false|false|C0031809|Physical Examination|physical
Finding|Intellectual Product|Impression|7590,7606|false|false|false|C1547999|Diagnostic Service Section ID - Physical Therapy|physical therapy
Procedure|Therapeutic or Preventive Procedure|Impression|7590,7606|false|false|false|C0949766|Physical therapy|physical therapy
Event|Event|Impression|7599,7606|false|false|false|||therapy
Finding|Finding|Impression|7599,7606|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|Impression|7599,7606|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|Impression|7599,7606|false|false|false|C0087111|Therapeutic procedure|therapy
Event|Event|Impression|7611,7622|false|false|false|||recommended
Event|Event|Impression|7623,7628|false|false|false|||rehab
Procedure|Therapeutic or Preventive Procedure|Impression|7623,7628|false|false|false|C0034991|Rehabilitation therapy|rehab
Event|Event|Impression|7636,7650|false|false|false|||recommendation
Finding|Idea or Concept|Impression|7636,7650|false|false|false|C0034866|Recommendation|recommendation
Event|Event|Impression|7655,7664|false|false|false|||discussed
Finding|Classification|Impression|7674,7680|false|false|true|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Impression|7674,7680|false|false|true|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Impression|7674,7680|false|false|true|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Impression|7674,7680|false|false|true|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Event|Event|Impression|7685,7690|false|false|false|||opted
Event|Event|Impression|7696,7705|false|false|false|||discharge
Finding|Body Substance|Impression|7696,7705|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Impression|7696,7705|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Impression|7696,7705|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Impression|7696,7705|false|false|false|C0030685|Patient Discharge|discharge
Procedure|Therapeutic or Preventive Procedure|Impression|7696,7713|false|false|false|C0184713|Discharge to home|discharge to home
Event|Event|Impression|7709,7713|false|false|false|||home
Finding|Idea or Concept|Impression|7709,7713|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Impression|7709,7713|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Impression|7709,7713|false|false|false|C1553498|home health encounter|home
Finding|Idea or Concept|Impression|7719,7723|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Impression|7719,7723|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Impression|7719,7723|false|false|false|C1553498|home health encounter|home
Finding|Finding|Impression|7724,7732|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Finding|Functional Concept|Impression|7724,7732|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Procedure|Health Care Activity|Impression|7724,7732|false|false|false|C0031809|Physical Examination|physical
Finding|Intellectual Product|Impression|7724,7740|false|false|false|C1547999|Diagnostic Service Section ID - Physical Therapy|physical therapy
Procedure|Therapeutic or Preventive Procedure|Impression|7724,7740|false|false|false|C0949766|Physical therapy|physical therapy
Event|Event|Impression|7733,7740|false|false|false|||therapy
Finding|Finding|Impression|7733,7740|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|Impression|7733,7740|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|Impression|7733,7740|false|false|false|C0087111|Therapeutic procedure|therapy
Drug|Biologically Active Substance|Impression|7756,7760|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Impression|7756,7760|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Substance|Impression|7756,7760|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Event|Event|Impression|7756,7760|false|false|false|||line
Finding|Intellectual Product|Impression|7756,7760|false|false|false|C1546701|line source specimen code|line
Finding|Body Substance|Impression|7771,7778|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Impression|7771,7778|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Impression|7771,7778|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Attribute|Clinical Attribute|Impression|7781,7786|false|false|false|C2979882||goals
Event|Event|Impression|7781,7786|false|false|false|||goals
Finding|Idea or Concept|Impression|7781,7786|false|false|false|C0018017;C0679840;C1546459|What subject filter - Goals;objective (goal);treatment goals|goals
Finding|Intellectual Product|Impression|7781,7786|false|false|false|C0018017;C0679840;C1546459|What subject filter - Goals;objective (goal);treatment goals|goals
Procedure|Health Care Activity|Impression|7781,7794|false|false|false|C2930505|Goals of Care|goals of care
Event|Activity|Impression|7790,7794|false|false|false|C1947933|care activity|care
Event|Event|Impression|7790,7794|false|false|false|||care
Finding|Finding|Impression|7790,7794|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Impression|7790,7794|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Idea or Concept|Impression|7797,7809|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Event|Event|Impression|7810,7816|false|false|false|||ISSUES
Event|Event|Impression|7821,7822|false|false|false|||f
Finding|Functional Concept|Impression|7825,7831|false|false|false|C0234621|Visual|visual
Finding|Sign or Symptom|Impression|7825,7845|false|false|false|C0233763|Hallucinations, Visual|visual hallucination
Disorder|Mental or Behavioral Dysfunction|Impression|7832,7845|false|false|false|C0018524|Hallucinations|hallucination
Event|Event|Impression|7832,7845|false|false|false|||hallucination
Event|Event|Impression|7846,7854|false|false|false|||symptoms
Finding|Functional Concept|Impression|7846,7854|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Impression|7846,7854|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Drug|Organic Chemical|Impression|7858,7866|false|false|false|C0287163|Seroquel|Seroquel
Drug|Pharmacologic Substance|Impression|7858,7866|false|false|false|C0287163|Seroquel|Seroquel
Event|Event|Impression|7858,7866|false|false|false|||Seroquel
Event|Event|Impression|7870,7871|false|false|false|||f
Finding|Finding|Impression|7874,7882|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Finding|Functional Concept|Impression|7874,7882|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Procedure|Health Care Activity|Impression|7874,7882|false|false|false|C0031809|Physical Examination|physical
Finding|Intellectual Product|Impression|7874,7890|false|false|false|C1547999|Diagnostic Service Section ID - Physical Therapy|physical therapy
Procedure|Therapeutic or Preventive Procedure|Impression|7874,7890|false|false|false|C0949766|Physical therapy|physical therapy
Event|Event|Impression|7883,7890|false|false|false|||therapy
Finding|Finding|Impression|7883,7890|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|Impression|7883,7890|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|Impression|7883,7890|false|false|false|C0087111|Therapeutic procedure|therapy
Finding|Finding|Impression|7891,7898|false|false|false|C4534363|At home|at home
Event|Event|Impression|7894,7898|false|false|false|||home
Finding|Idea or Concept|Impression|7894,7898|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Impression|7894,7898|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Impression|7894,7898|false|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|Impression|7901,7912|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Impression|7901,7912|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Impression|7901,7912|false|false|false|||Medications
Finding|Intellectual Product|Impression|7901,7912|false|false|false|C4284232|Medications|Medications
Finding|Finding|Impression|7901,7925|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Impression|7916,7925|false|false|false|||Admission
Procedure|Health Care Activity|Impression|7916,7925|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|Impression|7944,7954|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Impression|7944,7954|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|Impression|7944,7959|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|Impression|7955,7959|false|false|false|||list
Finding|Intellectual Product|Impression|7955,7959|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|Impression|7967,7977|false|false|false|||inaccurate
Event|Event|Impression|7982,7990|false|false|false|||requires
Event|Event|Impression|7999,8012|false|false|false|||investigation
Finding|Intellectual Product|Impression|7999,8012|false|false|false|C1552578|Act Class - investigation|investigation
Procedure|Health Care Activity|Impression|7999,8012|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|investigation
Drug|Organic Chemical|Impression|8017,8027|false|false|false|C0525678|rasagiline|Rasagiline
Drug|Pharmacologic Substance|Impression|8017,8027|false|false|false|C0525678|rasagiline|Rasagiline
Drug|Organic Chemical|Impression|8046,8057|false|false|false|C0074710|pramipexole|Pramipexole
Drug|Pharmacologic Substance|Impression|8046,8057|false|false|false|C0074710|pramipexole|Pramipexole
Event|Event|Impression|8070,8073|false|false|false|||TID
Drug|Organic Chemical|Impression|8078,8090|false|false|false|C0649350|rivastigmine|rivastigmine
Drug|Pharmacologic Substance|Impression|8078,8090|false|false|false|C0649350|rivastigmine|rivastigmine
Event|Event|Impression|8078,8090|false|false|false|||rivastigmine
Finding|Finding|Impression|8104,8115|false|false|false|C0040652;C0694643;C4521342|Transdermal (intended site);Transdermal Route of Administration;transdermal|transdermal
Finding|Functional Concept|Impression|8104,8115|false|false|false|C0040652;C0694643;C4521342|Transdermal (intended site);Transdermal Route of Administration;transdermal|transdermal
Drug|Organic Chemical|Impression|8126,8137|false|false|false|C0085542|pravastatin|Pravastatin
Drug|Pharmacologic Substance|Impression|8126,8137|false|false|false|C0085542|pravastatin|Pravastatin
Event|Event|Impression|8147,8150|false|false|false|||QPM
Drug|Organic Chemical|Impression|8155,8169|false|false|false|C0042845;C3714801|Cyanocobalamin Drug Class;vitamin B12|Cyanocobalamin
Drug|Pharmacologic Substance|Impression|8155,8169|false|false|false|C0042845;C3714801|Cyanocobalamin Drug Class;vitamin B12|Cyanocobalamin
Drug|Vitamin|Impression|8155,8169|false|false|false|C0042845;C3714801|Cyanocobalamin Drug Class;vitamin B12|Cyanocobalamin
Event|Event|Impression|8170,8174|false|false|false|||Dose
Drug|Amino Acid, Peptide, or Protein|Impression|8178,8185|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|Unknown
Drug|Immunologic Factor|Impression|8178,8185|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|Unknown
Drug|Pharmacologic Substance|Impression|8178,8185|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|Unknown
Event|Event|Impression|8178,8185|false|false|false|||Unknown
Finding|Finding|Impression|8178,8185|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|Unknown
Finding|Functional Concept|Impression|8178,8185|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|Unknown
Finding|Idea or Concept|Impression|8178,8185|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|Unknown
Finding|Intellectual Product|Impression|8178,8185|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|Unknown
Drug|Organic Chemical|Impression|8200,8210|false|false|false|C0065180|loratadine|Loratadine
Drug|Pharmacologic Substance|Impression|8200,8210|false|false|false|C0065180|loratadine|Loratadine
Event|Event|Impression|8230,8239|false|false|false|||Discharge
Finding|Body Substance|Impression|8230,8239|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Impression|8230,8239|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Impression|8230,8239|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Impression|8230,8239|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Impression|8230,8251|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Impression|8240,8251|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Impression|8240,8251|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Impression|8240,8251|false|false|false|||Medications
Finding|Intellectual Product|Impression|8240,8251|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Impression|8257,8267|false|false|false|C0123091|quetiapine|QUEtiapine
Drug|Pharmacologic Substance|Impression|8257,8267|false|false|false|C0123091|quetiapine|QUEtiapine
Event|Event|Impression|8257,8267|false|false|false|||QUEtiapine
Drug|Organic Chemical|Impression|8257,8276|false|false|false|C0724680|quetiapine fumarate|QUEtiapine Fumarate
Drug|Pharmacologic Substance|Impression|8257,8276|false|false|false|C0724680|quetiapine fumarate|QUEtiapine Fumarate
Drug|Organic Chemical|Impression|8268,8276|false|false|false|C0220833|fumarate|Fumarate
Drug|Pharmacologic Substance|Impression|8268,8276|false|false|false|C0220833|fumarate|Fumarate
Event|Event|Impression|8268,8276|false|false|false|||Fumarate
Drug|Organic Chemical|Impression|8295,8305|false|false|false|C0123091|quetiapine|quetiapine
Drug|Pharmacologic Substance|Impression|8295,8305|false|false|false|C0123091|quetiapine|quetiapine
Event|Event|Impression|8295,8305|false|false|false|||quetiapine
Drug|Biomedical or Dental Material|Impression|8314,8320|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Impression|8324,8332|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Impression|8327,8332|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Impression|8327,8332|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Biomedical or Dental Material|Impression|8353,8359|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Impression|8360,8367|false|false|false|||Refills
Finding|Idea or Concept|Impression|8360,8367|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Impression|8376,8386|false|false|false|C0065180|loratadine|Loratadine
Drug|Pharmacologic Substance|Impression|8376,8386|false|false|false|C0065180|loratadine|Loratadine
Drug|Organic Chemical|Impression|8408,8419|false|false|false|C0074710|pramipexole|Pramipexole
Drug|Pharmacologic Substance|Impression|8408,8419|false|false|false|C0074710|pramipexole|Pramipexole
Event|Event|Impression|8432,8435|false|false|false|||TID
Drug|Organic Chemical|Impression|8442,8453|false|false|false|C0085542|pravastatin|Pravastatin
Drug|Pharmacologic Substance|Impression|8442,8453|false|false|false|C0085542|pravastatin|Pravastatin
Event|Event|Impression|8463,8466|false|false|false|||QPM
Drug|Organic Chemical|Impression|8473,8483|false|false|false|C0525678|rasagiline|Rasagiline
Drug|Pharmacologic Substance|Impression|8473,8483|false|false|false|C0525678|rasagiline|Rasagiline
Drug|Organic Chemical|Impression|8504,8516|false|false|false|C0649350|rivastigmine|rivastigmine
Drug|Pharmacologic Substance|Impression|8504,8516|false|false|false|C0649350|rivastigmine|rivastigmine
Event|Event|Impression|8504,8516|false|false|false|||rivastigmine
Finding|Finding|Impression|8530,8541|false|false|false|C0040652;C0694643;C4521342|Transdermal (intended site);Transdermal Route of Administration;transdermal|transdermal
Finding|Functional Concept|Impression|8530,8541|false|false|false|C0040652;C0694643;C4521342|Transdermal (intended site);Transdermal Route of Administration;transdermal|transdermal
Event|Event|Impression|8553,8562|false|false|false|||Discharge
Finding|Body Substance|Impression|8553,8562|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Impression|8553,8562|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Impression|8553,8562|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Impression|8553,8562|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Impression|8553,8574|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Impression|8553,8574|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Impression|8563,8574|false|false|false|C2926604||Disposition
Event|Event|Impression|8563,8574|false|false|false|||Disposition
Procedure|Health Care Activity|Impression|8563,8574|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|Impression|8576,8580|false|false|false|||Home
Finding|Idea or Concept|Impression|8576,8580|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Impression|8576,8580|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Impression|8576,8580|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|Impression|8586,8593|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|Impression|8586,8593|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|Impression|8596,8604|false|false|false|||Facility
Finding|Intellectual Product|Impression|8596,8604|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|Impression|8612,8621|false|false|false|||Discharge
Finding|Body Substance|Impression|8612,8621|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Impression|8612,8621|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Impression|8612,8621|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Impression|8612,8621|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Impression|8612,8631|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Impression|8622,8631|false|false|false|C0945731||Diagnosis
Event|Event|Impression|8622,8631|false|false|false|||Diagnosis
Finding|Classification|Impression|8622,8631|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Impression|8622,8631|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Impression|8622,8631|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Mental or Behavioral Dysfunction|Impression|8637,8645|false|false|false|C0011265;C0497327|Dementia;Presenile dementia|Dementia
Event|Event|Impression|8637,8645|false|false|false|||Dementia
Finding|Mental Process|Discharge Condition|8669,8675|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|8669,8682|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|8669,8682|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|8676,8682|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|8676,8682|false|false|false|C1546481|What subject filter - Status|Status
Disorder|Mental or Behavioral Dysfunction|Discharge Condition|8684,8692|false|false|false|C0009676|Confusion|Confused
Event|Event|Discharge Condition|8684,8692|false|false|false|||Confused
Finding|Finding|Discharge Condition|8684,8692|false|false|false|C0683369;C1547301|Clouded consciousness;Precaution Code - Confused|Confused
Finding|Intellectual Product|Discharge Condition|8684,8692|false|false|false|C0683369;C1547301|Clouded consciousness;Precaution Code - Confused|Confused
Event|Event|Discharge Condition|8706,8711|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|8706,8728|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|8706,8728|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|8715,8728|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|8715,8728|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|8715,8728|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|8730,8735|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|8730,8735|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|8730,8735|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|8730,8735|false|false|false|||Alert
Finding|Finding|Discharge Condition|8730,8735|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|8730,8735|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|8730,8735|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|8740,8751|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|8740,8751|false|false|false|C1704675|Interaction|interactive
Finding|Gene or Genome|Discharge Instructions|8780,8784|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|Discharge Instructions|8805,8814|false|false|false|||privilege
Finding|Conceptual Entity|Discharge Instructions|8805,8814|false|false|false|C1547898;C1706335;C1706336|Privilege;Role Privilege;User Privilege|privilege
Finding|Idea or Concept|Discharge Instructions|8805,8814|false|false|false|C1547898;C1706335;C1706336|Privilege;Role Privilege;User Privilege|privilege
Event|Event|Discharge Instructions|8815,8821|false|false|false|||caring
Event|Event|Discharge Instructions|8844,8847|false|false|false|||WAS
Event|Event|Discharge Instructions|8857,8865|false|false|false|||HOSPITAL
Finding|Idea or Concept|Discharge Instructions|8857,8865|false|false|false|C1547192|Organization unit type - Hospital|HOSPITAL
Event|Event|Discharge Instructions|8879,8883|false|false|false|||sent
Event|Event|Discharge Instructions|8891,8900|false|false|false|||emergency
Finding|Finding|Discharge Instructions|8891,8900|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Idea or Concept|Discharge Instructions|8891,8900|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Intellectual Product|Discharge Instructions|8891,8900|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Pathologic Function|Discharge Instructions|8891,8900|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Phenomenon|Phenomenon or Process|Discharge Instructions|8891,8900|false|false|false|C0013956|Emergency Situation|emergency
Procedure|Health Care Activity|Discharge Instructions|8891,8900|false|false|false|C1553500|emergency encounter|emergency
Finding|Idea or Concept|Discharge Instructions|8891,8905|false|false|false|C1546435|Encounter Referral Source - emergency room|emergency room
Event|Event|Discharge Instructions|8935,8944|false|false|false|||concerned
Finding|Functional Concept|Discharge Instructions|8966,8972|false|false|false|C0234621|Visual|visual
Finding|Sign or Symptom|Discharge Instructions|8966,8987|false|false|false|C0233763|Hallucinations, Visual|visual hallucinations
Disorder|Mental or Behavioral Dysfunction|Discharge Instructions|8973,8987|false|false|false|C0018524|Hallucinations|hallucinations
Event|Event|Discharge Instructions|8973,8987|false|false|false|||hallucinations
Event|Event|Discharge Instructions|8990,8994|false|false|false|||WHAT
Event|Event|Discharge Instructions|9007,9009|false|false|false|||ME
Finding|Idea or Concept|Discharge Instructions|9017,9025|false|false|false|C1547192|Organization unit type - Hospital|HOSPITAL
Event|Event|Discharge Instructions|9039,9046|false|false|false|||started
Finding|Finding|Discharge Instructions|9052,9055|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Discharge Instructions|9052,9055|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Drug|Pharmacologic Substance|Discharge Instructions|9056,9066|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Discharge Instructions|9056,9066|false|false|false|||medication
Finding|Intellectual Product|Discharge Instructions|9056,9066|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Discharge Instructions|9070,9074|false|false|false|||help
Event|Event|Discharge Instructions|9075,9080|false|false|false|||treat
Event|Event|Discharge Instructions|9087,9095|false|false|false|||symptoms
Finding|Functional Concept|Discharge Instructions|9087,9095|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Discharge Instructions|9087,9095|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|Discharge Instructions|9103,9109|false|false|false|||SHOULD
Event|Event|Discharge Instructions|9133,9141|false|false|false|||HOSPITAL
Finding|Idea or Concept|Discharge Instructions|9133,9141|false|false|false|C1547192|Organization unit type - Hospital|HOSPITAL
Event|Event|Discharge Instructions|9146,9154|false|false|false|||Continue
Finding|Idea or Concept|Discharge Instructions|9146,9154|false|false|false|C0549178|Continuous|Continue
Event|Event|Discharge Instructions|9158,9162|false|false|false|||take
Drug|Pharmacologic Substance|Discharge Instructions|9172,9181|false|false|false|C0013227|Pharmaceutical Preparations|medicines
Event|Event|Discharge Instructions|9172,9181|false|false|false|||medicines
Event|Event|Discharge Instructions|9186,9190|false|false|false|||keep
Event|Activity|Discharge Instructions|9197,9209|false|false|false|C0003629|Appointments|appointments
Event|Event|Discharge Instructions|9197,9209|false|false|false|||appointments
Disorder|Disease or Syndrome|Discharge Instructions|9229,9233|false|false|false|C0339510|Vitelliform Macular Dystrophy|best
Event|Event|Discharge Instructions|9229,9233|false|false|false|||best
Finding|Gene or Genome|Discharge Instructions|9229,9233|false|false|false|C1826421;C5781213|BEST1 gene;BEST1 wt Allele|best
Procedure|Health Care Activity|Discharge Instructions|9266,9274|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|9275,9287|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|9275,9287|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|9275,9287|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

