 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|47,56|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|47,56|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|47,61|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|81,90|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|81,90|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|81,90|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|81,90|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|81,90|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|81,95|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|113,118|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|113,118|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|113,118|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|137,140|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|137,140|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|137,140|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|137,140|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|137,140|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|148,155|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|148,155|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|157,165|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|168,177|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|168,177|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|168,177|false|false|false|C0020517|Hypersensitivity|Allergies
Attribute|Clinical Attribute|SIMPLE_SEGMENT|189,198|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|189,198|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|189,198|false|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|201,223|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|209,213|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|SIMPLE_SEGMENT|209,213|false|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|SIMPLE_SEGMENT|209,223|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Event|Event|SIMPLE_SEGMENT|214,223|false|false|false|||Reactions
Event|Event|SIMPLE_SEGMENT|226,235|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|226,235|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|244,259|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|250,259|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|250,259|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|250,259|false|false|false|C5441521|Complaint (finding)|Complaint
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|278,284|false|false|false|C4255010||NSTEMI
Event|Event|SIMPLE_SEGMENT|278,284|false|false|false|||NSTEMI
Finding|Finding|SIMPLE_SEGMENT|278,284|false|false|false|C3537184||NSTEMI
Finding|Classification|SIMPLE_SEGMENT|287,292|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|293,301|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|293,301|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|305,323|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|314,323|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|314,323|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|314,323|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|314,323|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|314,323|false|false|false|C0184661|Interventional procedure|Procedure
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|327,334|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|327,334|false|false|false|C1314974|Cardiac attachment|cardiac
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|327,350|false|false|false|C0261588|Cardiac catheterisation as the cause of abnormal reaction of the patient, or of later complication, without mention of misadventure at the time of the procedure|cardiac catheterization
Finding|Intellectual Product|SIMPLE_SEGMENT|327,350|false|false|false|C1547981|Diagnostic Service Section ID - Cardiac Catheterization|cardiac catheterization
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|327,350|false|false|false|C0018795;C1548828|Cardiac Catheterization Procedures;Consent Type - Cardiac Catheterization|cardiac catheterization
Procedure|Health Care Activity|SIMPLE_SEGMENT|327,350|false|false|false|C0018795;C1548828|Cardiac Catheterization Procedures;Consent Type - Cardiac Catheterization|cardiac catheterization
Event|Event|SIMPLE_SEGMENT|335,350|false|false|false|||catheterization
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|335,350|false|false|false|C0007430|Catheterization|catheterization
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|356,359|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|356,359|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|SIMPLE_SEGMENT|356,359|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|SIMPLE_SEGMENT|356,359|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|SIMPLE_SEGMENT|356,359|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|356,359|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Event|Event|SIMPLE_SEGMENT|356,359|false|false|false|||DES
Finding|Gene or Genome|SIMPLE_SEGMENT|356,359|false|false|false|C1413980|DES gene|DES
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|371,380|false|false|false|C0001168|Complete obstruction|occlusion
Event|Event|SIMPLE_SEGMENT|371,380|false|false|false|||occlusion
Finding|Finding|SIMPLE_SEGMENT|371,380|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Functional Concept|SIMPLE_SEGMENT|371,380|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|371,380|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Pathologic Function|SIMPLE_SEGMENT|371,380|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Conceptual Entity|SIMPLE_SEGMENT|388,394|false|false|false|C0442038;C0920847|Circumpennate;Radial|radial
Event|Event|SIMPLE_SEGMENT|395,401|false|false|false|||access
Finding|Functional Concept|SIMPLE_SEGMENT|395,401|false|false|false|C1554204|Role Class - access|access
Event|Event|SIMPLE_SEGMENT|404,408|false|false|false|||IABP
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|404,408|false|false|false|C0021860|Intra-Aortic Balloon Pumping|IABP
Event|Event|SIMPLE_SEGMENT|409,418|false|false|false|||placement
Procedure|Health Care Activity|SIMPLE_SEGMENT|409,418|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|409,418|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Event|Activity|SIMPLE_SEGMENT|423,430|false|false|false|C1883720|Removing (action)|removal
Event|Event|SIMPLE_SEGMENT|423,430|false|false|false|||removal
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|423,430|false|false|false|C0015252;C0185115;C0728940|Excision;Extraction;removal technique|removal
Event|Event|SIMPLE_SEGMENT|433,440|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|433,440|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|433,440|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|433,440|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|433,443|false|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|433,459|false|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|433,459|false|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|444,451|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|444,451|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|444,459|false|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|452,459|false|false|false|C0221423|Illness (finding)|Illness
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|485,488|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|485,488|false|false|false|||HTN
Event|Event|SIMPLE_SEGMENT|490,493|false|false|false|||HLD
Event|Event|SIMPLE_SEGMENT|495,499|false|false|false|||DMII
Event|Event|SIMPLE_SEGMENT|520,527|false|false|false|||medical
Finding|Functional Concept|SIMPLE_SEGMENT|520,527|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|SIMPLE_SEGMENT|520,527|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|SIMPLE_SEGMENT|520,527|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|520,527|false|false|false|C0199168|Medical service|medical
Event|Event|SIMPLE_SEGMENT|528,538|false|false|false|||management
Event|Occupational Activity|SIMPLE_SEGMENT|528,538|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|SIMPLE_SEGMENT|528,538|false|false|false|C0376636|Disease Management|management
Event|Event|SIMPLE_SEGMENT|543,547|false|false|false|||cath
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|543,547|false|false|false|C0007430|Catheterization|cath
Event|Event|SIMPLE_SEGMENT|548,557|false|false|false|||presented
Event|Event|SIMPLE_SEGMENT|575,586|false|false|false|||transferred
Event|Event|SIMPLE_SEGMENT|598,613|false|false|false|||catheterization
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|598,613|false|false|false|C0007430|Catheterization|catheterization
Event|Event|SIMPLE_SEGMENT|618,625|false|false|false|||concern
Finding|Idea or Concept|SIMPLE_SEGMENT|618,625|false|false|false|C2699424|Concern|concern
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|630,635|false|false|false|C1536220|ST segment elevation myocardial infarction|STEMI
Event|Event|SIMPLE_SEGMENT|630,635|false|false|false|||STEMI
Finding|Finding|SIMPLE_SEGMENT|630,635|false|false|false|C3538872|ST Elevation Myocardial Infarction by ECG Finding|STEMI
Finding|Body Substance|SIMPLE_SEGMENT|639,646|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|639,646|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|639,646|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Functional Concept|SIMPLE_SEGMENT|639,650|false|false|false|C0332310|Has patient|Patient has
Attribute|Clinical Attribute|SIMPLE_SEGMENT|665,671|false|false|false|C2926611||angina
Event|Event|SIMPLE_SEGMENT|665,671|false|false|false|||angina
Finding|Finding|SIMPLE_SEGMENT|665,671|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Finding|Sign or Symptom|SIMPLE_SEGMENT|665,671|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Finding|Sign or Symptom|SIMPLE_SEGMENT|665,676|false|false|false|C0002962|Angina Pectoris|angina pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|672,676|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|672,676|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|672,676|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|672,676|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|680,688|false|false|false|||exertion
Finding|Organism Function|SIMPLE_SEGMENT|680,688|false|false|false|C0015264|Exertion|exertion
Finding|Intellectual Product|SIMPLE_SEGMENT|708,713|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Intellectual Product|SIMPLE_SEGMENT|708,719|false|false|false|C1272517|Sudden onset (contextual qualifier) (qualifier value)|acute onset
Event|Event|SIMPLE_SEGMENT|749,757|false|false|false|||resolved
Event|Event|SIMPLE_SEGMENT|767,770|false|false|false|||NTG
Finding|Finding|SIMPLE_SEGMENT|767,770|false|false|false|C1417953;C1847730;C5575300|GLAUCOMA, NORMAL TENSION, SUSCEPTIBILITY TO;OPA1 gene;OPA1 wt Allele|NTG
Finding|Gene or Genome|SIMPLE_SEGMENT|767,770|false|false|false|C1417953;C1847730;C5575300|GLAUCOMA, NORMAL TENSION, SUSCEPTIBILITY TO;OPA1 gene;OPA1 wt Allele|NTG
Event|Event|SIMPLE_SEGMENT|776,785|false|false|false|||persisted
Finding|Functional Concept|SIMPLE_SEGMENT|805,813|false|false|false|C0332287;C1883712|Add - instruction imperative;In addition to|addition
Event|Event|SIMPLE_SEGMENT|820,828|false|false|false|||episodes
Event|Event|SIMPLE_SEGMENT|833,841|false|false|false|||diarrhea
Finding|Finding|SIMPLE_SEGMENT|833,841|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|833,841|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Event|Event|SIMPLE_SEGMENT|846,854|false|false|false|||weakness
Finding|Sign or Symptom|SIMPLE_SEGMENT|846,854|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Event|Event|SIMPLE_SEGMENT|855,862|false|false|false|||malaise
Finding|Sign or Symptom|SIMPLE_SEGMENT|855,862|false|false|false|C0231218|Malaise|malaise
Event|Event|SIMPLE_SEGMENT|886,895|false|false|false|||orthopnea
Finding|Finding|SIMPLE_SEGMENT|886,895|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|886,895|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|897,900|false|false|false|C1956415|Paroxysmal nocturnal dyspnea|PND
Event|Event|SIMPLE_SEGMENT|897,900|false|false|false|||PND
Finding|Gene or Genome|SIMPLE_SEGMENT|897,900|false|false|false|C1417807;C4552608|NPPA gene;NPPA wt Allele|PND
Attribute|Clinical Attribute|SIMPLE_SEGMENT|906,911|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|906,911|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|906,911|false|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|913,925|false|false|false|||palpitations
Finding|Finding|SIMPLE_SEGMENT|913,925|false|false|false|C0030252|Palpitations|palpitations
Event|Event|SIMPLE_SEGMENT|930,933|false|false|false|||SOB
Finding|Sign or Symptom|SIMPLE_SEGMENT|930,933|false|false|false|C0013404|Dyspnea|SOB
Finding|Idea or Concept|SIMPLE_SEGMENT|948,955|false|false|false|C1555582|Initial (abbreviation)|initial
Event|Event|SIMPLE_SEGMENT|956,962|false|false|false|||vitals
Event|Event|SIMPLE_SEGMENT|971,975|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|971,975|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|971,975|false|false|false|C0582103|Medical Examination|Exam
Anatomy|Body Location or Region|SIMPLE_SEGMENT|977,982|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|SIMPLE_SEGMENT|977,982|false|false|false|C0741025|Chest problem|Chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|977,987|false|false|false|C2926613||Chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|977,987|false|false|false|C0008031|Chest Pain|Chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|983,987|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|983,987|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|983,987|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|983,987|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|1005,1009|false|false|false|||Labs
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1005,1009|false|false|false|C0587081|Laboratory test finding|Labs
Anatomy|Cell|SIMPLE_SEGMENT|1024,1027|false|false|false|C0023516|Leukocytes|WBC
Event|Event|SIMPLE_SEGMENT|1034,1037|false|false|false|||Hct
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1034,1037|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1034,1037|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Event|Event|SIMPLE_SEGMENT|1044,1047|false|false|false|||Plt
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1044,1047|false|false|false|C0201617|Primed lymphocyte test|Plt
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1053,1056|false|false|false|C0368980|Coagulation tissue factor induced.INR|INR
Event|Event|SIMPLE_SEGMENT|1053,1056|false|false|false|||INR
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1053,1056|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1053,1056|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1080,1083|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Drug|Inorganic Chemical|SIMPLE_SEGMENT|1080,1083|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Event|Event|SIMPLE_SEGMENT|1080,1083|false|false|false|||BUN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1080,1083|false|false|false|C0005845|Blood urea nitrogen measurement|BUN
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1087,1090|false|false|false|C0056182;C1721462|CR1 protein, human;Complement 3b Receptor|Cr1
Drug|Immunologic Factor|SIMPLE_SEGMENT|1087,1090|false|false|false|C0056182;C1721462|CR1 protein, human;Complement 3b Receptor|Cr1
Event|Event|SIMPLE_SEGMENT|1087,1090|false|false|false|||Cr1
Finding|Gene or Genome|SIMPLE_SEGMENT|1087,1090|false|false|false|C0056182;C1413694;C1721462|CR1 gene;CR1 protein, human;Complement 3b Receptor|Cr1
Finding|Receptor|SIMPLE_SEGMENT|1087,1090|false|false|false|C0056182;C1413694;C1721462|CR1 gene;CR1 protein, human;Complement 3b Receptor|Cr1
Event|Event|SIMPLE_SEGMENT|1094,1101|false|false|false|||Imaging
Finding|Finding|SIMPLE_SEGMENT|1094,1101|false|false|false|C0740845|Imaging problem|Imaging
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1094,1101|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|Imaging
Event|Event|SIMPLE_SEGMENT|1103,1106|false|false|false|||EKG
Finding|Intellectual Product|SIMPLE_SEGMENT|1103,1106|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1103,1106|false|false|false|C1623258|Electrocardiography|EKG
Event|Event|SIMPLE_SEGMENT|1107,1113|false|false|false|||showed
Event|Event|SIMPLE_SEGMENT|1117,1127|false|false|false|||elevations
Event|Event|SIMPLE_SEGMENT|1142,1152|false|false|false|||borderline
Event|Event|SIMPLE_SEGMENT|1154,1163|false|false|false|||elevation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1154,1163|false|false|false|C0439775|Elevation procedure|elevation
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1196,1207|false|false|false|C0011570|Mental Depression|depressions
Event|Event|SIMPLE_SEGMENT|1196,1207|false|false|false|||depressions
Event|Event|SIMPLE_SEGMENT|1218,1222|false|false|false|||ECHO
Procedure|Health Care Activity|SIMPLE_SEGMENT|1218,1222|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1218,1222|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1233,1244|false|false|false|C1980023|Wall motion|wall motion
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|1238,1244|false|false|false|C0026597|Motion|motion
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|1245,1258|false|false|false|C0000768|Congenital Abnormality|abnormalities
Event|Event|SIMPLE_SEGMENT|1245,1258|false|false|false|||abnormalities
Finding|Functional Concept|SIMPLE_SEGMENT|1245,1258|false|false|false|C0000769|teratologic|abnormalities
Event|Event|SIMPLE_SEGMENT|1260,1263|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1260,1263|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|SIMPLE_SEGMENT|1272,1277|false|false|false|||acute
Finding|Intellectual Product|SIMPLE_SEGMENT|1272,1277|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|1279,1292|false|false|false|C0000768|Congenital Abnormality|abnormalities
Event|Event|SIMPLE_SEGMENT|1279,1292|false|false|false|||abnormalities
Finding|Functional Concept|SIMPLE_SEGMENT|1279,1292|false|false|false|C0000769|teratologic|abnormalities
Finding|Body Substance|SIMPLE_SEGMENT|1295,1302|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1295,1302|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1295,1302|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1314,1321|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Drug|Organic Chemical|SIMPLE_SEGMENT|1314,1321|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1314,1321|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1322,1325|false|false|false|C1135868|Gestational Trophoblastic Neoplasms|gtt
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1322,1325|false|false|false|C0991568|Drops - Drug Form|gtt
Event|Event|SIMPLE_SEGMENT|1322,1325|false|false|false|||gtt
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1322,1325|false|false|false|C0017741|Glucose tolerance test|gtt
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1333,1336|false|false|false|C1135868|Gestational Trophoblastic Neoplasms|gtt
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1333,1336|false|false|false|C0991568|Drops - Drug Form|gtt
Event|Event|SIMPLE_SEGMENT|1333,1336|false|false|false|||gtt
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1333,1336|false|false|false|C0017741|Glucose tolerance test|gtt
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1338,1341|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Enzyme|SIMPLE_SEGMENT|1338,1341|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Organic Chemical|SIMPLE_SEGMENT|1338,1341|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1338,1341|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Event|Event|SIMPLE_SEGMENT|1338,1341|false|false|false|||ASA
Finding|Gene or Genome|SIMPLE_SEGMENT|1338,1341|false|false|false|C1412553|ARSA gene|ASA
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|1349,1359|false|false|false|C1999375|ticagrelor|Ticagrelor
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1349,1359|false|false|false|C1999375|ticagrelor|Ticagrelor
Event|Event|SIMPLE_SEGMENT|1349,1359|false|false|false|||Ticagrelor
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1375,1380|false|false|false|C0042313|vancomycin|Vanco
Drug|Antibiotic|SIMPLE_SEGMENT|1375,1380|false|false|false|C0042313|vancomycin|Vanco
Event|Event|SIMPLE_SEGMENT|1396,1407|false|false|false|||Transferred
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1419,1426|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|1419,1426|false|false|false|C1314974|Cardiac attachment|cardiac
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1419,1431|false|false|false|C0018795|Cardiac Catheterization Procedures|cardiac cath
Event|Event|SIMPLE_SEGMENT|1427,1431|false|false|false|||cath
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1427,1431|false|false|false|C0007430|Catheterization|cath
Event|Event|SIMPLE_SEGMENT|1433,1439|false|false|false|||Vitals
Event|Event|SIMPLE_SEGMENT|1443,1451|false|false|false|||transfer
Finding|Functional Concept|SIMPLE_SEGMENT|1443,1451|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|SIMPLE_SEGMENT|1443,1451|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|SIMPLE_SEGMENT|1443,1451|false|false|false|C4706767|Transfer (immobility management)|transfer
Event|Event|SIMPLE_SEGMENT|1483,1491|false|false|false|||afebrile
Finding|Finding|SIMPLE_SEGMENT|1483,1491|false|false|false|C0277797|Apyrexial|afebrile
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1492,1496|false|false|false|C0007430|Catheterization|Cath
Event|Event|SIMPLE_SEGMENT|1497,1500|false|false|false|||lab
Finding|Gene or Genome|SIMPLE_SEGMENT|1497,1500|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|lab
Finding|Intellectual Product|SIMPLE_SEGMENT|1497,1500|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|lab
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1510,1515|false|false|false|C1410088|Still|still
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1524,1528|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|1524,1528|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1524,1528|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1524,1528|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1532,1539|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|SIMPLE_SEGMENT|1532,1539|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1532,1539|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Event|Event|SIMPLE_SEGMENT|1532,1539|false|false|false|||heparin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1550,1553|false|false|false|C1135868|Gestational Trophoblastic Neoplasms|gtt
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1550,1553|false|false|false|C0991568|Drops - Drug Form|gtt
Event|Event|SIMPLE_SEGMENT|1550,1553|false|false|false|||gtt
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1550,1553|false|false|false|C0017741|Glucose tolerance test|gtt
Event|Event|SIMPLE_SEGMENT|1556,1571|false|false|false|||Catheterization
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1556,1571|false|false|false|C0007430|Catheterization|Catheterization
Event|Event|SIMPLE_SEGMENT|1572,1578|false|false|false|||showed
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|1594,1603|false|false|false|C0001168|Complete obstruction|occlusion
Event|Event|SIMPLE_SEGMENT|1594,1603|false|false|false|||occlusion
Finding|Finding|SIMPLE_SEGMENT|1594,1603|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Functional Concept|SIMPLE_SEGMENT|1594,1603|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|1594,1603|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Pathologic Function|SIMPLE_SEGMENT|1594,1603|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1613,1620|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|1613,1620|false|false|false|||disease
Drug|Organic Chemical|SIMPLE_SEGMENT|1638,1646|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1638,1646|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|1638,1646|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|SIMPLE_SEGMENT|1638,1646|false|false|false|||complete
Finding|Functional Concept|SIMPLE_SEGMENT|1638,1646|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|1638,1646|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|1647,1656|false|false|false|C0001168|Complete obstruction|occlusion
Event|Event|SIMPLE_SEGMENT|1647,1656|false|false|false|||occlusion
Finding|Finding|SIMPLE_SEGMENT|1647,1656|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Functional Concept|SIMPLE_SEGMENT|1647,1656|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|1647,1656|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Pathologic Function|SIMPLE_SEGMENT|1647,1656|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Event|Event|SIMPLE_SEGMENT|1660,1670|false|false|false|||circumflex
Event|Event|SIMPLE_SEGMENT|1696,1704|false|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|1696,1704|false|false|false|C1261287|Stenosis|stenosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1716,1719|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1716,1719|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1716,1719|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|SIMPLE_SEGMENT|1716,1719|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|SIMPLE_SEGMENT|1716,1719|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1716,1719|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Event|Event|SIMPLE_SEGMENT|1716,1719|false|false|false|||DES
Finding|Gene or Genome|SIMPLE_SEGMENT|1716,1719|false|false|false|C1413980|DES gene|DES
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|1731,1740|false|false|false|C0001168|Complete obstruction|occlusion
Event|Event|SIMPLE_SEGMENT|1731,1740|false|false|false|||occlusion
Finding|Finding|SIMPLE_SEGMENT|1731,1740|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Functional Concept|SIMPLE_SEGMENT|1731,1740|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|1731,1740|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Pathologic Function|SIMPLE_SEGMENT|1731,1740|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Conceptual Entity|SIMPLE_SEGMENT|1748,1754|false|false|false|C0442038;C0920847|Circumpennate;Radial|radial
Event|Event|SIMPLE_SEGMENT|1755,1761|false|false|false|||access
Finding|Functional Concept|SIMPLE_SEGMENT|1755,1761|false|false|false|C1554204|Role Class - access|access
Event|Event|SIMPLE_SEGMENT|1763,1774|false|false|false|||Hypotensive
Finding|Pathologic Function|SIMPLE_SEGMENT|1763,1774|false|false|false|C0857353|Hypotensive|Hypotensive
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|1801,1804|false|false|false|C0016520|Structure of interventricular foramen|IVF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1801,1804|false|false|false|C2751898|Ventricular Fibrillation, Paroxysmal Familial, 1|IVF
Event|Event|SIMPLE_SEGMENT|1801,1804|false|false|false|||IVF
Finding|Gene or Genome|SIMPLE_SEGMENT|1801,1804|false|false|false|C1419864;C4321334|SCN5A gene;SCN5A wt Allele|IVF
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1801,1804|false|false|false|C0015915;C0872104|Assisted Reproductive Technologies;Fertilization in Vitro|IVF
Finding|Sign or Symptom|SIMPLE_SEGMENT|1807,1815|false|false|false|C0010200|Coughing|Coughing
Event|Event|SIMPLE_SEGMENT|1816,1830|false|false|false|||post-procedure
Event|Event|SIMPLE_SEGMENT|1836,1841|false|false|false|||LVEDP
Finding|Finding|SIMPLE_SEGMENT|1836,1841|false|false|false|C0456190|Left ventricular end-diastolic pressure|LVEDP
Drug|Organic Chemical|SIMPLE_SEGMENT|1854,1859|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1854,1859|false|false|false|C0699992|Lasix|Lasix
Event|Event|SIMPLE_SEGMENT|1870,1873|false|false|false|||Was
Finding|Intellectual Product|SIMPLE_SEGMENT|1874,1878|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|SIMPLE_SEGMENT|1879,1891|false|false|false|||hypertensive
Finding|Finding|SIMPLE_SEGMENT|1879,1891|false|false|false|C0857121|Hypertensive (finding)|hypertensive
Drug|Organic Chemical|SIMPLE_SEGMENT|1916,1921|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1916,1921|false|false|false|C0699992|Lasix|Lasix
Event|Event|SIMPLE_SEGMENT|1932,1940|false|false|false|||Admitted
Event|Event|SIMPLE_SEGMENT|1944,1947|false|false|false|||CCU
Event|Event|SIMPLE_SEGMENT|1952,1963|false|false|false|||hypotension
Finding|Finding|SIMPLE_SEGMENT|1952,1963|false|false|false|C0020649|Hypotension|hypotension
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1975,1984|false|false|false|C0945766||procedure
Event|Event|SIMPLE_SEGMENT|1975,1984|false|false|false|||procedure
Event|Occupational Activity|SIMPLE_SEGMENT|1975,1984|false|false|false|C1546467|Act Class - procedure|procedure
Finding|Functional Concept|SIMPLE_SEGMENT|1975,1984|false|false|false|C2700391|Procedure (set of actions)|procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1975,1984|false|false|false|C0184661|Interventional procedure|procedure
Anatomy|Cell|SIMPLE_SEGMENT|1986,1989|false|false|false|C0023516|Leukocytes|WBC
Event|Event|SIMPLE_SEGMENT|2011,2015|false|false|false|||beds
Finding|Body Substance|SIMPLE_SEGMENT|2029,2036|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|2029,2036|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|2029,2036|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|2037,2044|false|false|false|||reports
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2048,2053|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|2048,2053|true|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2048,2058|true|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2048,2058|true|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2054,2058|true|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|2054,2058|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|2054,2058|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2054,2058|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|2064,2073|false|false|false|||continues
Finding|Finding|SIMPLE_SEGMENT|2082,2098|false|false|false|C0239134|Productive Cough|productive cough
Drug|Organic Chemical|SIMPLE_SEGMENT|2093,2098|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2093,2098|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|SIMPLE_SEGMENT|2093,2098|false|false|false|||cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|2093,2098|false|false|false|C0010200|Coughing|cough
Event|Event|SIMPLE_SEGMENT|2103,2111|false|false|false|||diarrhea
Finding|Finding|SIMPLE_SEGMENT|2103,2111|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|2103,2111|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Gene or Genome|SIMPLE_SEGMENT|2133,2136|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|SIMPLE_SEGMENT|2141,2150|false|false|false|||endoscopy
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2141,2150|false|false|false|C0014245;C0079278|Endoscopy (procedure);Endoscopy, Gastrointestinal|endoscopy
Event|Event|SIMPLE_SEGMENT|2155,2164|false|false|false|||diagnosed
Drug|Antibiotic|SIMPLE_SEGMENT|2194,2208|false|false|false|C0055856|clarithromycin|clarithromycin
Drug|Organic Chemical|SIMPLE_SEGMENT|2194,2208|false|false|false|C0055856|clarithromycin|clarithromycin
Event|Event|SIMPLE_SEGMENT|2194,2208|false|false|false|||clarithromycin
Drug|Antibiotic|SIMPLE_SEGMENT|2213,2224|false|false|false|C0002645|amoxicillin|amoxicillin
Drug|Organic Chemical|SIMPLE_SEGMENT|2213,2224|false|false|false|C0002645|amoxicillin|amoxicillin
Event|Event|SIMPLE_SEGMENT|2213,2224|false|false|false|||amoxicillin
Event|Event|SIMPLE_SEGMENT|2240,2249|false|false|false|||developed
Event|Event|SIMPLE_SEGMENT|2250,2258|false|false|false|||diarrhea
Finding|Finding|SIMPLE_SEGMENT|2250,2258|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|2250,2258|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2274,2280|false|false|false|C0944911||weight
Finding|Finding|SIMPLE_SEGMENT|2274,2280|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|2274,2280|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|2274,2280|false|false|false|C1305866|Weighing patient|weight
Finding|Finding|SIMPLE_SEGMENT|2274,2285|false|false|false|C1262477;C3540682|Losing Weight (question);Weight Loss|weight loss
Finding|Intellectual Product|SIMPLE_SEGMENT|2274,2285|false|false|false|C1262477;C3540682|Losing Weight (question);Weight Loss|weight loss
Event|Event|SIMPLE_SEGMENT|2281,2285|false|false|false|||loss
Finding|Finding|SIMPLE_SEGMENT|2281,2285|false|false|false|C5890125|Loss (adaptation)|loss
Finding|Finding|SIMPLE_SEGMENT|2308,2328|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|2313,2320|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|2313,2320|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|2313,2320|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|2313,2320|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2313,2320|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|2313,2328|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2321,2328|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2321,2328|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2321,2328|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2333,2336|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|2333,2336|false|false|false|||HTN
Event|Event|SIMPLE_SEGMENT|2340,2343|false|false|false|||HLD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2355,2358|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2355,2358|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|2355,2358|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|2355,2358|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|2355,2358|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2355,2358|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|2355,2358|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2355,2358|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|SIMPLE_SEGMENT|2378,2385|false|false|false|||managed
Event|Occupational Activity|SIMPLE_SEGMENT|2378,2385|false|false|false|C1273870|Management procedure|managed
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|2402,2417|false|false|false|C0037944;C1861329|Spinal Stenosis;Spinal canal stenosis|Spinal stenosis
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|2402,2417|false|false|false|C0037944;C1861329|Spinal Stenosis;Spinal canal stenosis|Spinal stenosis
Event|Event|SIMPLE_SEGMENT|2409,2417|false|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|2409,2417|false|false|false|C1261287|Stenosis|stenosis
Finding|Functional Concept|SIMPLE_SEGMENT|2420,2426|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|2420,2434|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|2427,2434|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2427,2434|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2427,2434|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2427,2434|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|2440,2446|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2440,2446|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|2440,2446|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|2440,2446|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|2440,2454|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|2447,2454|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2447,2454|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2447,2454|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2447,2454|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2456,2462|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|SIMPLE_SEGMENT|2456,2462|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Finding|SIMPLE_SEGMENT|2464,2472|false|false|false|C0332149|Possible|possible
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2481,2495|false|true|false|C0878544|Cardiomyopathies|cardiomyopathy
Event|Event|SIMPLE_SEGMENT|2481,2495|false|false|false|||cardiomyopathy
Finding|Classification|SIMPLE_SEGMENT|2499,2505|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2499,2505|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|2499,2505|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|2499,2505|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Finding|SIMPLE_SEGMENT|2499,2513|true|false|false|C0241889|Family Medical History|family history
Finding|Finding|SIMPLE_SEGMENT|2499,2516|true|false|false|C0241889|Family Medical History|family history of
Event|Event|SIMPLE_SEGMENT|2506,2513|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|2506,2513|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2506,2513|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|2506,2513|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2506,2516|true|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2527,2537|true|false|false|C0003811|Cardiac Arrhythmia|arrhythmia
Event|Event|SIMPLE_SEGMENT|2527,2537|false|false|false|||arrhythmia
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2549,2556|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|2549,2556|false|false|false|C1314974|Cardiac attachment|cardiac
Event|Event|SIMPLE_SEGMENT|2558,2563|false|false|false|||death
Finding|Finding|SIMPLE_SEGMENT|2558,2563|false|false|false|C0011065;C1306577;C1546949|Cessation of life;Death (finding);Event Consequence - Death|death
Finding|Idea or Concept|SIMPLE_SEGMENT|2558,2563|false|false|false|C0011065;C1306577;C1546949|Cessation of life;Death (finding);Event Consequence - Death|death
Finding|Organism Function|SIMPLE_SEGMENT|2558,2563|false|false|false|C0011065;C1306577;C1546949|Cessation of life;Death (finding);Event Consequence - Death|death
Event|Event|SIMPLE_SEGMENT|2575,2591|false|false|false|||non-contributory
Event|Event|SIMPLE_SEGMENT|2597,2605|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|2597,2605|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|2597,2605|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2597,2605|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|2597,2610|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2597,2610|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|2606,2610|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|2606,2610|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2606,2610|false|false|false|C0582103|Medical Examination|Exam
Event|Event|SIMPLE_SEGMENT|2615,2624|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|2615,2624|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|2646,2654|false|false|false|||afebrile
Finding|Finding|SIMPLE_SEGMENT|2646,2654|false|false|false|C0277797|Apyrexial|afebrile
Event|Event|SIMPLE_SEGMENT|2680,2694|false|false|false|||Non-rebreather
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2695,2701|false|false|false|C0944911||Weight
Event|Event|SIMPLE_SEGMENT|2695,2701|false|false|false|||Weight
Finding|Finding|SIMPLE_SEGMENT|2695,2701|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|Weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|2695,2701|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|Weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|2695,2701|false|false|false|C1305866|Weighing patient|Weight
Event|Event|SIMPLE_SEGMENT|2708,2712|false|false|false|||Tele
Finding|Gene or Genome|SIMPLE_SEGMENT|2708,2712|false|false|false|C1420621;C1515258|TCAP gene;Telephone Number|Tele
Finding|Intellectual Product|SIMPLE_SEGMENT|2708,2712|false|false|false|C1420621;C1515258|TCAP gene;Telephone Number|Tele
Event|Event|SIMPLE_SEGMENT|2714,2717|false|false|false|||NSR
Finding|Molecular Function|SIMPLE_SEGMENT|2714,2717|false|false|false|C1704493;C2700623|Neutral Sidebent Rotated|NSR
Finding|Pathologic Function|SIMPLE_SEGMENT|2714,2717|false|false|false|C1704493;C2700623|Neutral Sidebent Rotated|NSR
Finding|Classification|SIMPLE_SEGMENT|2718,2721|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Finding|Gene or Genome|SIMPLE_SEGMENT|2718,2721|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Finding|Finding|SIMPLE_SEGMENT|2732,2742|false|false|false|C0231835|Tachypnea|tachypneic
Finding|Sign or Symptom|SIMPLE_SEGMENT|2761,2769|false|false|false|C0043144|Wheezing|wheezing
Event|Event|SIMPLE_SEGMENT|2787,2796|false|false|false|||finishing
Event|Event|SIMPLE_SEGMENT|2797,2806|false|false|false|||sentences
Finding|Intellectual Product|SIMPLE_SEGMENT|2797,2806|false|false|false|C0876929|Sentence|sentences
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2808,2813|false|false|false|C1512338|HEENT|HEENT
Event|Event|SIMPLE_SEGMENT|2821,2827|false|false|false|||PERRLA
Finding|Finding|SIMPLE_SEGMENT|2821,2827|false|false|false|C2143306|PERRLA|PERRLA
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2829,2833|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|SIMPLE_SEGMENT|2829,2833|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|SIMPLE_SEGMENT|2829,2833|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|SIMPLE_SEGMENT|2838,2841|false|false|false|||JVD
Finding|Finding|SIMPLE_SEGMENT|2838,2841|true|false|false|C0425687|Jugular venous engorgement|JVD
Event|Event|SIMPLE_SEGMENT|2859,2868|false|false|false|||difficult
Finding|Finding|SIMPLE_SEGMENT|2859,2868|false|false|false|C0332218|Difficult (qualifier value)|difficult
Event|Event|SIMPLE_SEGMENT|2872,2882|false|false|false|||appreciate
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2883,2888|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2883,2888|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|2883,2888|false|false|false|C0795691|HEART PROBLEM|heart
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2883,2895|false|false|false|C4050434||heart sounds
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|2883,2895|false|false|false|C0018820|Heart Sounds|heart sounds
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2883,2895|false|false|false|C2230284|auscultation of heart sounds|heart sounds
Event|Event|SIMPLE_SEGMENT|2889,2895|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2889,2895|false|false|false|C0037709||sounds
Finding|Idea or Concept|SIMPLE_SEGMENT|2904,2915|false|false|false|C0750502|Significant|significant
Event|Event|SIMPLE_SEGMENT|2916,2923|false|false|false|||rhonchi
Finding|Finding|SIMPLE_SEGMENT|2916,2923|false|false|false|C0035508|Rhonchi|rhonchi
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2925,2930|false|false|false|C0024109|Lung|LUNGS
Event|Event|SIMPLE_SEGMENT|2936,2943|false|false|false|||rhonchi
Finding|Finding|SIMPLE_SEGMENT|2936,2943|false|false|false|C0035508|Rhonchi|rhonchi
Finding|Intellectual Product|SIMPLE_SEGMENT|2958,2962|false|false|false|C1547225|Mild Severity of Illness Code|mild
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2963,2966|false|false|false|C0082420|Endoglin, human|end
Drug|Immunologic Factor|SIMPLE_SEGMENT|2963,2966|false|false|false|C0082420|Endoglin, human|end
Finding|Functional Concept|SIMPLE_SEGMENT|2963,2966|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Finding|Gene or Genome|SIMPLE_SEGMENT|2963,2966|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Finding|Organism Function|SIMPLE_SEGMENT|2967,2977|false|false|false|C0231800|Expiration, Respiratory|expiratory
Finding|Sign or Symptom|SIMPLE_SEGMENT|2967,2986|false|false|false|C0231875|Expiratory wheezing|expiratory wheezing
Event|Event|SIMPLE_SEGMENT|2978,2986|false|false|false|||wheezing
Finding|Sign or Symptom|SIMPLE_SEGMENT|2978,2986|false|false|false|C0043144|Wheezing|wheezing
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2994,2998|false|false|false|C2987514|Anatomical base|base
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2994,2998|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|2994,2998|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|2994,2998|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Finding|Gene or Genome|SIMPLE_SEGMENT|2994,2998|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Finding|Idea or Concept|SIMPLE_SEGMENT|2994,2998|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Event|Event|SIMPLE_SEGMENT|2999,3007|false|false|false|||crackles
Finding|Finding|SIMPLE_SEGMENT|2999,3007|false|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3008,3011|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|ABD
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|3008,3011|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|ABD
Event|Event|SIMPLE_SEGMENT|3008,3011|false|false|false|||ABD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3013,3017|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|SIMPLE_SEGMENT|3013,3017|false|false|false|||Soft
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|3045,3048|false|false|false|C0015306|Hereditary Multiple Exostoses|EXT
Event|Event|SIMPLE_SEGMENT|3045,3048|false|false|false|||EXT
Finding|Gene or Genome|SIMPLE_SEGMENT|3045,3048|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|EXT
Finding|Conceptual Entity|SIMPLE_SEGMENT|3055,3061|false|false|false|C0442038;C0920847|Circumpennate;Radial|radial
Drug|Food|SIMPLE_SEGMENT|3062,3068|false|false|false|C5890763||pulses
Event|Event|SIMPLE_SEGMENT|3062,3068|false|false|false|||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|3062,3068|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|3062,3068|false|false|false|C0034107|Pulse taking|pulses
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3070,3075|false|false|false|C4048756|Right arm|R arm
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3072,3075|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|3072,3075|false|false|false|C3495676|Anorectal Malformations|arm
Event|Event|SIMPLE_SEGMENT|3072,3075|false|false|false|||arm
Finding|Gene or Genome|SIMPLE_SEGMENT|3072,3075|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3072,3075|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|SIMPLE_SEGMENT|3072,3075|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3072,3075|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Event|Activity|SIMPLE_SEGMENT|3087,3092|false|false|false|C1882509|put - instruction imperative|place
Event|Event|SIMPLE_SEGMENT|3087,3092|false|false|false|||place
Finding|Functional Concept|SIMPLE_SEGMENT|3087,3092|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|SIMPLE_SEGMENT|3087,3092|false|false|false|C1533810||place
Event|Event|SIMPLE_SEGMENT|3097,3103|false|false|false|||normal
Event|Event|SIMPLE_SEGMENT|3105,3110|false|false|false|||motor
Finding|Functional Concept|SIMPLE_SEGMENT|3105,3110|false|false|false|C1513492|motor movement|motor
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3111,3127|false|false|false|C0036658|Sensory perception|sensory function
Event|Event|SIMPLE_SEGMENT|3119,3127|false|false|false|||function
Finding|Finding|SIMPLE_SEGMENT|3119,3127|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|3119,3127|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|3119,3127|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|SIMPLE_SEGMENT|3119,3127|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Event|Event|SIMPLE_SEGMENT|3128,3134|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|3128,3134|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|SIMPLE_SEGMENT|3170,3181|false|false|false|||dopplerable
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3211,3215|false|false|false|C0009443;C0024117|Chronic Obstructive Airway Disease;Common Cold|cold
Drug|Organic Chemical|SIMPLE_SEGMENT|3211,3215|false|false|false|C0719425|Cold brand of chlorpheniramine-phenylpropanolamine|cold
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3211,3215|false|false|false|C0719425|Cold brand of chlorpheniramine-phenylpropanolamine|cold
Event|Event|SIMPLE_SEGMENT|3211,3215|false|false|false|||cold
Finding|Organism Function|SIMPLE_SEGMENT|3211,3215|false|false|false|C0234192|Cold Sensation|cold
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3211,3215|false|false|false|C0009264|Cold Temperature|cold
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3211,3215|false|false|false|C0010412|Cold Therapy|cold
Event|Event|SIMPLE_SEGMENT|3220,3226|false|false|false|||normal
Event|Event|SIMPLE_SEGMENT|3228,3237|false|false|false|||sensation
Finding|Finding|SIMPLE_SEGMENT|3228,3237|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3228,3237|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|SIMPLE_SEGMENT|3228,3237|false|false|false|C2229507|sensory exam|sensation
Finding|Functional Concept|SIMPLE_SEGMENT|3246,3251|false|false|false|C1513492|motor movement|motor
Event|Event|SIMPLE_SEGMENT|3252,3260|false|false|false|||strength
Finding|Idea or Concept|SIMPLE_SEGMENT|3252,3260|false|false|false|C0808080|Strength (attribute)|strength
Event|Event|SIMPLE_SEGMENT|3265,3268|false|false|false|||ROM
Finding|Finding|SIMPLE_SEGMENT|3265,3268|false|false|false|C0948106;C1419600|ROM1 gene;Rupture of Membranes|ROM
Finding|Gene or Genome|SIMPLE_SEGMENT|3265,3268|false|false|false|C0948106;C1419600|ROM1 gene;Rupture of Membranes|ROM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3265,3268|false|false|false|C1562926|Range of motion technique (procedure)|ROM
Anatomy|Body System|SIMPLE_SEGMENT|3269,3273|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3269,3273|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3269,3273|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|SIMPLE_SEGMENT|3269,3273|false|false|false|||SKIN
Finding|Body Substance|SIMPLE_SEGMENT|3269,3273|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|SIMPLE_SEGMENT|3269,3273|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Event|Event|SIMPLE_SEGMENT|3278,3284|false|false|false|||rashes
Finding|Sign or Symptom|SIMPLE_SEGMENT|3278,3284|true|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Event|Event|SIMPLE_SEGMENT|3288,3295|false|false|false|||chronic
Finding|Intellectual Product|SIMPLE_SEGMENT|3288,3295|true|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|3288,3295|true|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Finding|Pathologic Function|SIMPLE_SEGMENT|3296,3305|false|false|false|C0013604|Edema|edematous
Event|Event|SIMPLE_SEGMENT|3306,3313|false|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|3306,3313|true|false|false|C0392747|Changing|changes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3321,3326|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|3321,3326|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3321,3326|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|3321,3326|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|3321,3326|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|3321,3326|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|3321,3326|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|3331,3340|false|false|false|||attentive
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3355,3370|false|false|false|C0278454|All extremities|all extremities
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3359,3370|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Event|Event|SIMPLE_SEGMENT|3375,3384|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|3375,3384|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|3375,3384|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|3375,3384|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|3375,3384|false|false|false|C0030685|Patient Discharge|discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3401,3407|false|false|false|C0944911||Weight
Event|Event|SIMPLE_SEGMENT|3401,3407|false|false|false|||Weight
Finding|Finding|SIMPLE_SEGMENT|3401,3407|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|Weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|3401,3407|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|Weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|3401,3407|false|false|false|C1305866|Weighing patient|Weight
Event|Event|SIMPLE_SEGMENT|3506,3509|false|false|false|||Gen
Finding|Classification|SIMPLE_SEGMENT|3506,3509|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Finding|Gene or Genome|SIMPLE_SEGMENT|3506,3509|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Event|Event|SIMPLE_SEGMENT|3511,3516|false|false|false|||awake
Finding|Finding|SIMPLE_SEGMENT|3511,3516|false|false|false|C0234422|Awake (finding)|awake
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3518,3523|false|false|false|C5890168||alert
Drug|Organic Chemical|SIMPLE_SEGMENT|3518,3523|false|false|false|C0718338|Alert brand of caffeine|alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3518,3523|false|false|false|C0718338|Alert brand of caffeine|alert
Event|Event|SIMPLE_SEGMENT|3518,3523|false|false|false|||alert
Finding|Finding|SIMPLE_SEGMENT|3518,3523|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Functional Concept|SIMPLE_SEGMENT|3518,3523|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Intellectual Product|SIMPLE_SEGMENT|3518,3523|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Event|Event|SIMPLE_SEGMENT|3525,3533|false|false|false|||oriented
Finding|Finding|SIMPLE_SEGMENT|3525,3533|false|false|false|C1961028|Oriented to place|oriented
Event|Event|SIMPLE_SEGMENT|3537,3541|false|false|false|||self
Finding|Idea or Concept|SIMPLE_SEGMENT|3537,3541|false|false|false|C0036588;C1551994|Self;subscriber - self|self
Finding|Intellectual Product|SIMPLE_SEGMENT|3537,3541|false|false|false|C0036588;C1551994|Self;subscriber - self|self
Event|Event|SIMPLE_SEGMENT|3549,3557|false|false|false|||hospital
Finding|Idea or Concept|SIMPLE_SEGMENT|3549,3557|false|false|false|C1547192|Organization unit type - Hospital|hospital
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3558,3563|false|false|false|C1512338|HEENT|HEENT
Event|Event|SIMPLE_SEGMENT|3571,3577|false|false|false|||PERRLA
Finding|Finding|SIMPLE_SEGMENT|3571,3577|false|false|false|C2143306|PERRLA|PERRLA
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3579,3583|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|SIMPLE_SEGMENT|3579,3583|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|SIMPLE_SEGMENT|3579,3583|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|SIMPLE_SEGMENT|3588,3591|false|false|false|||JVD
Finding|Finding|SIMPLE_SEGMENT|3588,3591|true|false|false|C0425687|Jugular venous engorgement|JVD
Event|Event|SIMPLE_SEGMENT|3609,3618|false|false|false|||difficult
Finding|Finding|SIMPLE_SEGMENT|3609,3618|false|false|false|C0332218|Difficult (qualifier value)|difficult
Event|Event|SIMPLE_SEGMENT|3622,3632|false|false|false|||appreciate
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3633,3638|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3633,3638|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|3633,3638|false|false|false|C0795691|HEART PROBLEM|heart
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3633,3645|false|false|false|C4050434||heart sounds
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3633,3645|false|false|false|C0018820|Heart Sounds|heart sounds
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3633,3645|false|false|false|C2230284|auscultation of heart sounds|heart sounds
Event|Event|SIMPLE_SEGMENT|3639,3645|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3639,3645|false|false|false|C0037709||sounds
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3647,3652|false|false|false|C0024109|Lung|LUNGS
Event|Event|SIMPLE_SEGMENT|3665,3673|false|false|false|||crackles
Finding|Finding|SIMPLE_SEGMENT|3665,3673|false|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3674,3677|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|ABD
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|3674,3677|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|ABD
Event|Event|SIMPLE_SEGMENT|3674,3677|false|false|false|||ABD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3679,3683|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|SIMPLE_SEGMENT|3679,3683|false|false|false|||Soft
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|3711,3714|false|false|false|C0015306|Hereditary Multiple Exostoses|EXT
Event|Event|SIMPLE_SEGMENT|3711,3714|false|false|false|||EXT
Finding|Gene or Genome|SIMPLE_SEGMENT|3711,3714|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|EXT
Finding|Conceptual Entity|SIMPLE_SEGMENT|3723,3729|false|false|false|C0442038;C0920847|Circumpennate;Radial|radial
Drug|Food|SIMPLE_SEGMENT|3730,3736|false|false|false|C5890763||pulses
Event|Event|SIMPLE_SEGMENT|3730,3736|false|false|false|||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|3730,3736|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|3730,3736|false|false|false|C0034107|Pulse taking|pulses
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3738,3743|false|false|false|C4048756|Right arm|R arm
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3740,3743|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|3740,3743|false|false|false|C3495676|Anorectal Malformations|arm
Finding|Gene or Genome|SIMPLE_SEGMENT|3740,3743|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3740,3743|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|SIMPLE_SEGMENT|3740,3743|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3740,3743|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Event|Event|SIMPLE_SEGMENT|3745,3751|false|false|false|||normal
Finding|Functional Concept|SIMPLE_SEGMENT|3752,3757|false|false|false|C1513492|motor movement|motor
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3758,3774|false|true|false|C0036658|Sensory perception|sensory function
Event|Event|SIMPLE_SEGMENT|3766,3774|false|false|false|||function
Finding|Finding|SIMPLE_SEGMENT|3766,3774|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|3766,3774|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|3766,3774|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|SIMPLE_SEGMENT|3766,3774|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Event|Event|SIMPLE_SEGMENT|3776,3782|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|3776,3782|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|SIMPLE_SEGMENT|3830,3835|false|false|false|||trace
Finding|Functional Concept|SIMPLE_SEGMENT|3830,3835|false|false|false|C1883002|Sequence Chromatogram|trace
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3837,3842|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|3837,3842|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|3837,3842|false|false|false|C0013604|Edema|edema
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3865,3869|false|false|false|C0009443;C0024117|Chronic Obstructive Airway Disease;Common Cold|cold
Drug|Organic Chemical|SIMPLE_SEGMENT|3865,3869|false|false|false|C0719425|Cold brand of chlorpheniramine-phenylpropanolamine|cold
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3865,3869|false|false|false|C0719425|Cold brand of chlorpheniramine-phenylpropanolamine|cold
Event|Event|SIMPLE_SEGMENT|3865,3869|false|false|false|||cold
Finding|Organism Function|SIMPLE_SEGMENT|3865,3869|false|false|false|C0234192|Cold Sensation|cold
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3865,3869|false|false|false|C0009264|Cold Temperature|cold
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3865,3869|false|false|false|C0010412|Cold Therapy|cold
Event|Event|SIMPLE_SEGMENT|3881,3890|false|false|false|||sensation
Finding|Finding|SIMPLE_SEGMENT|3881,3890|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3881,3890|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|SIMPLE_SEGMENT|3881,3890|false|false|false|C2229507|sensory exam|sensation
Finding|Functional Concept|SIMPLE_SEGMENT|3900,3905|false|false|false|C1513492|motor movement|motor
Event|Event|SIMPLE_SEGMENT|3906,3914|false|false|false|||strength
Finding|Idea or Concept|SIMPLE_SEGMENT|3906,3914|false|false|false|C0808080|Strength (attribute)|strength
Event|Event|SIMPLE_SEGMENT|3919,3922|false|false|false|||ROM
Finding|Finding|SIMPLE_SEGMENT|3919,3922|false|false|false|C0948106;C1419600|ROM1 gene;Rupture of Membranes|ROM
Finding|Gene or Genome|SIMPLE_SEGMENT|3919,3922|false|false|false|C0948106;C1419600|ROM1 gene;Rupture of Membranes|ROM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3919,3922|false|false|false|C1562926|Range of motion technique (procedure)|ROM
Anatomy|Body System|SIMPLE_SEGMENT|3923,3927|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3923,3927|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3923,3927|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|SIMPLE_SEGMENT|3923,3927|false|false|false|||SKIN
Finding|Body Substance|SIMPLE_SEGMENT|3923,3927|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|SIMPLE_SEGMENT|3923,3927|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Event|Event|SIMPLE_SEGMENT|3932,3938|false|false|false|||rashes
Finding|Sign or Symptom|SIMPLE_SEGMENT|3932,3938|true|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Event|Event|SIMPLE_SEGMENT|3942,3949|false|false|false|||chronic
Finding|Intellectual Product|SIMPLE_SEGMENT|3942,3949|true|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|3942,3949|true|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Finding|Pathologic Function|SIMPLE_SEGMENT|3950,3959|false|false|false|C0013604|Edema|edematous
Event|Event|SIMPLE_SEGMENT|3960,3967|false|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|3960,3967|true|false|false|C0392747|Changing|changes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3975,3980|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|3975,3980|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3975,3980|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|3975,3980|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|3975,3980|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|3975,3980|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|3975,3980|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|3985,3994|false|false|false|||attentive
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4009,4024|false|false|false|C0278454|All extremities|all extremities
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4013,4024|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Event|Event|SIMPLE_SEGMENT|4047,4051|false|false|false|||Labs
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4047,4051|false|false|false|C0587081|Laboratory test finding|Labs
Event|Event|SIMPLE_SEGMENT|4055,4064|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|4055,4064|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Anatomy|Cell|SIMPLE_SEGMENT|4100,4103|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|4110,4113|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4110,4113|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4110,4113|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4120,4123|false|false|false|C0019046|Hemoglobin|HGB
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4120,4123|false|false|false|C0019046|Hemoglobin|HGB
Event|Event|SIMPLE_SEGMENT|4120,4123|false|false|false|||HGB
Finding|Gene or Genome|SIMPLE_SEGMENT|4120,4123|false|false|false|C1424337|CYGB gene|HGB
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4120,4123|false|false|false|C0019029|Hemoglobin concentration|HGB
Event|Event|SIMPLE_SEGMENT|4129,4132|false|false|false|||HCT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4129,4132|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4129,4132|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Disorder|Virus|SIMPLE_SEGMENT|4138,4141|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|4138,4141|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4138,4141|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4138,4141|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4138,4141|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|4146,4149|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4146,4149|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|4146,4149|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|4146,4149|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|4146,4149|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4146,4149|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|4155,4159|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4155,4159|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Event|Event|SIMPLE_SEGMENT|4199,4202|false|false|false|||PLT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4199,4202|false|false|false|C0201617|Primed lymphocyte test|PLT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4203,4206|false|false|false|C5441956|Megakaryocyte-Potentiating Factor, human|SMR
Drug|Immunologic Factor|SIMPLE_SEGMENT|4203,4206|false|false|false|C5441956|Megakaryocyte-Potentiating Factor, human|SMR
Event|Event|SIMPLE_SEGMENT|4203,4206|false|false|false|||SMR
Finding|Gene or Genome|SIMPLE_SEGMENT|4203,4206|false|false|false|C1334533;C1704868|MSLN gene;MSLN wt Allele|SMR
Event|Event|SIMPLE_SEGMENT|4214,4217|false|false|false|||PLT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4214,4217|false|false|false|C0201617|Primed lymphocyte test|PLT
Finding|Body Substance|SIMPLE_SEGMENT|4262,4268|false|false|false|C0024202|Lymph|LYMPHS
Drug|Antibiotic|SIMPLE_SEGMENT|4272,4277|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4272,4277|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Organic Chemical|SIMPLE_SEGMENT|4272,4277|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4280,4283|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|EOS
Event|Event|SIMPLE_SEGMENT|4280,4283|false|false|false|||EOS
Finding|Gene or Genome|SIMPLE_SEGMENT|4280,4283|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|EOS
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4397,4400|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|SIMPLE_SEGMENT|4397,4400|false|false|false|||PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4397,4400|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4425,4432|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|SIMPLE_SEGMENT|4425,4432|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4425,4432|false|false|false|C0017725|glucose|GLUCOSE
Event|Event|SIMPLE_SEGMENT|4425,4432|false|false|false|||GLUCOSE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4425,4432|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4425,4432|false|false|false|C0337438|Glucose measurement|GLUCOSE
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4438,4442|false|false|false|C0041942|urea|UREA
Drug|Organic Chemical|SIMPLE_SEGMENT|4438,4442|false|false|false|C0041942|urea|UREA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4438,4442|false|false|false|C0041942|urea|UREA
Event|Event|SIMPLE_SEGMENT|4438,4442|false|false|false|||UREA
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4438,4442|false|false|false|C0523961|Urea measurement|UREA
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4461,4467|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4461,4467|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4461,4467|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Event|Event|SIMPLE_SEGMENT|4461,4467|false|false|false|||SODIUM
Finding|Physiologic Function|SIMPLE_SEGMENT|4461,4467|false|false|false|C4553025|Sodium metabolic function|SODIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4461,4467|false|false|false|C0337443|Sodium measurement|SODIUM
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4473,4482|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4473,4482|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Food|SIMPLE_SEGMENT|4473,4482|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4473,4482|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4473,4482|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Finding|Physiologic Function|SIMPLE_SEGMENT|4473,4482|false|false|false|C4553027|Potassium metabolic function|POTASSIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4473,4482|false|false|false|C0202194|Potassium measurement|POTASSIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4487,4495|false|false|false|C0008203;C0596019|Chlorides;chloride ion|CHLORIDE
Event|Event|SIMPLE_SEGMENT|4487,4495|false|false|false|||CHLORIDE
Finding|Physiologic Function|SIMPLE_SEGMENT|4487,4495|false|false|false|C4553021|Chloride metabolic function|CHLORIDE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4487,4495|false|false|false|C0201952|Chloride measurement|CHLORIDE
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4505,4508|false|false|false|C0007012|carbon dioxide|CO2
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4505,4508|false|false|false|C0007012|carbon dioxide|CO2
Finding|Finding|SIMPLE_SEGMENT|4505,4508|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Finding|Gene or Genome|SIMPLE_SEGMENT|4505,4508|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4513,4518|false|false|false|C0003075|Anions|ANION
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4520,4523|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4520,4523|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Event|Event|SIMPLE_SEGMENT|4520,4523|false|false|false|||GAP
Finding|Gene or Genome|SIMPLE_SEGMENT|4520,4523|false|false|false|C1419277;C2984552|RASA1 gene;RASA1 wt Allele|GAP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4542,4549|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4542,4549|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4542,4549|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4542,4549|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Vitamin|SIMPLE_SEGMENT|4542,4549|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Event|Event|SIMPLE_SEGMENT|4542,4549|false|false|false|||CALCIUM
Finding|Physiologic Function|SIMPLE_SEGMENT|4542,4549|false|false|false|C4553026|Calcium metabolic function|CALCIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4542,4549|false|false|false|C0201925|Calcium measurement|CALCIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4555,4564|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4555,4564|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4555,4564|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4555,4564|false|false|false|C0523826|Phosphate measurement|PHOSPHATE
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4569,4578|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4569,4578|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4569,4578|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4569,4578|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4569,4578|false|false|false|C0373675|Magnesium measurement|MAGNESIUM
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4611,4616|false|false|false|C0019018|Glycosylated hemoglobin A|HbA1c
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4611,4616|false|false|false|C0019018|Glycosylated hemoglobin A|HbA1c
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4611,4616|false|false|false|C0202054|Glucohemoglobin measurement|HbA1c
Finding|Gene or Genome|SIMPLE_SEGMENT|4621,4624|false|false|false|C1416571|KCNH1 gene|eAG
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4643,4648|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|SIMPLE_SEGMENT|4643,4648|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|SIMPLE_SEGMENT|4643,4648|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4643,4648|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4694,4697|false|false|false|C0023821|High Density Lipoproteins|HDL
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4694,4697|false|false|false|C0023821|High Density Lipoproteins|HDL
Event|Event|SIMPLE_SEGMENT|4694,4697|false|false|false|||HDL
Finding|Gene or Genome|SIMPLE_SEGMENT|4694,4697|false|false|false|C3715113|HSD11B1 wt Allele|HDL
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4694,4697|false|false|false|C0392885|High density lipoprotein measurement|HDL
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4711,4714|false|false|false|C0023821|High Density Lipoproteins|HDL
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4711,4714|false|false|false|C0023821|High Density Lipoproteins|HDL
Event|Event|SIMPLE_SEGMENT|4711,4714|false|false|false|||HDL
Finding|Gene or Genome|SIMPLE_SEGMENT|4711,4714|false|false|false|C3715113|HSD11B1 wt Allele|HDL
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4711,4714|false|false|false|C0392885|High density lipoprotein measurement|HDL
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4720,4723|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Drug|Organic Chemical|SIMPLE_SEGMENT|4720,4723|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Event|Event|SIMPLE_SEGMENT|4720,4723|false|false|false|||LDL
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4720,4723|false|false|false|C0202117|Low density lipoprotein cholesterol measurement|LDL
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4724,4728|false|false|false|C4084820|Intracalcarine cortex|CALC
Finding|Gene or Genome|SIMPLE_SEGMENT|4724,4728|false|false|false|C1413147|MICU1 gene|CALC
Event|Event|SIMPLE_SEGMENT|4852,4856|false|false|false|||Labs
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4852,4856|false|false|false|C0587081|Laboratory test finding|Labs
Event|Event|SIMPLE_SEGMENT|4860,4869|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|4860,4869|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|4860,4869|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|4860,4869|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|4860,4869|false|false|false|C0030685|Patient Discharge|Discharge
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4903,4908|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4903,4908|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4903,4908|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|4909,4912|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|4919,4922|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4919,4922|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4919,4922|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4929,4932|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4929,4932|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|4929,4932|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4929,4932|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4939,4942|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4939,4942|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|4950,4953|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|4950,4953|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4950,4953|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4950,4953|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4950,4953|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|4957,4960|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4957,4960|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|4957,4960|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|4957,4960|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|4957,4960|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4957,4960|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|4966,4970|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4966,4970|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4997,5000|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5017,5022|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5017,5022|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5017,5022|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5041,5047|false|false|false|C0024202|Lymph|Lymphs
Drug|Antibiotic|SIMPLE_SEGMENT|5052,5057|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5052,5057|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|SIMPLE_SEGMENT|5052,5057|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5061,5064|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Event|Event|SIMPLE_SEGMENT|5061,5064|false|false|false|||Eos
Finding|Gene or Genome|SIMPLE_SEGMENT|5061,5064|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5175,5180|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5175,5180|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5175,5180|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5185,5188|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|SIMPLE_SEGMENT|5185,5188|false|false|false|||PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5185,5188|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5210,5215|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5210,5215|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5210,5215|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|5210,5223|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5210,5223|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5210,5223|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5216,5223|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|5216,5223|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5216,5223|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|5216,5223|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5216,5223|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5216,5223|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5270,5274|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5270,5274|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5270,5274|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5299,5304|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5299,5304|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5299,5304|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5305,5308|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5305,5308|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|5305,5308|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|5305,5308|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|5305,5308|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|5305,5308|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|5305,5308|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5305,5308|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5312,5315|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5312,5315|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5312,5315|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5312,5315|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|5312,5315|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|5312,5315|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|5312,5315|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5322,5325|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Drug|Enzyme|SIMPLE_SEGMENT|5322,5325|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Event|Event|SIMPLE_SEGMENT|5322,5325|false|false|false|||LDH
Finding|Finding|SIMPLE_SEGMENT|5322,5325|false|false|false|C0851148|Lifetime Drinking History|LDH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5322,5325|false|false|false|C0202113|Lactate dehydrogenase measurement|LDH
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5332,5339|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|SIMPLE_SEGMENT|5332,5339|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5368,5373|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5368,5373|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5368,5373|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5368,5381|false|false|false|C0853248|Blood albumin|BLOOD Albumin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5374,5381|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5374,5381|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5374,5381|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Event|Event|SIMPLE_SEGMENT|5374,5381|false|false|false|||Albumin
Finding|Gene or Genome|SIMPLE_SEGMENT|5374,5381|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Finding|Physiologic Function|SIMPLE_SEGMENT|5374,5381|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5374,5381|false|false|false|C0201838|Albumin measurement|Albumin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5387,5394|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|5387,5394|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5387,5394|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5387,5394|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|5387,5394|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|5387,5394|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|5387,5394|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5387,5394|false|false|false|C0201925|Calcium measurement|Calcium
Event|Event|SIMPLE_SEGMENT|5425,5432|false|false|false|||Imaging
Finding|Finding|SIMPLE_SEGMENT|5425,5432|false|false|false|C0740845|Imaging problem|Imaging
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5425,5432|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|Imaging
Event|Event|SIMPLE_SEGMENT|5452,5455|false|false|false|||TTE
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5452,5455|false|false|false|C0430462|Transthoracic echocardiography|TTE
Finding|Functional Concept|SIMPLE_SEGMENT|5465,5469|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5465,5476|false|false|false|C0225860|Left atrial structure|left atrium
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5470,5476|false|false|false|C0018792|Heart Atrium|atrium
Event|Event|SIMPLE_SEGMENT|5487,5494|false|false|false|||dilated
Finding|Functional Concept|SIMPLE_SEGMENT|5510,5515|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5516,5522|false|false|false|C0018792|Heart Atrium|atrial
Event|Event|SIMPLE_SEGMENT|5524,5532|false|false|false|||pressure
Finding|Finding|SIMPLE_SEGMENT|5524,5532|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|5524,5532|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5524,5532|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|5524,5532|false|false|false|C0033095||pressure
Finding|Functional Concept|SIMPLE_SEGMENT|5546,5550|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5546,5567|false|false|false|C0504053|Wall of left ventricle|Left ventricular wall
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5551,5562|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5551,5567|false|false|false|C0507618|Wall of ventricle|ventricular wall
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5585,5591|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|5585,5591|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5585,5591|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Event|Event|SIMPLE_SEGMENT|5592,5596|false|false|false|||size
Event|Event|SIMPLE_SEGMENT|5601,5607|false|false|false|||normal
Finding|Intellectual Product|SIMPLE_SEGMENT|5609,5616|false|false|false|C0282416|Overall Publication Type|Overall
Finding|Functional Concept|SIMPLE_SEGMENT|5617,5621|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5622,5633|false|false|false|C0018827|Heart Ventricle|ventricular
Event|Event|SIMPLE_SEGMENT|5634,5642|false|false|false|||systolic
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5634,5642|false|false|false|C0039155|Systole|systolic
Event|Event|SIMPLE_SEGMENT|5644,5652|false|false|false|||function
Finding|Finding|SIMPLE_SEGMENT|5644,5652|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|5644,5652|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|5644,5652|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|SIMPLE_SEGMENT|5644,5652|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Finding|SIMPLE_SEGMENT|5656,5666|false|false|false|C4085643;C5201148;C5962468|Moderate;Moderate Effect;Moderate Response|moderately
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|5667,5676|false|false|false|C0344315|Depressed mood|depressed
Event|Event|SIMPLE_SEGMENT|5667,5676|false|false|false|||depressed
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5678,5682|false|false|false|C0428772|Left ventricular ejection fraction|LVEF
Event|Event|SIMPLE_SEGMENT|5678,5682|false|false|false|||LVEF
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5678,5682|false|false|false|C3837267|LVEF (procedure)|LVEF
Event|Activity|SIMPLE_SEGMENT|5695,5705|false|false|false|C1516048|Assessed|assessment
Event|Event|SIMPLE_SEGMENT|5695,5705|false|false|false|||assessment
Finding|Intellectual Product|SIMPLE_SEGMENT|5695,5705|false|false|false|C0679207|Knowledge acquisition using a method of assessment|assessment
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5695,5705|false|false|false|C0028708;C0031809;C0220825;C0542573;C0549068;C0549070;C0549071;C0549072;C0549073;C0549074;C0549075;C0549076;C0549078;C0549079;C0549080;C1161151;C1261322;C2237115|Evaluation;Evaluation procedure;Nutrition Assessment;Personal care assessment;Physical Examination;assessment of cognitive functions|assessment
Procedure|Health Care Activity|SIMPLE_SEGMENT|5695,5705|false|false|false|C0028708;C0031809;C0220825;C0542573;C0549068;C0549070;C0549071;C0549072;C0549073;C0549074;C0549075;C0549076;C0549078;C0549079;C0549080;C1161151;C1261322;C2237115|Evaluation;Evaluation procedure;Nutrition Assessment;Personal care assessment;Physical Examination;assessment of cognitive functions|assessment
Event|Event|SIMPLE_SEGMENT|5707,5714|false|false|false|||limited
Finding|Finding|SIMPLE_SEGMENT|5718,5734|false|false|false|C2828075|Suboptimal Image Reason|suboptimal image
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5729,5734|false|false|false|C1846009|Intrauterine growth restriction, metaphyseal dysplasia, adrenal hypoplasia congenita, and genital anomaly syndrome|image
Event|Event|SIMPLE_SEGMENT|5729,5734|false|false|false|||image
Finding|Intellectual Product|SIMPLE_SEGMENT|5729,5734|false|false|false|C1696103;C1704254;C1704922;C3542466|Image;Image (foundation metadata concept);Medical Image;image - dosage form|image
Finding|Idea or Concept|SIMPLE_SEGMENT|5747,5758|false|false|false|C0750502|Significant|significant
Event|Event|SIMPLE_SEGMENT|5759,5763|false|false|false|||beat
Event|Event|SIMPLE_SEGMENT|5767,5771|false|false|false|||beat
Event|Event|SIMPLE_SEGMENT|5773,5784|false|false|false|||variability
Finding|Conceptual Entity|SIMPLE_SEGMENT|5773,5784|false|false|false|C2827666|Variability|variability
Event|Event|SIMPLE_SEGMENT|5796,5807|false|false|false|||hypokinesis
Finding|Finding|SIMPLE_SEGMENT|5796,5807|false|false|false|C0086439|Hypokinesia|hypokinesis
Event|Event|SIMPLE_SEGMENT|5829,5837|false|false|false|||segments
Anatomy|Cell Component|SIMPLE_SEGMENT|5843,5847|false|false|false|C3890171|dinoflagellate apex|apex
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5843,5847|false|false|false|C0140145|APEX1 protein, human|apex
Drug|Enzyme|SIMPLE_SEGMENT|5843,5847|false|false|false|C0140145|APEX1 protein, human|apex
Finding|Gene or Genome|SIMPLE_SEGMENT|5843,5847|false|false|false|C1332102|APEX1 gene|apex
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5861,5872|false|false|false|C0018827|Heart Ventricle|ventricular
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|5861,5886|true|false|false|C0018818|Ventricular Septal Defects|ventricular septal defect
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|5873,5886|true|false|false|C0018816;C5779791|Congenital septal defect of heart;Heart Septal Defects|septal defect
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|5873,5886|true|false|false|C0018816;C5779791|Congenital septal defect of heart;Heart Septal Defects|septal defect
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5880,5886|true|false|false|C1861101|THYROID HORMONE PLASMA MEMBRANE TRANSPORT DEFECT|defect
Event|Event|SIMPLE_SEGMENT|5880,5886|false|false|false|||defect
Finding|Functional Concept|SIMPLE_SEGMENT|5880,5886|true|false|false|C1457869|Defect|defect
Finding|Functional Concept|SIMPLE_SEGMENT|5888,5893|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5895,5906|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5907,5914|false|false|false|C0935616|chamber [body part]|chamber
Event|Event|SIMPLE_SEGMENT|5915,5919|false|false|false|||size
Event|Event|SIMPLE_SEGMENT|5924,5928|false|false|false|||free
Finding|Functional Concept|SIMPLE_SEGMENT|5924,5928|false|false|false|C0332296|Free of (attribute)|free
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5929,5940|false|false|false|C1980023|Wall motion|wall motion
Event|Event|SIMPLE_SEGMENT|5934,5940|false|false|false|||motion
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|5934,5940|false|false|false|C0026597|Motion|motion
Event|Event|SIMPLE_SEGMENT|5945,5951|false|false|false|||normal
Finding|Functional Concept|SIMPLE_SEGMENT|5958,5967|false|false|false|C1547175;C1962987|Ascend (action);Sequencing - Ascending|ascending
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5958,5973|false|false|false|C0003956|Ascending aorta structure|ascending aorta
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5968,5973|false|false|false|C0003483;C4037978|Aorta;Chest+Abdomen>Aorta|aorta
Procedure|Health Care Activity|SIMPLE_SEGMENT|5968,5973|false|false|false|C0869784|Procedure on aorta|aorta
Event|Event|SIMPLE_SEGMENT|5984,5991|false|false|false|||dilated
Event|Event|SIMPLE_SEGMENT|5997,6003|false|false|false|||number
Finding|Idea or Concept|SIMPLE_SEGMENT|5997,6003|false|false|false|C1554106|MDF AttributeType - Number|number
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6007,6013|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6007,6019|false|false|false|C0003501;C4533215|Aortic valve structure;Chest>Aortic valve|aortic valve
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6014,6019|false|false|false|C1186983|Anatomical valve|valve
Event|Event|SIMPLE_SEGMENT|6021,6029|false|false|false|||leaflets
Event|Event|SIMPLE_SEGMENT|6040,6050|false|false|false|||determined
Finding|Intellectual Product|SIMPLE_SEGMENT|6061,6065|false|false|false|C1547225|Mild Severity of Illness Code|mild
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6066,6072|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6066,6078|false|false|false|C0003501;C4533215|Aortic valve structure;Chest>Aortic valve|aortic valve
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6073,6078|false|false|false|C1186983|Anatomical valve|valve
Event|Event|SIMPLE_SEGMENT|6080,6088|false|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|6080,6088|false|false|false|C1261287|Stenosis|stenosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6090,6095|false|false|false|C1186983|Anatomical valve|valve
Finding|Finding|SIMPLE_SEGMENT|6090,6100|false|false|false|C4687749|Valve Area|valve area
Event|Governmental or Regulatory Activity|SIMPLE_SEGMENT|6096,6100|false|false|false|C1510751|Academic Research Enhancement Awards|area
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|6108,6111|false|false|false|C0555206|Chiari malformation type II|cm2
Event|Event|SIMPLE_SEGMENT|6108,6111|false|false|false|||cm2
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6117,6123|false|false|false|C0003483|Aorta|aortic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6117,6137|true|false|false|C0003504|Aortic Valve Insufficiency|aortic regurgitation
Event|Event|SIMPLE_SEGMENT|6124,6137|false|false|false|||regurgitation
Finding|Finding|SIMPLE_SEGMENT|6124,6137|true|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|SIMPLE_SEGMENT|6124,6137|true|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|6124,6137|true|false|false|C0460152|Regurgitation - mechanism|regurgitation
Event|Event|SIMPLE_SEGMENT|6142,6146|false|false|false|||seen
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6152,6164|false|false|false|C0026264|Mitral Valve|mitral valve
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6159,6164|false|false|false|C1186983|Anatomical valve|valve
Event|Event|SIMPLE_SEGMENT|6165,6172|false|false|false|||appears
Event|Event|SIMPLE_SEGMENT|6186,6192|false|false|false|||normal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6207,6227|false|false|false|C0026266|Mitral Valve Insufficiency|mitral regurgitation
Event|Event|SIMPLE_SEGMENT|6214,6227|false|false|false|||regurgitation
Finding|Finding|SIMPLE_SEGMENT|6214,6227|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|SIMPLE_SEGMENT|6214,6227|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|6214,6227|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6233,6242|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6233,6242|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|6233,6242|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6233,6249|false|false|false|C0034052|Pulmonary artery structure|pulmonary artery
Finding|Finding|SIMPLE_SEGMENT|6233,6267|false|false|false|C0428643|Pulmonary artery systolic pressure|pulmonary artery systolic pressure
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6243,6249|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|6243,6249|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|6250,6258|false|false|false|C0039155|Systole|systolic
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6250,6267|false|false|false|C0871470|Systolic Pressure|systolic pressure
Event|Event|SIMPLE_SEGMENT|6259,6267|false|false|false|||pressure
Finding|Finding|SIMPLE_SEGMENT|6259,6267|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|6259,6267|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|6259,6267|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|6259,6267|false|false|false|C0033095||pressure
Event|Event|SIMPLE_SEGMENT|6282,6292|false|false|false|||determined
Finding|Functional Concept|SIMPLE_SEGMENT|6313,6324|false|false|false|C0205463|Physiological|physiologic
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6326,6337|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6326,6337|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6326,6346|false|false|false|C0031039|Pericardial effusion|pericardial effusion
Finding|Body Substance|SIMPLE_SEGMENT|6326,6346|false|false|false|C1253937|Pericardial effusion body substance|pericardial effusion
Event|Event|SIMPLE_SEGMENT|6338,6346|false|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|6338,6346|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|6338,6346|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|6338,6346|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Event|Event|SIMPLE_SEGMENT|6382,6387|false|false|false|||study
Finding|Intellectual Product|SIMPLE_SEGMENT|6382,6387|false|false|false|C1705923|Study Object|study
Procedure|Research Activity|SIMPLE_SEGMENT|6382,6387|false|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|study
Event|Event|SIMPLE_SEGMENT|6396,6404|false|false|false|||reviewed
Finding|Functional Concept|SIMPLE_SEGMENT|6415,6419|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6420,6431|false|false|false|C0018827|Heart Ventricle|ventricular
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|6432,6440|false|false|false|C0039155|Systole|systolic
Event|Event|SIMPLE_SEGMENT|6441,6449|false|false|false|||function
Finding|Finding|SIMPLE_SEGMENT|6441,6449|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|6441,6449|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|6441,6449|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|SIMPLE_SEGMENT|6441,6449|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Finding|SIMPLE_SEGMENT|6453,6461|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|probably
Finding|Idea or Concept|SIMPLE_SEGMENT|6453,6461|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|probably
Finding|Finding|SIMPLE_SEGMENT|6481,6497|false|false|false|C2828075|Suboptimal Image Reason|suboptimal image
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6492,6497|false|false|false|C1846009|Intrauterine growth restriction, metaphyseal dysplasia, adrenal hypoplasia congenita, and genital anomaly syndrome|image
Event|Event|SIMPLE_SEGMENT|6492,6497|false|false|false|||image
Finding|Intellectual Product|SIMPLE_SEGMENT|6492,6497|false|false|false|C1696103;C1704254;C1704922;C3542466|Image;Image (foundation metadata concept);Medical Image;image - dosage form|image
Event|Event|SIMPLE_SEGMENT|6498,6505|false|false|false|||quality
Event|Event|SIMPLE_SEGMENT|6514,6521|false|false|false|||studies
Procedure|Research Activity|SIMPLE_SEGMENT|6514,6521|false|false|false|C0947630|Scientific Study|studies
Event|Event|SIMPLE_SEGMENT|6523,6532|false|false|false|||precludes
Event|Activity|SIMPLE_SEGMENT|6542,6552|false|false|false|C1707455|Comparison|comparison
Event|Event|SIMPLE_SEGMENT|6542,6552|false|false|false|||comparison
Event|Event|SIMPLE_SEGMENT|6561,6564|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6561,6564|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|SIMPLE_SEGMENT|6567,6577|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|6567,6577|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|6567,6577|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Event|Event|SIMPLE_SEGMENT|6596,6607|false|false|false|||improvement
Finding|Conceptual Entity|SIMPLE_SEGMENT|6596,6607|false|false|false|C2986411|Improvement|improvement
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6611,6621|false|false|false|C0225754|Bilateral lungs|both lungs
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6616,6621|false|false|false|C0024109|Lung|lungs
Finding|Finding|SIMPLE_SEGMENT|6625,6633|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|probably
Finding|Idea or Concept|SIMPLE_SEGMENT|6625,6633|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|probably
Event|Event|SIMPLE_SEGMENT|6642,6650|false|false|false|||decrease
Finding|Finding|SIMPLE_SEGMENT|6642,6650|false|false|false|C0392756|Reduced|decrease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6654,6663|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6654,6663|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|6654,6663|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6665,6670|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|6665,6670|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|6665,6670|false|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|6676,6680|false|false|false|||mild
Finding|Intellectual Product|SIMPLE_SEGMENT|6676,6680|false|false|false|C1547225|Mild Severity of Illness Code|mild
Event|Event|SIMPLE_SEGMENT|6686,6694|false|false|false|||decrease
Finding|Finding|SIMPLE_SEGMENT|6686,6694|false|false|false|C0392756|Reduced|decrease
Finding|Finding|SIMPLE_SEGMENT|6707,6715|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|6707,6715|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Functional Concept|SIMPLE_SEGMENT|6716,6721|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Tissue|SIMPLE_SEGMENT|6722,6729|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6722,6729|false|false|false|C0032226|Pleural Diseases|pleural
Event|Event|SIMPLE_SEGMENT|6731,6739|false|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|6731,6739|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|6731,6739|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|6731,6739|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6752,6757|false|false|false|C1410088|Still|still
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6770,6783|false|false|false|C0521530|Lung consolidation|consolidation
Event|Event|SIMPLE_SEGMENT|6770,6783|false|false|false|||consolidation
Finding|Functional Concept|SIMPLE_SEGMENT|6791,6796|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6791,6807|false|false|false|C1261074|Structure of right upper lobe of lung|right upper lobe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6797,6807|false|false|false|C0225756|Structure of upper lobe of lung|upper lobe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6803,6807|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|SIMPLE_SEGMENT|6803,6807|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Finding|Finding|SIMPLE_SEGMENT|6809,6817|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|probably
Finding|Idea or Concept|SIMPLE_SEGMENT|6809,6817|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|probably
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6819,6828|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|SIMPLE_SEGMENT|6819,6828|false|false|false|||pneumonia
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6847,6852|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|6847,6852|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6847,6857|false|false|false|C0225758|Structure of lower lobe of lung|lower lobe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6853,6857|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|SIMPLE_SEGMENT|6853,6857|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Event|Event|SIMPLE_SEGMENT|6874,6882|false|false|false|||improved
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6886,6891|false|false|false|C0018787;C4037974|Chest>Heart;Heart|Heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6886,6891|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|Heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|6886,6891|false|false|false|C0795691|HEART PROBLEM|Heart
Finding|Finding|SIMPLE_SEGMENT|6886,6896|false|false|false|C0744689|heart size|Heart size
Event|Event|SIMPLE_SEGMENT|6892,6896|false|false|false|||size
Event|Event|SIMPLE_SEGMENT|6902,6908|false|false|false|||normal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6914,6926|true|false|false|C0032326|Pneumothorax|pneumothorax
Event|Event|SIMPLE_SEGMENT|6914,6926|false|false|false|||pneumothorax
Event|Event|SIMPLE_SEGMENT|6930,6935|false|false|false|||MICRO
Finding|Conceptual Entity|SIMPLE_SEGMENT|6930,6935|false|false|false|C3811161;C4049106|Micro (prefix);Microbiology - Laboratory Class|MICRO
Finding|Intellectual Product|SIMPLE_SEGMENT|6930,6935|false|false|false|C3811161;C4049106|Micro (prefix);Microbiology - Laboratory Class|MICRO
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6930,6935|false|false|false|C0085672|Microbiology procedure|MICRO
Finding|Idea or Concept|SIMPLE_SEGMENT|6945,6950|false|false|false|C1546485|Diagnosis Type - Final|FINAL
Finding|Intellectual Product|SIMPLE_SEGMENT|6945,6957|false|false|false|C0460114|Final report|FINAL REPORT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6951,6957|false|false|false|C4255046||REPORT
Event|Event|SIMPLE_SEGMENT|6951,6957|false|false|false|||REPORT
Finding|Intellectual Product|SIMPLE_SEGMENT|6951,6957|false|false|false|C0684224|Report (document)|REPORT
Procedure|Health Care Activity|SIMPLE_SEGMENT|6951,6957|false|false|false|C0700287|Reporting|REPORT
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6979,6982|false|false|false|C0012854|DNA|DNA
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|6979,6982|false|false|false|C0012854|DNA|DNA
Finding|Genetic Function|SIMPLE_SEGMENT|6979,6996|false|false|false|C0683230|dna amplification|DNA amplification
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|6983,6996|false|false|false|C1705759|Gene Amplification Abnormality|amplification
Event|Event|SIMPLE_SEGMENT|6983,6996|false|false|false|||amplification
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|6983,6996|false|false|false|C1521871|Amplification|amplification
Procedure|Molecular Biology Research Technique|SIMPLE_SEGMENT|6983,6996|false|false|false|C1517480|Gene Amplification Technique|amplification
Event|Event|SIMPLE_SEGMENT|6997,7002|false|false|false|||assay
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6997,7002|false|false|false|C0005507;C1510438|Assay;Biological Assay|assay
Finding|Idea or Concept|SIMPLE_SEGMENT|7004,7009|false|false|false|C1546485|Diagnosis Type - Final|Final
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|7055,7063|false|false|false|C4727483|BRAF Gene Rearrangement|Positive
Event|Event|SIMPLE_SEGMENT|7055,7063|false|false|false|||Positive
Finding|Classification|SIMPLE_SEGMENT|7055,7063|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|Positive
Finding|Finding|SIMPLE_SEGMENT|7055,7063|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|Positive
Finding|Finding|SIMPLE_SEGMENT|7055,7067|false|false|false|C1446409|Positive|Positive for
Finding|Intellectual Product|SIMPLE_SEGMENT|7068,7077|false|false|false|C0445332|Toxigenic|toxigenic
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7110,7113|false|false|false|C0012854|DNA|DNA
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|7110,7113|false|false|false|C0012854|DNA|DNA
Event|Event|SIMPLE_SEGMENT|7110,7113|false|false|false|||DNA
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|7123,7136|false|false|false|C1705759|Gene Amplification Abnormality|amplification
Event|Event|SIMPLE_SEGMENT|7123,7136|false|false|false|||amplification
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|7123,7136|false|false|false|C1521871|Amplification|amplification
Procedure|Molecular Biology Research Technique|SIMPLE_SEGMENT|7123,7136|false|false|false|C1517480|Gene Amplification Technique|amplification
Finding|Conceptual Entity|SIMPLE_SEGMENT|7150,7159|false|false|false|C1514811;C1561577;C1706462;C3244318;C4266518|Bibliographic Reference;Reference - HL7UpdateMode;Reference - MdfHmdMetSourceType;Reference Object;Reference source|Reference
Finding|Idea or Concept|SIMPLE_SEGMENT|7150,7159|false|false|false|C1514811;C1561577;C1706462;C3244318;C4266518|Bibliographic Reference;Reference - HL7UpdateMode;Reference - MdfHmdMetSourceType;Reference Object;Reference source|Reference
Finding|Intellectual Product|SIMPLE_SEGMENT|7150,7159|false|false|false|C1514811;C1561577;C1706462;C3244318;C4266518|Bibliographic Reference;Reference - HL7UpdateMode;Reference - MdfHmdMetSourceType;Reference Object;Reference source|Reference
Finding|Intellectual Product|SIMPLE_SEGMENT|7160,7165|false|false|false|C3542016|Concept model range (foundation metadata concept)|Range
Event|Event|SIMPLE_SEGMENT|7166,7174|false|false|false|||Negative
Finding|Classification|SIMPLE_SEGMENT|7166,7174|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Finding|Finding|SIMPLE_SEGMENT|7166,7174|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7166,7174|false|false|false|C5237010|Expression Negative|Negative
Finding|Body Substance|SIMPLE_SEGMENT|7192,7198|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|SPUTUM
Finding|Intellectual Product|SIMPLE_SEGMENT|7192,7198|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|SPUTUM
Event|Event|SIMPLE_SEGMENT|7204,7210|false|false|false|||Source
Finding|Finding|SIMPLE_SEGMENT|7204,7210|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|Source
Finding|Functional Concept|SIMPLE_SEGMENT|7204,7210|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|Source
Finding|Intellectual Product|SIMPLE_SEGMENT|7204,7210|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|Source
Event|Event|SIMPLE_SEGMENT|7212,7224|false|false|false|||Expectorated
Finding|Finding|SIMPLE_SEGMENT|7212,7224|false|false|false|C0566528|Does expectorate|Expectorated
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|7231,7241|false|false|false|C0061856|Gram's stain|GRAM STAIN
Drug|Organic Chemical|SIMPLE_SEGMENT|7231,7241|false|false|false|C0061856|Gram's stain|GRAM STAIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7231,7241|false|false|false|C0200966|Bacterial stain, routine|GRAM STAIN
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|7236,7241|false|false|false|C0038128|Stains|STAIN
Event|Event|SIMPLE_SEGMENT|7236,7241|false|false|false|||STAIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7236,7241|false|false|false|C0487602|Staining method|STAIN
Finding|Idea or Concept|SIMPLE_SEGMENT|7243,7248|false|false|false|C1546485|Diagnosis Type - Final|Final
Anatomy|Cell|SIMPLE_SEGMENT|7278,7294|false|false|false|C0014597|Epithelial Cells|epithelial cells
Anatomy|Cell|SIMPLE_SEGMENT|7289,7294|false|false|false|C0007634|Cells|cells
Event|Event|SIMPLE_SEGMENT|7300,7305|false|false|false|||field
Finding|Conceptual Entity|SIMPLE_SEGMENT|7300,7305|false|false|false|C1521738;C2346620;C2349184|Field;Force Field;Knowledge Field|field
Procedure|Health Care Activity|SIMPLE_SEGMENT|7300,7305|false|false|false|C1553496|field - patient encounter|field
Event|Event|SIMPLE_SEGMENT|7333,7338|false|false|false|||FIELD
Finding|Conceptual Entity|SIMPLE_SEGMENT|7333,7338|true|false|false|C1521738;C2346620;C2349184|Field;Force Field;Knowledge Field|FIELD
Procedure|Health Care Activity|SIMPLE_SEGMENT|7333,7338|true|false|false|C1553496|field - patient encounter|FIELD
Finding|Classification|SIMPLE_SEGMENT|7348,7356|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Finding|Finding|SIMPLE_SEGMENT|7348,7356|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7348,7356|false|false|false|C5237010|Expression Negative|NEGATIVE
Anatomy|Cell|SIMPLE_SEGMENT|7357,7360|false|false|false|C0206427|Rod Photoreceptors|ROD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7357,7360|true|false|false|C0035086|Renal Osteodystrophy|ROD
Event|Event|SIMPLE_SEGMENT|7357,7360|false|false|false|||ROD
Finding|Gene or Genome|SIMPLE_SEGMENT|7357,7360|true|false|false|C1424852|KNTC1 gene|ROD
Event|Event|SIMPLE_SEGMENT|7391,7396|false|false|false|||FIELD
Finding|Conceptual Entity|SIMPLE_SEGMENT|7391,7396|false|false|false|C1521738;C2346620;C2349184|Field;Force Field;Knowledge Field|FIELD
Procedure|Health Care Activity|SIMPLE_SEGMENT|7391,7396|false|false|false|C1553496|field - patient encounter|FIELD
Event|Event|SIMPLE_SEGMENT|7401,7408|false|false|false|||BUDDING
Finding|Cell Function|SIMPLE_SEGMENT|7401,7408|false|false|false|C1155616|Cell budding|BUDDING
Drug|Food|SIMPLE_SEGMENT|7409,7414|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Immunologic Factor|SIMPLE_SEGMENT|7409,7414|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|7409,7414|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7409,7414|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Event|Event|SIMPLE_SEGMENT|7409,7414|false|false|false|||YEAST
Event|Event|SIMPLE_SEGMENT|7423,7430|false|false|false|||QUALITY
Drug|Substance|SIMPLE_SEGMENT|7434,7442|false|false|false|C0370003|Specimen|SPECIMEN
Event|Event|SIMPLE_SEGMENT|7434,7442|false|false|false|||SPECIMEN
Finding|Body Substance|SIMPLE_SEGMENT|7434,7442|false|false|false|C1561495;C2347026|Biospecimen;Role Class - specimen|SPECIMEN
Finding|Functional Concept|SIMPLE_SEGMENT|7434,7442|false|false|false|C1561495;C2347026|Biospecimen;Role Class - specimen|SPECIMEN
Event|Event|SIMPLE_SEGMENT|7450,7452|false|false|false|||BE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7468,7479|false|false|false|C0231832|Respiratory rate|RESPIRATORY
Finding|Body Substance|SIMPLE_SEGMENT|7468,7479|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|RESPIRATORY
Finding|Functional Concept|SIMPLE_SEGMENT|7468,7479|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|RESPIRATORY
Finding|Intellectual Product|SIMPLE_SEGMENT|7468,7479|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|RESPIRATORY
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7468,7487|false|false|false|C4282127|Respiratory culture|RESPIRATORY CULTURE
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7480,7487|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|SIMPLE_SEGMENT|7480,7487|false|false|false|||CULTURE
Finding|Functional Concept|SIMPLE_SEGMENT|7480,7487|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|7480,7487|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7480,7487|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|SIMPLE_SEGMENT|7518,7528|false|false|false|||incubation
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7518,7528|false|false|false|C5453732|Incubation|incubation
Event|Event|SIMPLE_SEGMENT|7529,7537|false|false|false|||required
Event|Event|SIMPLE_SEGMENT|7541,7550|false|false|false|||determine
Event|Event|SIMPLE_SEGMENT|7555,7563|false|false|false|||presence
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7555,7563|false|false|false|C0392148|Providing presence (regime/therapy)|presence
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|7568,7575|false|false|false|C1689985|Absence (morphologic abnormality)|absence
Event|Event|SIMPLE_SEGMENT|7568,7575|false|false|false|||absence
Finding|Functional Concept|SIMPLE_SEGMENT|7568,7575|false|false|false|C0332197|Absent|absence
Finding|Functional Concept|SIMPLE_SEGMENT|7568,7578|false|false|false|C0332197|Absent|absence of
Finding|Functional Concept|SIMPLE_SEGMENT|7585,7594|false|false|false|C0231202|Symbiotic|commensal
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7595,7606|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|SIMPLE_SEGMENT|7595,7606|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|SIMPLE_SEGMENT|7595,7606|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|SIMPLE_SEGMENT|7595,7606|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Event|Event|SIMPLE_SEGMENT|7607,7612|false|false|false|||flora
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7621,7631|false|false|false|C0519030|Pneumonia due to Klebsiella pneumoniae|KLEBSIELLA
Event|Event|SIMPLE_SEGMENT|7621,7631|false|false|false|||KLEBSIELLA
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7621,7642|false|false|false|C2712605|Infection by Klebsiella pneumoniae in conditions classified elsewhere and of unspecified site|KLEBSIELLA PNEUMONIAE
Event|Event|SIMPLE_SEGMENT|7632,7642|false|false|false|||PNEUMONIAE
Event|Event|SIMPLE_SEGMENT|7654,7660|false|false|false|||GROWTH
Finding|Finding|SIMPLE_SEGMENT|7654,7660|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|7654,7660|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organism Function|SIMPLE_SEGMENT|7654,7660|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Physiologic Function|SIMPLE_SEGMENT|7654,7660|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|7654,7660|false|false|false|C2911660|Growth action|GROWTH
Drug|Antibiotic|SIMPLE_SEGMENT|7672,7681|false|false|false|C0007546|cefazolin|Cefazolin
Drug|Organic Chemical|SIMPLE_SEGMENT|7672,7681|false|false|false|C0007546|cefazolin|Cefazolin
Event|Event|SIMPLE_SEGMENT|7697,7705|false|false|false|||criteria
Finding|Idea or Concept|SIMPLE_SEGMENT|7697,7705|false|false|false|C0243161|criteria|criteria
Event|Event|SIMPLE_SEGMENT|7729,7736|false|false|false|||regimen
Finding|Intellectual Product|SIMPLE_SEGMENT|7729,7736|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7729,7736|false|false|false|C0040808|Treatment Protocols|regimen
Event|Event|SIMPLE_SEGMENT|7769,7773|false|false|false|||GRAM
Finding|Classification|SIMPLE_SEGMENT|7774,7782|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Finding|Finding|SIMPLE_SEGMENT|7774,7782|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7774,7782|false|false|false|C5237010|Expression Negative|NEGATIVE
Anatomy|Cell|SIMPLE_SEGMENT|7783,7786|false|false|false|C0206427|Rod Photoreceptors|ROD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7783,7786|false|false|false|C0035086|Renal Osteodystrophy|ROD
Event|Event|SIMPLE_SEGMENT|7783,7786|false|false|false|||ROD
Finding|Gene or Genome|SIMPLE_SEGMENT|7783,7786|false|false|false|C1424852|KNTC1 gene|ROD
Event|Event|SIMPLE_SEGMENT|7801,7807|false|false|false|||GROWTH
Finding|Finding|SIMPLE_SEGMENT|7801,7807|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|7801,7807|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organism Function|SIMPLE_SEGMENT|7801,7807|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Physiologic Function|SIMPLE_SEGMENT|7801,7807|false|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|7801,7807|false|false|false|C2911660|Growth action|GROWTH
Event|Event|SIMPLE_SEGMENT|7841,7854|false|false|false|||SENSITIVITIES
Finding|Finding|SIMPLE_SEGMENT|7841,7854|false|false|false|C0427965|Antimicrobial susceptibility|SENSITIVITIES
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7856,7859|false|false|false|C2732473|Ductal Carcinoma In Situ with Microinvasion|MIC
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|7856,7859|false|false|false|C0066256|methyl isocyanate|MIC
Drug|Organic Chemical|SIMPLE_SEGMENT|7856,7859|false|false|false|C0066256|methyl isocyanate|MIC
Event|Event|SIMPLE_SEGMENT|7856,7859|false|false|false|||MIC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7856,7859|false|false|false|C0281162;C0427978|Minimum Inhibitory Concentration Test;cisplatin/ifosfamide/mitomycin protocol|MIC
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7856,7859|false|false|false|C0281162;C0427978|Minimum Inhibitory Concentration Test;cisplatin/ifosfamide/mitomycin protocol|MIC
Event|Event|SIMPLE_SEGMENT|7874,7877|false|false|false|||MCG
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7991,8001|false|false|false|C0519030|Pneumonia due to Klebsiella pneumoniae|KLEBSIELLA
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7991,8012|false|false|false|C2712605|Infection by Klebsiella pneumoniae in conditions classified elsewhere and of unspecified site|KLEBSIELLA PNEUMONIAE
Event|Event|SIMPLE_SEGMENT|8002,8012|false|false|false|||PNEUMONIAE
Drug|Antibiotic|SIMPLE_SEGMENT|8047,8057|false|false|false|C0002680;C2095775|ampicillin;ampicillins|AMPICILLIN
Drug|Organic Chemical|SIMPLE_SEGMENT|8047,8057|false|false|false|C0002680;C2095775|ampicillin;ampicillins|AMPICILLIN
Event|Event|SIMPLE_SEGMENT|8047,8057|false|false|false|||AMPICILLIN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8047,8067|false|false|false|C2930041|Ampicillin / Sulbactam|AMPICILLIN/SULBACTAM
Drug|Antibiotic|SIMPLE_SEGMENT|8058,8067|false|false|false|C0038665|sulbactam|SULBACTAM
Drug|Organic Chemical|SIMPLE_SEGMENT|8058,8067|false|false|false|C0038665|sulbactam|SULBACTAM
Drug|Antibiotic|SIMPLE_SEGMENT|8078,8087|false|false|false|C0007546|cefazolin|CEFAZOLIN
Drug|Organic Chemical|SIMPLE_SEGMENT|8078,8087|false|false|false|C0007546|cefazolin|CEFAZOLIN
Drug|Antibiotic|SIMPLE_SEGMENT|8109,8117|false|false|false|C0055003|cefepime|CEFEPIME
Drug|Organic Chemical|SIMPLE_SEGMENT|8109,8117|false|false|false|C0055003|cefepime|CEFEPIME
Drug|Antibiotic|SIMPLE_SEGMENT|8140,8151|false|false|false|C0007559|ceftazidime|CEFTAZIDIME
Drug|Organic Chemical|SIMPLE_SEGMENT|8140,8151|false|false|false|C0007559|ceftazidime|CEFTAZIDIME
Drug|Antibiotic|SIMPLE_SEGMENT|8171,8182|false|false|false|C0007561|ceftriaxone|CEFTRIAXONE
Drug|Organic Chemical|SIMPLE_SEGMENT|8171,8182|false|false|false|C0007561|ceftriaxone|CEFTRIAXONE
Drug|Organic Chemical|SIMPLE_SEGMENT|8202,8215|false|false|false|C0008809|ciprofloxacin|CIPROFLOXACIN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8202,8215|false|false|false|C0008809|ciprofloxacin|CIPROFLOXACIN
Drug|Antibiotic|SIMPLE_SEGMENT|8233,8243|false|false|false|C3854019|gentamicin|GENTAMICIN
Drug|Organic Chemical|SIMPLE_SEGMENT|8233,8243|false|false|false|C3854019|gentamicin|GENTAMICIN
Event|Event|SIMPLE_SEGMENT|8233,8243|false|false|false|||GENTAMICIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8233,8243|false|false|false|C0202391|Gentamicin measurement|GENTAMICIN
Drug|Antibiotic|SIMPLE_SEGMENT|8264,8273|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|MEROPENEM
Drug|Clinical Drug|SIMPLE_SEGMENT|8264,8273|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|MEROPENEM
Drug|Organic Chemical|SIMPLE_SEGMENT|8264,8273|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|MEROPENEM
Drug|Antibiotic|SIMPLE_SEGMENT|8295,8307|false|false|false|C0031955|piperacillin|PIPERACILLIN
Drug|Organic Chemical|SIMPLE_SEGMENT|8295,8307|false|false|false|C0031955|piperacillin|PIPERACILLIN
Drug|Antibiotic|SIMPLE_SEGMENT|8308,8312|false|false|false|C0075870|tazobactam|TAZO
Drug|Organic Chemical|SIMPLE_SEGMENT|8308,8312|false|false|false|C0075870|tazobactam|TAZO
Drug|Antibiotic|SIMPLE_SEGMENT|8326,8336|false|false|false|C0040341|tobramycin|TOBRAMYCIN
Drug|Organic Chemical|SIMPLE_SEGMENT|8326,8336|false|false|false|C0040341|tobramycin|TOBRAMYCIN
Event|Event|SIMPLE_SEGMENT|8326,8336|false|false|false|||TOBRAMYCIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8326,8336|false|false|false|C0202490|Tobramycin measurement|TOBRAMYCIN
Drug|Antibiotic|SIMPLE_SEGMENT|8357,8369|false|false|false|C0041041|trimethoprim|TRIMETHOPRIM
Drug|Organic Chemical|SIMPLE_SEGMENT|8357,8369|false|false|false|C0041041|trimethoprim|TRIMETHOPRIM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8370,8375|false|false|false|C0749139|sulfa|SULFA
Finding|Intellectual Product|SIMPLE_SEGMENT|8391,8396|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|8397,8405|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8397,8412|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|8397,8412|false|false|false|C0489547|Hospital course|Hospital Course
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8436,8439|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|8436,8439|false|false|false|||HTN
Event|Event|SIMPLE_SEGMENT|8441,8444|false|false|false|||HLD
Event|Event|SIMPLE_SEGMENT|8446,8450|false|false|false|||DMII
Event|Event|SIMPLE_SEGMENT|8456,8459|false|false|false|||old
Event|Event|SIMPLE_SEGMENT|8463,8474|false|false|false|||transferred
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8488,8494|false|false|false|C4255010||NSTEMI
Event|Event|SIMPLE_SEGMENT|8488,8494|false|false|false|||NSTEMI
Finding|Finding|SIMPLE_SEGMENT|8488,8494|false|false|false|C3537184||NSTEMI
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8508,8514|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8508,8514|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8515,8522|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|8515,8522|false|false|false|||disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8527,8530|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8527,8530|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8527,8530|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|SIMPLE_SEGMENT|8527,8530|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|SIMPLE_SEGMENT|8527,8530|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8527,8530|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Event|Event|SIMPLE_SEGMENT|8527,8530|false|false|false|||DES
Finding|Gene or Genome|SIMPLE_SEGMENT|8527,8530|false|false|false|C1413980|DES gene|DES
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|8543,8552|false|false|false|C0001168|Complete obstruction|occlusion
Event|Event|SIMPLE_SEGMENT|8543,8552|false|false|false|||occlusion
Finding|Finding|SIMPLE_SEGMENT|8543,8552|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Functional Concept|SIMPLE_SEGMENT|8543,8552|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|8543,8552|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Pathologic Function|SIMPLE_SEGMENT|8543,8552|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Event|Event|SIMPLE_SEGMENT|8553,8558|false|false|false|||found
Finding|Finding|SIMPLE_SEGMENT|8567,8573|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|8567,8573|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8613,8619|false|false|false|C4255010||NSTEMI
Event|Event|SIMPLE_SEGMENT|8613,8619|false|false|false|||NSTEMI
Finding|Finding|SIMPLE_SEGMENT|8613,8619|false|false|false|C3537184||NSTEMI
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8621,8627|false|false|false|C4255010||NSTEMI
Event|Event|SIMPLE_SEGMENT|8621,8627|false|false|false|||NSTEMI
Finding|Finding|SIMPLE_SEGMENT|8621,8627|false|false|false|C3537184||NSTEMI
Event|Event|SIMPLE_SEGMENT|8637,8640|false|false|false|||STE
Finding|Gene or Genome|SIMPLE_SEGMENT|8637,8640|false|false|false|C1420459;C3811127|SULT1E1 gene;SULT1E1 wt Allele|STE
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8663,8674|false|false|false|C0011570|Mental Depression|depressions
Event|Event|SIMPLE_SEGMENT|8663,8674|false|false|false|||depressions
Finding|Idea or Concept|SIMPLE_SEGMENT|8679,8690|false|false|false|C0750502|Significant|significant
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8697,8703|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8697,8703|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8704,8711|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|8704,8711|false|false|false|||disease
Finding|Idea or Concept|SIMPLE_SEGMENT|8716,8727|false|true|false|C0750502|Significant|significant
Event|Event|SIMPLE_SEGMENT|8728,8736|false|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|8728,8736|false|true|false|C1261287|Stenosis|stenosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8740,8743|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8740,8743|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|SIMPLE_SEGMENT|8740,8743|false|false|false|||LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|8740,8743|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8749,8752|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8749,8752|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8749,8752|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|SIMPLE_SEGMENT|8749,8752|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|SIMPLE_SEGMENT|8749,8752|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8749,8752|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Event|Event|SIMPLE_SEGMENT|8749,8752|false|false|false|||DES
Finding|Gene or Genome|SIMPLE_SEGMENT|8749,8752|false|false|false|C1413980|DES gene|DES
Finding|Finding|SIMPLE_SEGMENT|8758,8766|false|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Finding|Functional Concept|SIMPLE_SEGMENT|8758,8766|false|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Event|Event|SIMPLE_SEGMENT|8767,8776|false|false|false|||diagnonal
Finding|Functional Concept|SIMPLE_SEGMENT|8778,8784|false|false|false|C0205341;C1705914|Repeat;Repeat Object|Repeat
Event|Event|SIMPLE_SEGMENT|8785,8789|false|false|false|||cath
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8785,8789|false|false|false|C0007430|Catheterization|cath
Event|Event|SIMPLE_SEGMENT|8790,8799|false|false|false|||unchanged
Finding|Finding|SIMPLE_SEGMENT|8790,8799|false|false|false|C0442739||unchanged
Event|Event|SIMPLE_SEGMENT|8809,8816|false|false|false|||started
Drug|Organic Chemical|SIMPLE_SEGMENT|8820,8826|false|false|false|C0633084|Plavix|plavix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8820,8826|false|false|false|C0633084|Plavix|plavix
Event|Event|SIMPLE_SEGMENT|8820,8826|false|false|false|||plavix
Drug|Organic Chemical|SIMPLE_SEGMENT|8828,8840|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8828,8840|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|SIMPLE_SEGMENT|8828,8840|false|false|false|||atorvastatin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8842,8845|false|false|false|C1452534|ACE protein, human|ACE
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8842,8845|false|false|false|C1452534|ACE protein, human|ACE
Event|Event|SIMPLE_SEGMENT|8842,8845|false|false|false|||ACE
Finding|Gene or Genome|SIMPLE_SEGMENT|8842,8845|false|false|false|C1413931;C4284014|ACE gene;Adverse Childhood Experience questionnaire|ACE
Finding|Intellectual Product|SIMPLE_SEGMENT|8842,8845|false|false|false|C1413931;C4284014|ACE gene;Adverse Childhood Experience questionnaire|ACE
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8842,8845|false|false|false|C0050385;C0108844;C0279078;C1879921|CDE Regimen;CDE protocol;cisplatin, cytarabine, and etoposide chemotherapy protocol;cyclophosphamide/doxorubicin protocol|ACE
Drug|Organic Chemical|SIMPLE_SEGMENT|8853,8863|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8853,8863|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|SIMPLE_SEGMENT|8853,8863|false|false|false|||metoprolol
Procedure|Health Care Activity|SIMPLE_SEGMENT|8865,8869|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|Echo
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8865,8869|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|Echo
Event|Event|SIMPLE_SEGMENT|8871,8877|false|false|false|||showed
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8878,8882|false|false|false|C0428772|Left ventricular ejection fraction|LVEF
Event|Event|SIMPLE_SEGMENT|8878,8882|false|false|false|||LVEF
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8878,8882|false|false|false|C3837267|LVEF (procedure)|LVEF
Event|Event|SIMPLE_SEGMENT|8895,8906|false|false|false|||hypokinesis
Finding|Finding|SIMPLE_SEGMENT|8895,8906|false|false|false|C0086439|Hypokinesia|hypokinesis
Event|Event|SIMPLE_SEGMENT|8924,8932|false|false|false|||segments
Anatomy|Cell Component|SIMPLE_SEGMENT|8938,8942|false|false|false|C3890171|dinoflagellate apex|apex
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8938,8942|false|false|false|C0140145|APEX1 protein, human|apex
Drug|Enzyme|SIMPLE_SEGMENT|8938,8942|false|false|false|C0140145|APEX1 protein, human|apex
Finding|Gene or Genome|SIMPLE_SEGMENT|8938,8942|false|false|false|C1332102|APEX1 gene|apex
Event|Event|SIMPLE_SEGMENT|8951,8958|false|false|false|||started
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8959,8970|false|false|false|C0851145|on warfarin|on warfarin
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|8962,8970|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|SIMPLE_SEGMENT|8962,8970|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8962,8970|false|false|false|C0043031|warfarin|warfarin
Event|Event|SIMPLE_SEGMENT|8962,8970|false|false|false|||warfarin
Event|Event|SIMPLE_SEGMENT|8979,8990|false|false|false|||hypokinetic
Finding|Finding|SIMPLE_SEGMENT|8979,8990|false|false|false|C0086439|Hypokinesia|hypokinetic
Event|Event|SIMPLE_SEGMENT|8998,9002|false|false|false|||well
Finding|Finding|SIMPLE_SEGMENT|8998,9002|false|false|false|C5575035|Well (answer to question)|well
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9010,9016|false|false|false|C0018792|Heart Atrium|atrial
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9010,9029|false|false|false|C2926591||atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9010,9029|false|false|false|C0004238|Atrial Fibrillation|atrial fibrillation
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|9010,9029|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9017,9029|false|false|false|C0232197|Fibrillation|fibrillation
Event|Event|SIMPLE_SEGMENT|9017,9029|false|false|false|||fibrillation
Event|Event|SIMPLE_SEGMENT|9033,9042|false|false|false|||discussed
Finding|Finding|SIMPLE_SEGMENT|9057,9065|false|false|false|C0332149|Possible|Possibly
Event|Event|SIMPLE_SEGMENT|9103,9108|false|false|false|||mixed
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9109,9115|false|false|false|C0042449|Veins|venous
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9133,9137|false|false|false|C0034094|Pulmonary Wedge Pressure|PCWP
Event|Event|SIMPLE_SEGMENT|9133,9137|false|false|false|||PCWP
Event|Event|SIMPLE_SEGMENT|9155,9163|false|false|false|||required
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9164,9172|false|false|false|C0237795|Pressors|pressors
Event|Event|SIMPLE_SEGMENT|9164,9172|false|false|false|||pressors
Event|Event|SIMPLE_SEGMENT|9177,9184|false|false|false|||balloon
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9177,9184|false|false|false|C0004704|Balloon Dilatation|balloon
Event|Event|SIMPLE_SEGMENT|9186,9190|false|false|false|||pump
Finding|Molecular Function|SIMPLE_SEGMENT|9186,9190|false|false|false|C1150186|matrix metalloproteinase 7 activity|pump
Finding|Intellectual Product|SIMPLE_SEGMENT|9199,9203|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|SIMPLE_SEGMENT|9217,9223|false|false|false|||weaned
Event|Event|SIMPLE_SEGMENT|9237,9245|false|false|false|||remained
Finding|Finding|SIMPLE_SEGMENT|9247,9269|false|false|false|C0578150|Hemodynamically stable|hemodynamically stable
Event|Event|SIMPLE_SEGMENT|9263,9269|false|false|false|||stable
Finding|Intellectual Product|SIMPLE_SEGMENT|9263,9269|false|false|false|C1547311|Patient Condition Code - Stable|stable
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9277,9281|false|false|false|C1742913|REST protein, human|rest
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9277,9281|false|false|false|C1742913|REST protein, human|rest
Event|Event|SIMPLE_SEGMENT|9277,9281|false|false|false|||rest
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|9277,9281|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Gene or Genome|SIMPLE_SEGMENT|9277,9281|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Molecular Function|SIMPLE_SEGMENT|9277,9281|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Idea or Concept|SIMPLE_SEGMENT|9285,9293|false|false|false|C1547192|Organization unit type - Hospital|hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9285,9300|false|false|false|C0488549||hospital course
Finding|Finding|SIMPLE_SEGMENT|9285,9300|false|false|false|C0489547|Hospital course|hospital course
Event|Event|SIMPLE_SEGMENT|9294,9300|false|false|false|||course
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9306,9312|false|false|false|C0018792|Heart Atrium|Atrial
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9306,9325|false|false|false|C2926591||Atrial Fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9306,9325|false|false|false|C0004238|Atrial Fibrillation|Atrial Fibrillation
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|9306,9325|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Atrial Fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9313,9325|false|false|false|C0232197|Fibrillation|Fibrillation
Event|Event|SIMPLE_SEGMENT|9313,9325|false|false|false|||Fibrillation
Finding|Body Substance|SIMPLE_SEGMENT|9326,9333|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|9326,9333|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|9326,9333|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|9350,9357|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|9350,9357|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|9350,9357|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|9350,9357|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|9350,9360|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9372,9376|false|false|false|C0004238|Atrial Fibrillation|afib
Event|Event|SIMPLE_SEGMENT|9372,9376|false|false|false|||afib
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|9372,9376|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|afib
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9385,9388|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9385,9388|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|9385,9388|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9385,9388|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|9385,9388|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|9385,9388|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|9385,9388|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9385,9388|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|9385,9388|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|9385,9388|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|9385,9388|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|SIMPLE_SEGMENT|9407,9417|false|false|false|||maintained
Drug|Organic Chemical|SIMPLE_SEGMENT|9421,9428|false|false|false|C0012265|digoxin|digoxin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9421,9428|false|false|false|C0012265|digoxin|digoxin
Event|Event|SIMPLE_SEGMENT|9421,9428|false|false|false|||digoxin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9421,9428|false|false|false|C0337449|Digoxin measurement|digoxin
Finding|Finding|SIMPLE_SEGMENT|9432,9436|false|false|false|C5575035|Well (answer to question)|well
Drug|Organic Chemical|SIMPLE_SEGMENT|9440,9447|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9440,9447|false|false|false|C0004057|aspirin|aspirin
Event|Event|SIMPLE_SEGMENT|9440,9447|false|false|false|||aspirin
Event|Event|SIMPLE_SEGMENT|9455,9457|false|false|false|||PO
Event|Event|SIMPLE_SEGMENT|9473,9482|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|9473,9482|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|9492,9497|false|false|false|||found
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9507,9513|false|false|false|C0018792|Heart Atrium|atrial
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9515,9527|false|false|false|C0232197|Fibrillation|fibrillation
Event|Event|SIMPLE_SEGMENT|9515,9527|false|false|false|||fibrillation
Event|Event|SIMPLE_SEGMENT|9535,9544|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|9535,9544|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|9553,9561|false|false|false|||decision
Finding|Mental Process|SIMPLE_SEGMENT|9553,9561|false|false|false|C0679006|Decision|decision
Event|Event|SIMPLE_SEGMENT|9575,9588|false|false|false|||anticoagulate
Drug|Organic Chemical|SIMPLE_SEGMENT|9594,9602|false|false|false|C0699129|Coumadin|Coumadin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9594,9602|false|false|false|C0699129|Coumadin|Coumadin
Event|Event|SIMPLE_SEGMENT|9594,9602|false|false|false|||Coumadin
Event|Event|SIMPLE_SEGMENT|9612,9621|false|false|false|||continued
Finding|Idea or Concept|SIMPLE_SEGMENT|9625,9629|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|9625,9629|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|9625,9629|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|9630,9634|false|false|false|||dose
Drug|Organic Chemical|SIMPLE_SEGMENT|9636,9643|false|false|false|C0012265|digoxin|digoxin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9636,9643|false|false|false|C0012265|digoxin|digoxin
Event|Event|SIMPLE_SEGMENT|9636,9643|false|false|false|||digoxin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9636,9643|false|false|false|C0337449|Digoxin measurement|digoxin
Finding|Idea or Concept|SIMPLE_SEGMENT|9650,9654|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|9650,9654|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|9650,9654|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|9660,9667|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9660,9667|false|false|false|C0004057|aspirin|aspirin
Event|Event|SIMPLE_SEGMENT|9660,9667|false|false|false|||aspirin
Event|Event|SIMPLE_SEGMENT|9672,9681|false|false|false|||decreased
Event|Event|SIMPLE_SEGMENT|9685,9694|false|false|false|||discussed
Finding|Idea or Concept|SIMPLE_SEGMENT|9695,9700|false|false|false|C1552828|Table Frame - above|above
Event|Event|SIMPLE_SEGMENT|9707,9717|false|false|false|||initiation
Finding|Functional Concept|SIMPLE_SEGMENT|9707,9717|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Finding|Genetic Function|SIMPLE_SEGMENT|9707,9717|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Finding|Mental Process|SIMPLE_SEGMENT|9707,9717|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Drug|Organic Chemical|SIMPLE_SEGMENT|9721,9729|false|false|false|C0699129|Coumadin|Coumadin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9721,9729|false|false|false|C0699129|Coumadin|Coumadin
Event|Event|SIMPLE_SEGMENT|9721,9729|false|false|false|||Coumadin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9734,9743|false|false|false|C0018965|Hematuria|Hematuria
Event|Event|SIMPLE_SEGMENT|9734,9743|false|false|false|||Hematuria
Finding|Finding|SIMPLE_SEGMENT|9746,9752|false|true|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Idea or Concept|SIMPLE_SEGMENT|9746,9752|false|true|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Event|Event|SIMPLE_SEGMENT|9753,9762|false|false|false|||traumatic
Finding|Functional Concept|SIMPLE_SEGMENT|9753,9762|false|true|false|C0332663|Traumatic|traumatic
Finding|Functional Concept|SIMPLE_SEGMENT|9777,9785|false|false|false|C0205373;C5849094|Systemic;Systemic Route of Administration|systemic
Event|Event|SIMPLE_SEGMENT|9786,9801|false|false|false|||anticoagulation
Finding|Finding|SIMPLE_SEGMENT|9786,9801|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|SIMPLE_SEGMENT|9786,9801|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9786,9801|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Finding|Body Substance|SIMPLE_SEGMENT|9807,9814|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|9807,9814|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|9807,9814|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|9815,9821|false|false|false|||pulled
Event|Event|SIMPLE_SEGMENT|9830,9838|false|false|false|||Cytology
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9830,9838|false|false|false|C0010818;C1305671|Cytological Techniques;Cytology--Technique|Cytology
Event|Event|SIMPLE_SEGMENT|9843,9851|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|9843,9851|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|9843,9851|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|9843,9851|false|false|false|C5237010|Expression Negative|negative
Event|Event|SIMPLE_SEGMENT|9861,9869|false|false|false|||followup
Event|Event|SIMPLE_SEGMENT|9871,9881|false|false|false|||outpatient
Finding|Classification|SIMPLE_SEGMENT|9871,9881|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|9871,9881|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|SIMPLE_SEGMENT|9887,9894|false|false|false|||urology
Finding|Finding|SIMPLE_SEGMENT|9899,9906|false|false|false|C0013404;C2024878|Dyspnea|Dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|9899,9906|false|false|false|C0013404;C2024878|Dyspnea|Dyspnea
Finding|Body Substance|SIMPLE_SEGMENT|9909,9916|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|9909,9916|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|9909,9916|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|9921,9926|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|SIMPLE_SEGMENT|9927,9935|false|false|false|||episodes
Event|Event|SIMPLE_SEGMENT|9939,9946|false|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|9939,9946|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|9939,9946|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Event|Event|SIMPLE_SEGMENT|9966,9976|false|false|false|||attributed
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9980,9989|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9980,9989|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|9980,9989|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|9980,9995|false|false|false|C0034063|Pulmonary Edema|pulmonary edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9990,9995|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|9990,9995|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|9990,9995|false|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|10000,10008|false|false|false|||improved
Finding|Finding|SIMPLE_SEGMENT|10000,10008|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Finding|Intellectual Product|SIMPLE_SEGMENT|10000,10008|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Event|Event|SIMPLE_SEGMENT|10014,10022|false|false|false|||diruesis
Event|Event|SIMPLE_SEGMENT|10040,10043|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10040,10043|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|SIMPLE_SEGMENT|10044,10050|false|false|false|||showed
Finding|Finding|SIMPLE_SEGMENT|10051,10059|false|false|false|C0332149|Possible|possible
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10060,10073|false|true|false|C0521530|Lung consolidation|consolidation
Event|Event|SIMPLE_SEGMENT|10060,10073|false|false|false|||consolidation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10077,10080|false|false|false|C1261074|Structure of right upper lobe of lung|RUL
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|10098,10108|false|false|false|C1720922|Respiratory Aspiration|aspiration
Event|Event|SIMPLE_SEGMENT|10098,10108|false|false|false|||aspiration
Finding|Finding|SIMPLE_SEGMENT|10098,10108|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|aspiration
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|10098,10108|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|aspiration
Finding|Pathologic Function|SIMPLE_SEGMENT|10098,10108|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|aspiration
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10098,10108|false|false|false|C0349707||aspiration
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10098,10118|false|false|false|C0032290;C1761609|Aspiration Pneumonia;Aspiration pneumonitis|aspiration pneumonia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10109,10118|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|SIMPLE_SEGMENT|10109,10118|false|false|false|||pneumonia
Event|Event|SIMPLE_SEGMENT|10129,10138|false|false|false|||treatment
Finding|Conceptual Entity|SIMPLE_SEGMENT|10129,10138|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|SIMPLE_SEGMENT|10129,10138|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|SIMPLE_SEGMENT|10129,10138|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10129,10138|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Event|Event|SIMPLE_SEGMENT|10144,10152|false|false|false|||deferred
Event|Event|SIMPLE_SEGMENT|10178,10183|false|false|false|||signs
Finding|Finding|SIMPLE_SEGMENT|10178,10183|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|10178,10183|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10187,10197|false|false|false|C0009450|Communicable Diseases|infectious
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|10198,10201|false|false|false|C0600500|Peptide Nucleic Acids|pna
Event|Event|SIMPLE_SEGMENT|10198,10201|false|false|false|||pna
Finding|Body Substance|SIMPLE_SEGMENT|10217,10223|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Finding|Intellectual Product|SIMPLE_SEGMENT|10217,10223|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Event|Event|SIMPLE_SEGMENT|10224,10232|false|false|false|||cultures
Finding|Idea or Concept|SIMPLE_SEGMENT|10224,10232|false|true|false|C0010453|Culture (Anthropological)|cultures
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10244,10254|false|false|false|C0519030|Pneumonia due to Klebsiella pneumoniae|Klebsiella
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10244,10264|false|false|false|C0519030|Pneumonia due to Klebsiella pneumoniae|Klebsiella pneumonia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10255,10264|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|SIMPLE_SEGMENT|10255,10264|false|false|false|||pneumonia
Event|Event|SIMPLE_SEGMENT|10273,10283|false|false|false|||discussion
Finding|Social Behavior|SIMPLE_SEGMENT|10273,10283|false|false|false|C2584313|Discussion (communication)|discussion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10273,10283|false|false|false|C0557061|Discussion (procedure)|discussion
Event|Event|SIMPLE_SEGMENT|10293,10297|false|false|false|||felt
Event|Event|SIMPLE_SEGMENT|10311,10318|false|false|false|||warrant
Event|Event|SIMPLE_SEGMENT|10323,10332|false|false|false|||treatment
Finding|Conceptual Entity|SIMPLE_SEGMENT|10323,10332|true|false|true|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|SIMPLE_SEGMENT|10323,10332|true|false|true|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|SIMPLE_SEGMENT|10323,10332|true|false|true|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10323,10332|true|false|true|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Event|Event|SIMPLE_SEGMENT|10344,10356|false|false|false|||asymptomatic
Finding|Finding|SIMPLE_SEGMENT|10344,10356|false|false|false|C0231221;C0332151|Asymptomatic (finding);Asymptomatic diagnosis of|asymptomatic
Event|Event|SIMPLE_SEGMENT|10366,10376|false|false|false|||discharged
Drug|Organic Chemical|SIMPLE_SEGMENT|10383,10388|false|false|false|C0699992|Lasix|lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10383,10388|false|false|false|C0699992|Lasix|lasix
Finding|Idea or Concept|SIMPLE_SEGMENT|10407,10411|false|false|false|C1552851|next - HtmlLinkType|next
Drug|Inorganic Chemical|SIMPLE_SEGMENT|10412,10424|false|false|false|C0013832;C3536863|Electrolyte [EPC];Electrolytes|electrolytes
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10412,10424|false|false|false|C0013832;C3536863|Electrolyte [EPC];Electrolytes|electrolytes
Event|Event|SIMPLE_SEGMENT|10412,10424|false|false|false|||electrolytes
Event|Event|SIMPLE_SEGMENT|10431,10438|false|false|false|||checked
Event|Event|SIMPLE_SEGMENT|10457,10463|false|false|false|||severe
Finding|Finding|SIMPLE_SEGMENT|10457,10463|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|10457,10463|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Sign or Symptom|SIMPLE_SEGMENT|10470,10481|false|false|false|C2129214|Loose stool|loose stool
Event|Event|SIMPLE_SEGMENT|10476,10481|false|false|false|||stool
Finding|Body Substance|SIMPLE_SEGMENT|10476,10481|false|true|false|C0015733|Feces|stool
Event|Event|SIMPLE_SEGMENT|10485,10492|false|false|false|||setting
Finding|Mental Process|SIMPLE_SEGMENT|10485,10492|false|false|false|C0542559|contextual factors|setting
Drug|Antibiotic|SIMPLE_SEGMENT|10496,10506|false|false|false|C0003232|Antibiotics|antibiotic
Event|Event|SIMPLE_SEGMENT|10534,10544|false|false|false|||outpatient
Finding|Classification|SIMPLE_SEGMENT|10534,10544|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|10534,10544|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Anatomy|Cell|SIMPLE_SEGMENT|10553,10556|false|false|false|C0023516|Leukocytes|WBC
Event|Event|SIMPLE_SEGMENT|10553,10556|false|false|false|||WBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10567,10570|false|false|false|C1114365||age
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10567,10570|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|SIMPLE_SEGMENT|10567,10570|false|false|false|C0162574|Glycation End Products, Advanced|age
Event|Event|SIMPLE_SEGMENT|10567,10570|false|false|false|||age
Event|Event|SIMPLE_SEGMENT|10576,10583|false|false|false|||treated
Event|Event|SIMPLE_SEGMENT|10588,10594|false|false|false|||severe
Finding|Finding|SIMPLE_SEGMENT|10588,10594|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|10588,10594|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Body Substance|SIMPLE_SEGMENT|10596,10603|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|10596,10603|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|10596,10603|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|10608,10615|false|false|false|||started
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10619,10629|false|false|false|C0042313|vancomycin|vancomycin
Drug|Antibiotic|SIMPLE_SEGMENT|10619,10629|false|false|false|C0042313|vancomycin|vancomycin
Event|Event|SIMPLE_SEGMENT|10619,10629|false|false|false|||vancomycin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10619,10629|false|false|false|C0489941|Vancomycin measurement|vancomycin
Finding|Idea or Concept|SIMPLE_SEGMENT|10651,10654|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|10651,10654|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Idea or Concept|SIMPLE_SEGMENT|10663,10666|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|10663,10666|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Idea or Concept|SIMPLE_SEGMENT|10677,10680|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|10677,10680|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Anatomy|Body Location or Region|SIMPLE_SEGMENT|10691,10707|false|false|false|C0744316|gastroesophageal|GASTROESOPHAGEAL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10691,10714|false|false|false|C0017168|Gastroesophageal reflux disease|GASTROESOPHAGEAL REFLUX
Finding|Finding|SIMPLE_SEGMENT|10691,10714|false|false|false|C3813607;C4317146|Acid reflux;Infantile Gastroesophageal Reflux|GASTROESOPHAGEAL REFLUX
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10691,10722|false|false|false|C0017168|Gastroesophageal reflux disease|GASTROESOPHAGEAL REFLUX DISEASE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10691,10729|false|false|false|C0017168|Gastroesophageal reflux disease|GASTROESOPHAGEAL REFLUX DISEASE (GERD)
Event|Event|SIMPLE_SEGMENT|10708,10714|false|false|false|||REFLUX
Finding|Pathologic Function|SIMPLE_SEGMENT|10708,10714|false|false|false|C0232483|Reflux|REFLUX
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10715,10722|false|false|false|C0012634|Disease|DISEASE
Event|Event|SIMPLE_SEGMENT|10715,10722|false|false|false|||DISEASE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10724,10728|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|SIMPLE_SEGMENT|10724,10728|false|false|false|||GERD
Event|Event|SIMPLE_SEGMENT|10732,10741|false|false|false|||Endoscopy
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10732,10741|false|false|false|C0014245;C0079278|Endoscopy (procedure);Endoscopy, Gastrointestinal|Endoscopy
Event|Event|SIMPLE_SEGMENT|10742,10751|false|false|false|||confirmed
Event|Event|SIMPLE_SEGMENT|10761,10768|false|false|false|||treated
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10774,10777|false|false|false|C0358591|Proton Pump Inhibitors|PPI
Event|Event|SIMPLE_SEGMENT|10774,10777|false|false|false|||PPI
Finding|Physiologic Function|SIMPLE_SEGMENT|10774,10777|false|false|false|C0871125|Prepulse Inhibition|PPI
Drug|Antibiotic|SIMPLE_SEGMENT|10781,10795|false|false|false|C0055856|clarithromycin|clarithromycin
Drug|Organic Chemical|SIMPLE_SEGMENT|10781,10795|false|false|false|C0055856|clarithromycin|clarithromycin
Event|Event|SIMPLE_SEGMENT|10781,10795|false|false|false|||clarithromycin
Drug|Antibiotic|SIMPLE_SEGMENT|10796,10807|false|false|false|C0002645|amoxicillin|amoxicillin
Drug|Organic Chemical|SIMPLE_SEGMENT|10796,10807|false|false|false|C0002645|amoxicillin|amoxicillin
Event|Event|SIMPLE_SEGMENT|10796,10807|false|false|false|||amoxicillin
Drug|Organic Chemical|SIMPLE_SEGMENT|10831,10841|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10831,10841|false|false|false|C0028978|omeprazole|Omeprazole
Event|Event|SIMPLE_SEGMENT|10847,10856|false|false|false|||continued
Drug|Antibiotic|SIMPLE_SEGMENT|10858,10869|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|Antibiotics
Event|Event|SIMPLE_SEGMENT|10858,10869|false|false|false|||Antibiotics
Event|Event|SIMPLE_SEGMENT|10870,10874|false|false|false|||held
Finding|Mental Process|SIMPLE_SEGMENT|10878,10885|false|false|false|C0542559|contextual factors|setting
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10889,10905|false|false|false|C0343386|Clostridium difficile infection|c.diff infection
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10896,10905|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|10896,10905|false|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|10896,10905|false|false|false|C3714514|Infection|infection
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|10911,10919|false|false|false|C0011206|Delirium|Delirium
Event|Event|SIMPLE_SEGMENT|10911,10919|false|false|false|||Delirium
Finding|Body Substance|SIMPLE_SEGMENT|10922,10929|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|10922,10929|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|10922,10929|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|10944,10954|false|false|false|C1142436|Sundowning|sundowning
Event|Event|SIMPLE_SEGMENT|10944,10954|false|false|false|||sundowning
Event|Event|SIMPLE_SEGMENT|10962,10977|false|false|false|||hospitalization
Procedure|Health Care Activity|SIMPLE_SEGMENT|10962,10977|false|false|false|C0019993|Hospitalization|hospitalization
Event|Event|SIMPLE_SEGMENT|10979,10988|false|false|false|||requiring
Drug|Organic Chemical|SIMPLE_SEGMENT|10989,10997|false|false|false|C0287163|Seroquel|Seroquel
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10989,10997|false|false|false|C0287163|Seroquel|Seroquel
Finding|Intellectual Product|SIMPLE_SEGMENT|11003,11010|false|false|false|C1547296|Chronic - Admission Level of Care Code|CHRONIC
Procedure|Health Care Activity|SIMPLE_SEGMENT|11003,11010|false|false|false|C1555457|Provision of recurring care for chronic illness|CHRONIC
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|11036,11051|false|false|false|C0037944;C1861329|Spinal Stenosis;Spinal canal stenosis|Spinal Stenosis
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|11036,11051|false|false|false|C0037944;C1861329|Spinal Stenosis;Spinal canal stenosis|Spinal Stenosis
Event|Event|SIMPLE_SEGMENT|11043,11051|false|false|false|||Stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|11043,11051|false|false|false|C1261287|Stenosis|Stenosis
Drug|Organic Chemical|SIMPLE_SEGMENT|11063,11073|false|false|false|C0060926|gabapentin|gabapentin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11063,11073|false|false|false|C0060926|gabapentin|gabapentin
Event|Event|SIMPLE_SEGMENT|11063,11073|false|false|false|||gabapentin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11077,11080|false|false|false|C0011989;C4551571|Camurati-Engelmann Syndrome;Cranioectodermal dysplasia|ced
Drug|Antibiotic|SIMPLE_SEGMENT|11077,11080|false|false|false|C0007738|cephradine|ced
Drug|Organic Chemical|SIMPLE_SEGMENT|11077,11080|false|false|false|C0007738|cephradine|ced
Event|Event|SIMPLE_SEGMENT|11077,11080|false|false|false|||ced
Finding|Functional Concept|SIMPLE_SEGMENT|11077,11080|false|false|false|C1366557;C1704974;C3890738|Convection-Enhanced Delivery;TGFB1 gene;TGFB1 wt Allele|ced
Finding|Gene or Genome|SIMPLE_SEGMENT|11077,11080|false|false|false|C1366557;C1704974;C3890738|Convection-Enhanced Delivery;TGFB1 gene;TGFB1 wt Allele|ced
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11077,11080|false|false|false|C0108844;C0280001|CDE protocol;cisplatin/dexamethasone/etoposide protocol|ced
Drug|Organic Chemical|SIMPLE_SEGMENT|11081,11089|false|false|false|C0027396|naproxen|naproxen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11081,11089|false|false|false|C0027396|naproxen|naproxen
Event|Event|SIMPLE_SEGMENT|11081,11089|false|false|false|||naproxen
Event|Event|SIMPLE_SEGMENT|11101,11109|false|false|false|||complain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11113,11117|false|true|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|11113,11117|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|11113,11117|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|11113,11117|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Idea or Concept|SIMPLE_SEGMENT|11129,11137|false|false|false|C1547192|Organization unit type - Hospital|hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11129,11144|true|false|false|C0488549||hospital course
Finding|Finding|SIMPLE_SEGMENT|11129,11144|true|false|false|C0489547|Hospital course|hospital course
Event|Event|SIMPLE_SEGMENT|11138,11144|false|false|false|||course
Event|Event|SIMPLE_SEGMENT|11172,11176|false|false|false|||take
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11186,11192|false|true|false|C0003211;C0358845|Analgesics and non-steroidal anti-inflammatory drugs;Anti-Inflammatory Agents, Non-Steroidal|NSAIDS
Event|Event|SIMPLE_SEGMENT|11186,11192|false|false|false|||NSAIDS
Event|Event|SIMPLE_SEGMENT|11196,11203|false|false|false|||setting
Finding|Mental Process|SIMPLE_SEGMENT|11196,11203|false|false|false|C0542559|contextual factors|setting
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|11214,11217|false|false|false|C0262187|anterior calcarine sulcus (human only)|ACS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11214,11217|false|false|false|C0742343;C0796147|Acrocallosal Syndrome;Acute Chest Syndrome|ACS
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11214,11217|false|false|false|C4042561|ACSS2 protein, human|ACS
Drug|Enzyme|SIMPLE_SEGMENT|11214,11217|false|false|false|C4042561|ACSS2 protein, human|ACS
Event|Event|SIMPLE_SEGMENT|11214,11217|false|false|false|||ACS
Finding|Gene or Genome|SIMPLE_SEGMENT|11214,11217|false|false|false|C1150760;C1424787;C1825842;C1842089;C2266615;C4318612;C5400867;C5551036|ACCS gene;ACS - Activity Card Sort;ACSS2 gene;ACSS2 wt Allele;American Community Survey;CO-methylating acetyl-CoA synthase activity;PLA2G15 gene;acetate-CoA ligase activity|ACS
Finding|Intellectual Product|SIMPLE_SEGMENT|11214,11217|false|false|false|C1150760;C1424787;C1825842;C1842089;C2266615;C4318612;C5400867;C5551036|ACCS gene;ACS - Activity Card Sort;ACSS2 gene;ACSS2 wt Allele;American Community Survey;CO-methylating acetyl-CoA synthase activity;PLA2G15 gene;acetate-CoA ligase activity|ACS
Finding|Molecular Function|SIMPLE_SEGMENT|11214,11217|false|false|false|C1150760;C1424787;C1825842;C1842089;C2266615;C4318612;C5400867;C5551036|ACCS gene;ACS - Activity Card Sort;ACSS2 gene;ACSS2 wt Allele;American Community Survey;CO-methylating acetyl-CoA synthase activity;PLA2G15 gene;acetate-CoA ligase activity|ACS
Drug|Organic Chemical|SIMPLE_SEGMENT|11230,11238|false|false|false|C0699129|Coumadin|Coumadin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11230,11238|false|false|false|C0699129|Coumadin|Coumadin
Drug|Organic Chemical|SIMPLE_SEGMENT|11240,11246|false|false|false|C0633084|Plavix|Plavix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11240,11246|false|false|false|C0633084|Plavix|Plavix
Event|Event|SIMPLE_SEGMENT|11240,11246|false|false|false|||Plavix
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11251,11254|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|asa
Drug|Enzyme|SIMPLE_SEGMENT|11251,11254|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|asa
Drug|Organic Chemical|SIMPLE_SEGMENT|11251,11254|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|asa
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11251,11254|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|asa
Event|Event|SIMPLE_SEGMENT|11251,11254|false|false|false|||asa
Finding|Gene or Genome|SIMPLE_SEGMENT|11251,11254|false|false|false|C1412553|ARSA gene|asa
Event|Event|SIMPLE_SEGMENT|11263,11273|false|false|false|||maintained
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|11277,11280|false|false|false|C1845118|SHORT STATURE, IDIOPATHIC, X-LINKED|ISS
Event|Event|SIMPLE_SEGMENT|11277,11280|false|false|false|||ISS
Event|Event|SIMPLE_SEGMENT|11288,11297|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|11288,11297|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|11302,11312|false|false|false|||discharged
Event|Event|SIMPLE_SEGMENT|11316,11320|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|11316,11320|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|11316,11320|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|11316,11320|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|11322,11331|false|false|false|C0017642|glipizide|glipizide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11322,11331|false|false|false|C0017642|glipizide|glipizide
Event|Event|SIMPLE_SEGMENT|11322,11331|false|false|false|||glipizide
Drug|Organic Chemical|SIMPLE_SEGMENT|11336,11345|false|false|false|C0025598|metformin|metformin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11336,11345|false|false|false|C0025598|metformin|metformin
Event|Event|SIMPLE_SEGMENT|11336,11345|false|false|false|||metformin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11348,11351|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|11348,11351|false|false|false|||HTN
Event|Event|SIMPLE_SEGMENT|11353,11357|false|false|false|||Home
Finding|Idea or Concept|SIMPLE_SEGMENT|11353,11357|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|11353,11357|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|11353,11357|false|false|false|C1553498|home health encounter|Home
Drug|Organic Chemical|SIMPLE_SEGMENT|11363,11373|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11363,11373|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|SIMPLE_SEGMENT|11363,11373|false|false|false|||metoprolol
Event|Event|SIMPLE_SEGMENT|11374,11384|false|false|false|||uptitrated
Event|Event|SIMPLE_SEGMENT|11387,11391|false|false|false|||Home
Finding|Idea or Concept|SIMPLE_SEGMENT|11387,11391|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|11387,11391|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|11387,11391|false|false|false|C1553498|home health encounter|Home
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11397,11407|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11397,11407|false|false|false|C0065374|lisinopril|lisinopril
Event|Event|SIMPLE_SEGMENT|11397,11407|false|false|false|||lisinopril
Event|Event|SIMPLE_SEGMENT|11409,11418|false|false|false|||decreased
Event|Event|SIMPLE_SEGMENT|11421,11425|false|false|false|||Home
Finding|Idea or Concept|SIMPLE_SEGMENT|11421,11425|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|11421,11425|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|11421,11425|false|false|false|C1553498|home health encounter|Home
Drug|Organic Chemical|SIMPLE_SEGMENT|11431,11436|false|false|false|C0590690|Imdur|imdur
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11431,11436|false|false|false|C0590690|Imdur|imdur
Event|Event|SIMPLE_SEGMENT|11431,11436|false|false|false|||imdur
Event|Event|SIMPLE_SEGMENT|11437,11449|false|false|false|||discontinued
Event|Event|SIMPLE_SEGMENT|11453,11456|false|false|false|||HLD
Event|Event|SIMPLE_SEGMENT|11471,11475|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|11471,11475|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|11471,11475|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|11471,11475|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|11481,11492|false|false|false|C0074554|simvastatin|simvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11481,11492|false|false|false|C0074554|simvastatin|simvastatin
Event|Event|SIMPLE_SEGMENT|11481,11492|false|false|false|||simvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|11496,11508|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11496,11508|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|SIMPLE_SEGMENT|11496,11508|false|false|false|||atorvastatin
Finding|Idea or Concept|SIMPLE_SEGMENT|11510,11522|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Event|Event|SIMPLE_SEGMENT|11554,11563|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|11554,11563|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|11554,11563|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|11554,11563|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|11554,11563|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11564,11570|false|false|false|C0944911||weight
Event|Event|SIMPLE_SEGMENT|11564,11570|false|false|false|||weight
Finding|Finding|SIMPLE_SEGMENT|11564,11570|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|11564,11570|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|11564,11570|false|false|false|C1305866|Weighing patient|weight
Finding|Body Substance|SIMPLE_SEGMENT|11582,11589|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|11582,11589|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|11582,11589|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|11595,11602|false|false|false|||require
Event|Event|SIMPLE_SEGMENT|11611,11619|false|false|false|||followup
Procedure|Health Care Activity|SIMPLE_SEGMENT|11611,11619|false|false|false|C1522577|follow-up|followup
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11626,11635|false|false|false|C0018965|Hematuria|hematuria
Event|Event|SIMPLE_SEGMENT|11626,11635|false|false|false|||hematuria
Event|Event|SIMPLE_SEGMENT|11644,11653|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|11644,11653|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Body Substance|SIMPLE_SEGMENT|11656,11661|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Functional Concept|SIMPLE_SEGMENT|11656,11661|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Intellectual Product|SIMPLE_SEGMENT|11656,11661|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Finding|SIMPLE_SEGMENT|11656,11670|false|false|false|C0587953|Urine cytology (finding)|Urine cytology
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11656,11670|false|false|false|C2979983|Urine cytology|Urine cytology
Event|Event|SIMPLE_SEGMENT|11662,11670|false|false|false|||cytology
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11662,11670|false|false|false|C0010818;C1305671|Cytological Techniques;Cytology--Technique|cytology
Event|Event|SIMPLE_SEGMENT|11671,11679|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|11671,11679|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|11671,11679|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|11671,11679|false|false|false|C5237010|Expression Negative|negative
Finding|Body Substance|SIMPLE_SEGMENT|11683,11690|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|11683,11690|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|11683,11690|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|11696,11700|false|false|false|||need
Event|Event|SIMPLE_SEGMENT|11707,11714|false|false|false|||treated
Event|Event|SIMPLE_SEGMENT|11719,11726|false|false|false|||hpylori
Event|Event|SIMPLE_SEGMENT|11748,11754|false|false|false|||course
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11761,11771|false|false|false|C0042313|vancomycin|Vancomycin
Drug|Antibiotic|SIMPLE_SEGMENT|11761,11771|false|false|false|C0042313|vancomycin|Vancomycin
Event|Event|SIMPLE_SEGMENT|11761,11771|false|false|false|||Vancomycin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11761,11771|false|false|false|C0489941|Vancomycin measurement|Vancomycin
Finding|Finding|SIMPLE_SEGMENT|11776,11782|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Finding|Intellectual Product|SIMPLE_SEGMENT|11776,11782|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Event|Event|SIMPLE_SEGMENT|11783,11788|false|false|false|||CDiff
Event|Event|SIMPLE_SEGMENT|11798,11803|false|false|false|||check
Drug|Inorganic Chemical|SIMPLE_SEGMENT|11804,11816|false|false|false|C0013832;C3536863|Electrolyte [EPC];Electrolytes|electrolytes
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11804,11816|false|false|false|C0013832;C3536863|Electrolyte [EPC];Electrolytes|electrolytes
Event|Event|SIMPLE_SEGMENT|11804,11816|false|false|false|||electrolytes
Drug|Organic Chemical|SIMPLE_SEGMENT|11835,11843|false|false|false|C0699129|Coumadin|Coumadin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11835,11843|false|false|false|C0699129|Coumadin|Coumadin
Event|Event|SIMPLE_SEGMENT|11835,11843|false|false|false|||Coumadin
Event|Event|SIMPLE_SEGMENT|11844,11853|false|false|false|||initiated
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|11860,11866|false|false|false|C0018792|Heart Atrium|atrial
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11860,11879|false|false|false|C2926591||atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11860,11879|false|false|false|C0004238|Atrial Fibrillation|atrial fibrillation
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|11860,11879|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|11867,11879|false|false|false|C0232197|Fibrillation|fibrillation
Event|Event|SIMPLE_SEGMENT|11867,11879|false|false|false|||fibrillation
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11881,11884|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Enzyme|SIMPLE_SEGMENT|11881,11884|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Organic Chemical|SIMPLE_SEGMENT|11881,11884|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11881,11884|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Event|Event|SIMPLE_SEGMENT|11881,11884|false|false|false|||ASA
Finding|Gene or Genome|SIMPLE_SEGMENT|11881,11884|false|false|false|C1412553|ARSA gene|ASA
Event|Event|SIMPLE_SEGMENT|11885,11894|false|false|false|||decreased
Event|Event|SIMPLE_SEGMENT|11925,11932|false|false|false|||Started
Drug|Organic Chemical|SIMPLE_SEGMENT|11936,11942|false|false|false|C0633084|Plavix|Plavix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11936,11942|false|false|false|C0633084|Plavix|Plavix
Event|Event|SIMPLE_SEGMENT|11936,11942|false|false|false|||Plavix
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11956,11971|false|false|false|C2348535|Stenting|stent placement
Event|Event|SIMPLE_SEGMENT|11962,11971|false|false|false|||placement
Procedure|Health Care Activity|SIMPLE_SEGMENT|11962,11971|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11962,11971|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Drug|Organic Chemical|SIMPLE_SEGMENT|11973,11985|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11973,11985|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|SIMPLE_SEGMENT|11973,11985|false|false|false|||atorvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|12002,12013|false|false|false|C0074554|simvastatin|simvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12002,12013|false|false|false|C0074554|simvastatin|simvastatin
Event|Event|SIMPLE_SEGMENT|12002,12013|false|false|false|||simvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|12020,12025|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12020,12025|false|false|false|C0699992|Lasix|Lasix
Event|Event|SIMPLE_SEGMENT|12043,12047|false|false|false|||Home
Finding|Idea or Concept|SIMPLE_SEGMENT|12043,12047|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|12043,12047|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|12043,12047|false|false|false|C1553498|home health encounter|Home
Drug|Organic Chemical|SIMPLE_SEGMENT|12048,12058|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12048,12058|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|SIMPLE_SEGMENT|12048,12058|false|false|false|||metoprolol
Event|Event|SIMPLE_SEGMENT|12063,12072|false|false|false|||increased
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12107,12117|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12107,12117|false|false|false|C0065374|lisinopril|lisinopril
Event|Event|SIMPLE_SEGMENT|12107,12117|false|false|false|||lisinopril
Event|Event|SIMPLE_SEGMENT|12118,12127|false|false|false|||decreased
Finding|Idea or Concept|SIMPLE_SEGMENT|12151,12155|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|12151,12155|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|12151,12155|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|12156,12161|false|false|false|C0590690|Imdur|imdur
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12156,12161|false|false|false|C0590690|Imdur|imdur
Event|Event|SIMPLE_SEGMENT|12156,12161|false|false|false|||imdur
Event|Event|SIMPLE_SEGMENT|12167,12179|false|false|false|||discontinued
Finding|Body Substance|SIMPLE_SEGMENT|12182,12189|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|12182,12189|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|12182,12189|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|12195,12199|false|false|false|||need
Event|Event|SIMPLE_SEGMENT|12203,12211|false|false|false|||continue
Finding|Idea or Concept|SIMPLE_SEGMENT|12217,12220|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|12217,12220|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|12221,12227|false|false|false|||course
Finding|Idea or Concept|SIMPLE_SEGMENT|12240,12243|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|12240,12243|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Idea or Concept|SIMPLE_SEGMENT|12259,12262|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|12259,12262|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12277,12286|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|12277,12286|false|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|12277,12286|false|false|false|C3714514|Infection|infection
Finding|Body Substance|SIMPLE_SEGMENT|12289,12296|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|12289,12296|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|12289,12296|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|12297,12307|false|false|false|||instructed
Event|Event|SIMPLE_SEGMENT|12315,12319|false|false|false|||take
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12324,12330|true|false|false|C0003211;C0358845|Analgesics and non-steroidal anti-inflammatory drugs;Anti-Inflammatory Agents, Non-Steroidal|NSAIDS
Event|Event|SIMPLE_SEGMENT|12324,12330|false|false|false|||NSAIDS
Finding|Gene or Genome|SIMPLE_SEGMENT|12333,12336|false|false|false|C1412999;C4283853|C4A gene;C4A wt Allele|SLP
Event|Event|SIMPLE_SEGMENT|12337,12346|false|false|false|||treatment
Finding|Conceptual Entity|SIMPLE_SEGMENT|12337,12346|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|SIMPLE_SEGMENT|12337,12346|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|SIMPLE_SEGMENT|12337,12346|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12337,12346|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12350,12355|false|false|false|C0034991|Rehabilitation therapy|rehab
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12360,12370|false|false|false|C0031354|Pharyngeal structure|pharyngeal
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12371,12394|false|false|false|C0452260|Muscular strength development exercise|strengthening exercises
Event|Event|SIMPLE_SEGMENT|12385,12394|false|false|false|||exercises
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|12385,12394|false|false|false|C0015259|Exercise|exercises
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12385,12394|false|false|false|C0452240|Physical therapy exercises|exercises
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12397,12408|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12397,12408|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|12397,12408|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|12397,12408|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|12397,12421|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|SIMPLE_SEGMENT|12412,12421|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|12412,12421|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12440,12450|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|12440,12450|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|12440,12455|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|SIMPLE_SEGMENT|12451,12455|false|false|false|||list
Finding|Intellectual Product|SIMPLE_SEGMENT|12451,12455|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|SIMPLE_SEGMENT|12459,12467|false|false|false|||accurate
Drug|Organic Chemical|SIMPLE_SEGMENT|12472,12480|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12472,12480|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|12472,12480|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|SIMPLE_SEGMENT|12472,12480|false|false|false|||complete
Finding|Functional Concept|SIMPLE_SEGMENT|12472,12480|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|12472,12480|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|SIMPLE_SEGMENT|12485,12495|false|false|false|C0060926|gabapentin|Gabapentin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12485,12495|false|false|false|C0060926|gabapentin|Gabapentin
Event|Event|SIMPLE_SEGMENT|12506,12509|false|false|false|||TID
Drug|Organic Chemical|SIMPLE_SEGMENT|12514,12522|false|false|false|C0027396|naproxen|Naproxen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12514,12522|false|false|false|C0027396|naproxen|Naproxen
Drug|Organic Chemical|SIMPLE_SEGMENT|12543,12552|false|false|false|C0025598|metformin|MetFORMIN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12543,12552|false|false|false|C0025598|metformin|MetFORMIN
Drug|Organic Chemical|SIMPLE_SEGMENT|12554,12564|false|false|false|C0591573|Glucophage|Glucophage
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12554,12564|false|false|false|C0591573|Glucophage|Glucophage
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|12576,12579|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12576,12579|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12576,12579|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|12576,12579|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|12576,12579|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|12584,12594|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12584,12594|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|12584,12604|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12584,12604|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|12595,12604|false|false|false|C0038617;C0220918|Succinates;succinate|Succinate
Event|Event|SIMPLE_SEGMENT|12595,12604|false|false|false|||Succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|12627,12636|false|false|false|C0017642|glipizide|GlipiZIDE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12627,12636|false|false|false|C0017642|glipizide|GlipiZIDE
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|12647,12650|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12647,12650|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12647,12650|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|12647,12650|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|12647,12650|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|12655,12666|false|false|false|C0074554|simvastatin|Simvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12655,12666|false|false|false|C0074554|simvastatin|Simvastatin
Event|Event|SIMPLE_SEGMENT|12676,12679|false|false|false|||QPM
Drug|Organic Chemical|SIMPLE_SEGMENT|12684,12694|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12684,12694|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|SIMPLE_SEGMENT|12684,12706|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12684,12706|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Event|Event|SIMPLE_SEGMENT|12695,12706|false|false|false|||Mononitrate
Finding|Finding|SIMPLE_SEGMENT|12708,12716|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|12708,12716|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|SIMPLE_SEGMENT|12717,12724|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|12717,12724|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|12717,12724|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12717,12724|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12745,12755|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12745,12755|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Organic Chemical|SIMPLE_SEGMENT|12775,12782|false|false|false|C0012265|digoxin|Digoxin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12775,12782|false|false|false|C0012265|digoxin|Digoxin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12775,12782|false|false|false|C0337449|Digoxin measurement|Digoxin
Drug|Organic Chemical|SIMPLE_SEGMENT|12806,12813|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12806,12813|false|false|false|C0004057|aspirin|Aspirin
Event|Event|SIMPLE_SEGMENT|12834,12843|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|12834,12843|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|12834,12843|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|12834,12843|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|12834,12843|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|12834,12855|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12844,12855|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12844,12855|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|12844,12855|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|12844,12855|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|12860,12867|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12860,12867|false|false|false|C0004057|aspirin|Aspirin
Event|Event|SIMPLE_SEGMENT|12860,12867|false|false|false|||Aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|12860,12870|false|false|false|C5874014|Aspirin EC|Aspirin EC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12860,12870|false|false|false|C5874014|Aspirin EC|Aspirin EC
Drug|Organic Chemical|SIMPLE_SEGMENT|12890,12897|false|false|false|C0012265|digoxin|Digoxin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12890,12897|false|false|false|C0012265|digoxin|Digoxin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12890,12897|false|false|false|C0337449|Digoxin measurement|Digoxin
Drug|Organic Chemical|SIMPLE_SEGMENT|12920,12930|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12920,12930|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|12920,12940|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12920,12940|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|12931,12940|false|false|false|C0038617;C0220918|Succinates;succinate|Succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|12963,12975|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12963,12975|false|false|false|C0286651|atorvastatin|Atorvastatin
Event|Event|SIMPLE_SEGMENT|12985,12988|false|false|false|||QPM
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|12993,13001|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|SIMPLE_SEGMENT|12993,13001|false|false|false|C0043031|warfarin|Warfarin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12993,13001|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|SIMPLE_SEGMENT|13022,13031|false|false|false|C0017642|glipizide|GlipiZIDE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13022,13031|false|false|false|C0017642|glipizide|GlipiZIDE
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|13042,13045|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13042,13045|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|13042,13045|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|13042,13045|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|13042,13045|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|13050,13061|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13050,13061|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Organic Chemical|SIMPLE_SEGMENT|13081,13091|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13081,13091|false|false|false|C0028978|omeprazole|Omeprazole
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|13101,13104|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13101,13104|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|13101,13104|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|13101,13104|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|13101,13104|false|false|false|C1332410|BID gene|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13109,13119|false|false|false|C0042313|vancomycin|Vancomycin
Drug|Antibiotic|SIMPLE_SEGMENT|13109,13119|false|false|false|C0042313|vancomycin|Vancomycin
Event|Event|SIMPLE_SEGMENT|13109,13119|false|false|false|||Vancomycin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|13109,13119|false|false|false|C0489941|Vancomycin measurement|Vancomycin
Drug|Clinical Drug|SIMPLE_SEGMENT|13109,13124|false|false|false|C0360373||Vancomycin Oral
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|13120,13124|false|false|false|C0226896|Oral cavity|Oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13120,13124|false|false|false|C1272919|Oral Dosage Form|Oral
Finding|Finding|SIMPLE_SEGMENT|13120,13124|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Finding|Functional Concept|SIMPLE_SEGMENT|13120,13124|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13120,13131|false|false|false|C1273619|Oral Liquid Product|Oral Liquid
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|13125,13131|false|false|false|C0302908;C1697794|Liquid Dosage Form;Liquid substance|Liquid
Drug|Substance|SIMPLE_SEGMENT|13125,13131|false|false|false|C0302908;C1697794|Liquid Dosage Form;Liquid substance|Liquid
Event|Event|SIMPLE_SEGMENT|13125,13131|false|false|false|||Liquid
Finding|Finding|SIMPLE_SEGMENT|13125,13131|false|false|false|C1304698|Liquid (finding)|Liquid
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|13125,13131|false|false|false|C0301571|Liquid diet|Liquid
Drug|Organic Chemical|SIMPLE_SEGMENT|13151,13160|false|false|false|C0025598|metformin|MetFORMIN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13151,13160|false|false|false|C0025598|metformin|MetFORMIN
Drug|Organic Chemical|SIMPLE_SEGMENT|13162,13172|false|false|false|C0591573|Glucophage|Glucophage
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13162,13172|false|false|false|C0591573|Glucophage|Glucophage
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|13184,13187|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13184,13187|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|13184,13187|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|13184,13187|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|13184,13187|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|13193,13203|false|false|false|C0060926|gabapentin|Gabapentin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13193,13203|false|false|false|C0060926|gabapentin|Gabapentin
Event|Event|SIMPLE_SEGMENT|13214,13217|false|false|false|||TID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|13223,13233|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13223,13233|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Organic Chemical|SIMPLE_SEGMENT|13255,13265|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13255,13265|false|false|false|C0016860|furosemide|Furosemide
Event|Event|SIMPLE_SEGMENT|13285,13294|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|13285,13294|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|13285,13294|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|13285,13294|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|13285,13294|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13285,13306|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|13285,13306|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13295,13306|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|13295,13306|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|13295,13306|false|false|false|C0184758|Patient disposition|Disposition
Finding|Finding|SIMPLE_SEGMENT|13308,13316|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|13308,13316|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Procedure|Health Care Activity|SIMPLE_SEGMENT|13308,13321|false|false|false|C0023977|long-term care|Extended Care
Event|Activity|SIMPLE_SEGMENT|13317,13321|false|false|false|C1947933|care activity|Care
Event|Event|SIMPLE_SEGMENT|13317,13321|false|false|false|||Care
Finding|Finding|SIMPLE_SEGMENT|13317,13321|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|SIMPLE_SEGMENT|13317,13321|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Event|Event|SIMPLE_SEGMENT|13324,13332|false|false|false|||Facility
Finding|Intellectual Product|SIMPLE_SEGMENT|13324,13332|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|SIMPLE_SEGMENT|13340,13349|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|13340,13349|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|13340,13349|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|13340,13349|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|13340,13349|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|13340,13359|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13350,13359|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|13350,13359|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|13350,13359|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|13350,13359|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|13350,13359|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13361,13367|false|false|false|C4255010||NSTEMI
Event|Event|SIMPLE_SEGMENT|13361,13367|false|false|false|||NSTEMI
Finding|Finding|SIMPLE_SEGMENT|13361,13367|false|false|false|C3537184||NSTEMI
Finding|Finding|SIMPLE_SEGMENT|13377,13383|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|13377,13383|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Finding|SIMPLE_SEGMENT|13384,13389|false|true|false|C0205430;C3160715|Mixed (Normal and Tumor);Mixed (qualifier value)|mixed
Finding|Functional Concept|SIMPLE_SEGMENT|13384,13389|false|true|false|C0205430;C3160715|Mixed (Normal and Tumor);Mixed (qualifier value)|mixed
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13416,13425|false|false|false|C0018965|Hematuria|Hematuria
Event|Event|SIMPLE_SEGMENT|13416,13425|false|false|false|||Hematuria
Finding|Finding|SIMPLE_SEGMENT|13426,13433|false|false|false|C0013404;C2024878|Dyspnea|Dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|13426,13433|false|false|false|C0013404;C2024878|Dyspnea|Dyspnea
Finding|Gene or Genome|SIMPLE_SEGMENT|13437,13440|false|false|false|C0812246;C1710304|TNF gene;TNF wt Allele|dif
Event|Event|SIMPLE_SEGMENT|13442,13448|false|false|false|||severe
Finding|Finding|SIMPLE_SEGMENT|13442,13448|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|13442,13448|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13449,13453|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|SIMPLE_SEGMENT|13449,13453|false|false|false|||GERD
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|13454,13462|false|false|false|C0011206|Delirium|Delirium
Event|Event|SIMPLE_SEGMENT|13454,13462|false|false|false|||Delirium
Event|Event|SIMPLE_SEGMENT|13466,13475|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|13466,13475|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|13466,13475|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|13466,13475|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|13466,13475|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13476,13485|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13476,13485|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|13476,13485|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|13476,13485|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|13487,13493|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13487,13500|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|13487,13500|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13494,13500|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|13494,13500|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|13502,13507|false|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|13502,13507|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|13512,13520|false|false|false|||coherent
Finding|Finding|SIMPLE_SEGMENT|13512,13520|false|false|false|C4068804|Coherent|coherent
Event|Event|SIMPLE_SEGMENT|13522,13527|false|false|false|||Level
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13522,13544|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|13522,13544|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|SIMPLE_SEGMENT|13531,13544|false|false|false|||Consciousness
Finding|Finding|SIMPLE_SEGMENT|13531,13544|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|13531,13544|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13546,13551|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|13546,13551|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13546,13551|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|13546,13551|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|13546,13551|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|13546,13551|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|13546,13551|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|13556,13567|false|false|false|||interactive
Finding|Functional Concept|SIMPLE_SEGMENT|13556,13567|false|false|false|C1704675|Interaction|interactive
Event|Event|SIMPLE_SEGMENT|13571,13580|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|13571,13580|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|13571,13580|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|13571,13580|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|13571,13580|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13571,13593|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|13571,13593|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|13571,13593|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13581,13593|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|13581,13593|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|13581,13593|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Finding|Gene or Genome|SIMPLE_SEGMENT|13595,13599|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|SIMPLE_SEGMENT|13619,13627|false|false|false|||admitted
Anatomy|Body Location or Region|SIMPLE_SEGMENT|13665,13670|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|13665,13670|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13672,13676|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|13672,13676|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|13672,13676|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|13672,13676|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|13686,13691|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|13686,13691|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|13686,13691|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13686,13698|false|false|false|C0027051|Myocardial Infarction|heart attack
Event|Event|SIMPLE_SEGMENT|13692,13698|false|false|false|||attack
Finding|Finding|SIMPLE_SEGMENT|13692,13698|false|false|false|C1261512;C1304680|Attack (finding);Attack behavior|attack
Finding|Social Behavior|SIMPLE_SEGMENT|13692,13698|false|false|false|C1261512;C1304680|Attack (finding);Attack behavior|attack
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|13707,13711|false|false|false|C0007430|Catheterization|cath
Finding|Gene or Genome|SIMPLE_SEGMENT|13712,13715|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|lab
Finding|Intellectual Product|SIMPLE_SEGMENT|13712,13715|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|lab
Event|Event|SIMPLE_SEGMENT|13725,13730|false|false|false|||found
Event|Event|SIMPLE_SEGMENT|13740,13748|false|false|false|||blockage
Finding|Finding|SIMPLE_SEGMENT|13740,13748|false|false|false|C1706968;C1879887;C2237319|Blockage (obstruction - finding);Partial Blockage within Medical Device|blockage
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|13757,13765|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Anatomy|Body System|SIMPLE_SEGMENT|13757,13765|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Procedure|Health Care Activity|SIMPLE_SEGMENT|13757,13765|false|false|false|C0397581|Procedure on artery|arteries
Event|Event|SIMPLE_SEGMENT|13773,13778|false|false|false|||stent
Event|Event|SIMPLE_SEGMENT|13783,13789|false|false|false|||placed
Event|Event|SIMPLE_SEGMENT|13800,13807|false|false|false|||managed
Finding|Finding|SIMPLE_SEGMENT|13813,13816|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|SIMPLE_SEGMENT|13813,13816|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Finding|SIMPLE_SEGMENT|13813,13831|false|false|false|C0020649|Hypotension|low blood pressure
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13817,13822|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|13817,13822|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|13817,13822|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|SIMPLE_SEGMENT|13817,13831|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Finding|Organism Function|SIMPLE_SEGMENT|13817,13831|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Procedure|Health Care Activity|SIMPLE_SEGMENT|13817,13831|false|false|false|C0005824|Blood pressure determination|blood pressure
Event|Event|SIMPLE_SEGMENT|13823,13831|false|false|false|||pressure
Finding|Finding|SIMPLE_SEGMENT|13823,13831|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|13823,13831|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|13823,13831|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|13823,13831|false|false|false|C0033095||pressure
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13833,13843|false|false|false|C0009450|Communicable Diseases|infectious
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13833,13852|false|false|false|C0013369|Dysentery|infectious diarrhea
Event|Event|SIMPLE_SEGMENT|13844,13852|false|false|false|||diarrhea
Finding|Finding|SIMPLE_SEGMENT|13844,13852|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|13844,13852|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|13858,13864|false|false|false|C1368081;C3263723;C3714660|Physical trauma;Trauma;Traumatic injury|trauma
Event|Event|SIMPLE_SEGMENT|13858,13864|false|false|false|||trauma
Procedure|Health Care Activity|SIMPLE_SEGMENT|13858,13864|false|false|false|C0548346|Trauma assessment and care|trauma
Event|Event|SIMPLE_SEGMENT|13877,13886|false|false|false|||placement
Procedure|Health Care Activity|SIMPLE_SEGMENT|13877,13886|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|13877,13886|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Event|Event|SIMPLE_SEGMENT|13892,13901|false|false|false|||responded
Finding|Finding|SIMPLE_SEGMENT|13902,13906|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|13917,13925|false|false|false|||continue
Event|Event|SIMPLE_SEGMENT|13926,13932|false|false|false|||taking
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13938,13949|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13938,13949|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|13938,13949|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|13938,13949|false|false|false|C4284232|Medications|medications
Event|Event|SIMPLE_SEGMENT|13953,13963|false|false|false|||prescribed
Event|Event|SIMPLE_SEGMENT|13981,13988|false|false|false|||started
Drug|Organic Chemical|SIMPLE_SEGMENT|13992,14000|false|false|false|C0699129|Coumadin|coumadin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13992,14000|false|false|false|C0699129|Coumadin|coumadin
Event|Event|SIMPLE_SEGMENT|13992,14000|false|false|false|||coumadin
Event|Event|SIMPLE_SEGMENT|14017,14021|false|false|false|||take
Event|Event|SIMPLE_SEGMENT|14026,14039|false|false|false|||non-steroidal
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14041,14057|false|false|false|C0003209|Anti-Inflammatory Agents|antiinflammatory
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14058,14063|false|false|false|C0013227|Pharmaceutical Preparations|drugs
Event|Event|SIMPLE_SEGMENT|14058,14063|false|false|false|||drugs
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|14058,14063|false|false|false|C3687832|Drugs - dental services|drugs
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14065,14071|false|false|false|C0003211;C0358845|Analgesics and non-steroidal anti-inflammatory drugs;Anti-Inflammatory Agents, Non-Steroidal|NSAIDS
Event|Event|SIMPLE_SEGMENT|14065,14071|false|false|false|||NSAIDS
Drug|Organic Chemical|SIMPLE_SEGMENT|14081,14090|false|false|false|C0020740|ibuprofen|ibuprofen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14081,14090|false|false|false|C0020740|ibuprofen|ibuprofen
Event|Event|SIMPLE_SEGMENT|14081,14090|false|false|false|||ibuprofen
Drug|Organic Chemical|SIMPLE_SEGMENT|14092,14097|false|false|false|C0593507|Advil|advil
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14092,14097|false|false|false|C0593507|Advil|advil
Event|Event|SIMPLE_SEGMENT|14092,14097|false|false|false|||advil
Finding|Gene or Genome|SIMPLE_SEGMENT|14092,14097|false|false|false|C1422473|AVIL gene|advil
Drug|Organic Chemical|SIMPLE_SEGMENT|14100,14106|false|false|false|C0699203|Motrin|motrin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14100,14106|false|false|false|C0699203|Motrin|motrin
Event|Event|SIMPLE_SEGMENT|14100,14106|false|false|false|||motrin
Drug|Organic Chemical|SIMPLE_SEGMENT|14108,14113|false|false|false|C0718343|Aleve|aleve
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14108,14113|false|false|false|C0718343|Aleve|aleve
Event|Event|SIMPLE_SEGMENT|14108,14113|false|false|false|||aleve
Drug|Organic Chemical|SIMPLE_SEGMENT|14115,14123|false|false|false|C0027396|naproxen|naproxen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14115,14123|false|false|false|C0027396|naproxen|naproxen
Event|Event|SIMPLE_SEGMENT|14115,14123|false|false|false|||naproxen
Event|Event|SIMPLE_SEGMENT|14138,14144|false|false|false|||follow
Anatomy|Body System|SIMPLE_SEGMENT|14159,14169|false|false|false|C0007226|Cardiovascular system|cardiology
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|14174,14177|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|14174,14177|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|14174,14177|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|14174,14177|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|14174,14177|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|14174,14177|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|14174,14177|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|14174,14177|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|14174,14177|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|14174,14177|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|14174,14177|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Activity|SIMPLE_SEGMENT|14178,14190|false|false|false|C0003629|Appointments|appointments
Event|Event|SIMPLE_SEGMENT|14178,14190|false|false|false|||appointments
Event|Event|SIMPLE_SEGMENT|14194,14203|false|false|false|||scheduled
Event|Event|SIMPLE_SEGMENT|14214,14222|false|false|false|||pleasure
Finding|Intellectual Product|SIMPLE_SEGMENT|14214,14222|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|SIMPLE_SEGMENT|14214,14222|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|SIMPLE_SEGMENT|14230,14234|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|14230,14234|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|14230,14234|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|14230,14234|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|14230,14237|false|false|false|C1555558|care of - AddressPartType|care of
Event|Activity|SIMPLE_SEGMENT|14252,14256|false|false|false|C1947933|care activity|Care
Finding|Finding|SIMPLE_SEGMENT|14252,14256|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|SIMPLE_SEGMENT|14252,14256|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14252,14261|false|false|false|C4321316||Care Team
Finding|Finding|SIMPLE_SEGMENT|14252,14261|false|false|false|C4321315|Care team|Care Team
Procedure|Health Care Activity|SIMPLE_SEGMENT|14264,14272|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|14273,14285|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|14273,14285|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|14273,14285|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

