 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|33,37
No|38,40
:|40,41
_|44,45
_|45,46
_|46,47
<EOL>|47,48
<EOL>|49,50
Admission|50,59
Date|60,64
:|64,65
_|67,68
_|68,69
_|69,70
Discharge|84,93
Date|94,98
:|98,99
_|102,103
_|103,104
_|104,105
<EOL>|105,106
<EOL>|107,108
Date|108,112
of|113,115
Birth|116,121
:|121,122
_|124,125
_|125,126
_|126,127
Sex|140,143
:|143,144
F|147,148
<EOL>|148,149
<EOL>|150,151
Service|151,158
:|158,159
MEDICINE|160,168
<EOL>|168,169
<EOL>|170,171
Allergies|171,180
:|180,181
<EOL>|182,183
Percocet|183,191
/|192,193
Vicodin|194,201
<EOL>|201,202
<EOL>|203,204
Attending|204,213
:|213,214
_|215,216
_|216,217
_|217,218
.|218,219
<EOL>|219,220
<EOL>|221,222
Chief|222,227
Complaint|228,237
:|237,238
<EOL>|238,239
Abdominal|239,248
pain|249,253
<EOL>|253,254
<EOL>|255,256
Major|256,261
Surgical|262,270
or|271,273
Invasive|274,282
Procedure|283,292
:|292,293
<EOL>|293,294
_|294,295
_|295,296
_|296,297
Paracentesis|298,310
<EOL>|310,311
<EOL>|311,312
<EOL>|313,314
History|314,321
of|322,324
Present|325,332
Illness|333,340
:|340,341
<EOL>|341,342
_|342,343
_|343,344
_|344,345
w|346,347
/|347,348
HIV|349,352
on|353,355
HAART|356,361
,|361,362
COPD|363,367
on|368,370
3L|371,373
home|374,378
O2|379,381
(|382,383
though|383,389
sat|390,393
'|393,394
ing|394,397
fine|398,402
on|403,405
<EOL>|406,407
RA|407,409
on|410,412
admission|413,422
)|422,423
,|423,424
HCV|425,428
cirrhosis|429,438
c|439,440
/|440,441
b|441,442
ascites|443,450
requiring|451,460
biweekly|461,469
<EOL>|470,471
therapeutic|471,482
paracenteses|483,495
,|495,496
hepatic|497,504
encephalopathy|505,519
;|519,520
not|521,524
on|525,527
<EOL>|528,529
transplant|529,539
list|540,544
_|545,546
_|546,547
_|547,548
comorbidities|549,562
)|562,563
p|564,565
/|565,566
w|566,567
worsening|568,577
girth|578,583
and|584,587
abd|588,591
<EOL>|592,593
pain|593,597
.|597,598
She|599,602
'd|602,604
been|605,609
having|610,616
pain|617,621
from|622,626
her|627,630
ascites|631,638
,|638,639
and|640,643
felt|644,648
overdue|649,656
<EOL>|657,658
for|658,661
a|662,663
paracentesis|664,676
.|676,677
She|678,681
last|682,686
had|687,690
paracentesis|691,703
on|704,706
the|707,710
_|711,712
_|712,713
_|713,714
.|714,715
<EOL>|716,717
She|717,720
reported|721,729
that|730,734
she|735,738
began|739,744
feeling|745,752
worsening|753,762
abdominal|763,772
pain|773,777
<EOL>|778,779
(|779,780
constant|780,788
,|788,789
epigastric|790,800
and|801,804
radiates|805,813
to|814,816
back|817,821
,|821,822
not|823,826
a|827,828
/|828,829
w|829,830
food|831,835
)|835,836
on|837,839
<EOL>|840,841
_|841,842
_|842,843
_|843,844
,|844,845
which|846,851
increased|852,861
in|862,864
severity|865,873
throughout|874,884
the|885,888
course|889,895
of|896,898
the|899,902
<EOL>|903,904
day|904,907
.|907,908
She|909,912
was|913,916
brought|917,924
to|925,927
the|928,931
ED|932,934
by|935,937
her|938,941
son|942,945
because|946,953
of|954,956
this|957,961
pain|962,966
.|966,967
<EOL>|968,969
She|969,972
had|973,976
no|977,979
confusion|980,989
and|990,993
was|994,997
alert|998,1003
and|1004,1007
oriented|1008,1016
x3|1017,1019
.|1019,1020
The|1021,1024
patient|1025,1032
<EOL>|1033,1034
also|1034,1038
reported|1039,1047
she|1048,1051
recently|1052,1060
ran|1061,1064
out|1065,1068
of|1069,1071
most|1072,1076
of|1077,1079
her|1080,1083
home|1084,1088
<EOL>|1089,1090
medications|1090,1101
.|1101,1102
She|1103,1106
denied|1107,1113
any|1114,1117
fever|1118,1123
,|1123,1124
chills|1125,1131
,|1131,1132
shortness|1133,1142
of|1143,1145
breath|1146,1152
,|1152,1153
<EOL>|1154,1155
cough|1155,1160
,|1160,1161
dysuria|1162,1169
.|1169,1170
She|1171,1174
reported|1175,1183
loose|1184,1189
stool|1190,1195
a|1196,1197
bit|1198,1201
more|1202,1206
than|1207,1211
usual|1212,1217
,|1217,1218
<EOL>|1219,1220
but|1220,1223
attributed|1224,1234
it|1235,1237
to|1238,1240
lactulose|1241,1250
use|1251,1254
.|1254,1255
In|1256,1258
the|1259,1262
ED|1263,1265
,|1265,1266
vitals|1267,1273
were|1274,1278
:|1278,1279
99.4|1280,1284
<EOL>|1285,1286
105|1286,1289
106|1290,1293
/|1293,1294
57|1294,1296
18|1297,1299
96|1300,1302
%|1302,1303
ra|1304,1306
.|1306,1307
Labs|1308,1312
were|1313,1317
significant|1318,1329
for|1330,1333
Na|1334,1336
127|1337,1340
K|1341,1342
5.3|1343,1346
<EOL>|1347,1348
lactate|1348,1355
2.1|1356,1359
INR|1360,1363
1.7|1364,1367
.|1367,1368
ALT|1369,1372
135|1373,1376
AST|1377,1380
244|1381,1384
AP|1385,1387
123|1388,1391
.|1391,1392
no|1393,1395
leukocytosis|1396,1408
.|1408,1409
<EOL>|1410,1411
Ascitic|1411,1418
fluid|1419,1424
showed|1425,1431
220|1432,1435
WBC|1436,1439
.|1439,1440
She|1441,1444
was|1445,1448
given|1449,1454
Morphine|1455,1463
Sulfate|1464,1471
5|1472,1473
<EOL>|1474,1475
mg|1475,1477
IV|1478,1480
ONCE|1481,1485
MR1|1486,1489
,|1489,1490
and|1491,1494
a|1495,1496
GI|1497,1499
cocktail|1500,1508
.|1508,1509
<EOL>|1509,1510
<EOL>|1511,1512
Past|1512,1516
Medical|1517,1524
History|1525,1532
:|1532,1533
<EOL>|1533,1534
-|1534,1535
HCV|1536,1539
Cirrhosis|1540,1549
:|1549,1550
genotype|1551,1559
3a|1560,1562
<EOL>|1564,1565
-|1565,1566
HIV|1567,1570
:|1570,1571
on|1572,1574
HAART|1575,1580
,|1580,1581
_|1582,1583
_|1583,1584
_|1584,1585
CD4|1586,1589
count|1590,1595
173|1596,1599
,|1599,1600
_|1601,1602
_|1602,1603
_|1603,1604
HIV|1605,1608
viral|1609,1614
load|1615,1619
<EOL>|1620,1621
undetectable|1621,1633
<EOL>|1635,1636
-|1636,1637
COPD|1638,1642
:|1642,1643
_|1644,1645
_|1645,1646
_|1646,1647
PFT|1648,1651
showed|1652,1658
FVC|1659,1662
1.95|1663,1667
(|1668,1669
65|1669,1671
%|1671,1672
)|1672,1673
,|1673,1674
FEV1|1675,1679
0.88|1680,1684
(|1685,1686
37|1686,1688
%|1688,1689
)|1689,1690
,|1690,1691
<EOL>|1692,1693
FEFmax|1693,1699
2.00|1700,1704
(|1705,1706
33|1706,1708
%|1708,1709
)|1709,1710
<EOL>|1712,1713
-|1713,1714
Bipolar|1715,1722
Affective|1723,1732
Disorder|1733,1741
<EOL>|1743,1744
-|1744,1745
PTSD|1746,1750
<EOL>|1752,1753
-|1753,1754
Hx|1755,1757
of|1758,1760
cocaine|1761,1768
and|1769,1772
heroin|1773,1779
abuse|1780,1785
<EOL>|1787,1788
-|1788,1789
Hx|1790,1792
of|1793,1795
skin|1796,1800
cancer|1801,1807
per|1808,1811
patient|1812,1819
report|1820,1826
<EOL>|1828,1829
<EOL>|1830,1831
Social|1831,1837
History|1838,1845
:|1845,1846
<EOL>|1846,1847
_|1847,1848
_|1848,1849
_|1849,1850
<EOL>|1850,1851
Family|1851,1857
History|1858,1865
:|1865,1866
<EOL>|1866,1867
She|1867,1870
a|1871,1872
total|1873,1878
of|1879,1881
five|1882,1886
siblings|1887,1895
,|1895,1896
but|1897,1900
she|1901,1904
is|1905,1907
not|1908,1911
talking|1913,1920
to|1921,1923
most|1924,1928
of|1929,1931
<EOL>|1932,1933
them|1933,1937
.|1937,1938
She|1939,1942
only|1943,1947
has|1948,1951
one|1952,1955
brother|1956,1963
that|1964,1968
she|1969,1972
is|1973,1975
in|1976,1978
touch|1979,1984
with|1985,1989
and|1990,1993
<EOL>|1994,1995
lives|1995,2000
in|2001,2003
_|2004,2005
_|2005,2006
_|2006,2007
.|2007,2008
She|2009,2012
is|2013,2015
not|2016,2019
aware|2020,2025
of|2026,2028
any|2029,2032
known|2033,2038
GI|2039,2041
or|2042,2044
liver|2045,2050
<EOL>|2051,2052
disease|2052,2059
in|2060,2062
her|2063,2066
family|2067,2073
.|2073,2074
<EOL>|2076,2077
<EOL>|2078,2079
Physical|2079,2087
Exam|2088,2092
:|2092,2093
<EOL>|2093,2094
ADMISSION|2094,2103
PHYSICAL|2104,2112
EXAM|2113,2117
<EOL>|2117,2118
=|2118,2119
=|2119,2120
=|2120,2121
=|2121,2122
=|2122,2123
=|2123,2124
=|2124,2125
=|2125,2126
=|2126,2127
=|2127,2128
=|2128,2129
=|2129,2130
=|2130,2131
=|2131,2132
=|2132,2133
=|2133,2134
=|2134,2135
=|2135,2136
=|2136,2137
=|2137,2138
=|2138,2139
=|2139,2140
=|2140,2141
<EOL>|2141,2142
Vitals|2142,2148
-|2149,2150
T|2151,2152
97|2153,2155
,|2155,2156
BP|2157,2159
98|2160,2162
/|2162,2163
65|2163,2165
,|2165,2166
HR|2167,2169
103|2170,2173
,|2173,2174
RR|2175,2177
18|2178,2180
,|2180,2181
O2|2182,2184
94RA|2185,2189
,|2189,2190
Glucose|2191,2198
128|2199,2202
.|2202,2203
<EOL>|2205,2206
GENERAL|2206,2213
:|2213,2214
NAD|2215,2218
,|2218,2219
lying|2220,2225
on|2226,2228
her|2229,2232
right|2233,2238
side|2239,2243
.|2243,2244
<EOL>|2244,2245
HEENT|2245,2250
:|2250,2251
AT|2252,2254
/|2254,2255
NC|2255,2257
,|2257,2258
EOMI|2259,2263
,|2263,2264
PERRL|2265,2270
,|2270,2271
anicteric|2272,2281
sclera|2282,2288
,|2288,2289
pink|2290,2294
conjunctiva|2295,2306
,|2306,2307
<EOL>|2308,2309
MMM|2309,2312
,|2312,2313
good|2314,2318
dentition|2319,2328
<EOL>|2330,2331
NECK|2331,2335
:|2335,2336
nontender|2337,2346
supple|2347,2353
neck|2354,2358
,|2358,2359
no|2360,2362
LAD|2363,2366
,|2366,2367
no|2368,2370
JVD|2371,2374
<EOL>|2376,2377
CARDIAC|2377,2384
:|2384,2385
RRR|2386,2389
,|2389,2390
S1|2391,2393
/|2393,2394
S2|2394,2396
,|2396,2397
no|2398,2400
murmurs|2401,2408
,|2408,2409
gallops|2410,2417
,|2417,2418
or|2419,2421
rubs|2422,2426
<EOL>|2428,2429
LUNG|2429,2433
:|2433,2434
CTAB|2435,2439
,|2439,2440
no|2441,2443
wheezes|2444,2451
,|2451,2452
rales|2453,2458
,|2458,2459
rhonchi|2460,2467
,|2467,2468
breathing|2469,2478
comfortably|2479,2490
<EOL>|2491,2492
without|2492,2499
use|2500,2503
of|2504,2506
accessory|2507,2516
muscles|2517,2524
<EOL>|2526,2527
ABDOMEN|2527,2534
:|2534,2535
distended|2536,2545
,|2545,2546
+|2547,2548
fluid|2549,2554
wave|2555,2559
,|2559,2560
not|2561,2564
tense|2565,2570
.|2570,2571
NABS|2572,2576
,|2576,2577
nontender|2578,2587
<EOL>|2589,2590
EXTREMITIES|2590,2601
:|2601,2602
no|2603,2605
cyanosis|2606,2614
,|2614,2615
clubbing|2616,2624
or|2625,2627
edema|2628,2633
,|2633,2634
moving|2635,2641
all|2642,2645
4|2646,2647
<EOL>|2648,2649
extremities|2649,2660
with|2661,2665
purpose|2666,2673
<EOL>|2673,2674
PULSES|2674,2680
:|2680,2681
2|2682,2683
+|2683,2684
DP|2685,2687
pulses|2688,2694
bilaterally|2695,2706
<EOL>|2708,2709
NEURO|2709,2714
:|2714,2715
CN|2716,2718
II|2719,2721
-|2721,2722
XII|2722,2725
intact|2726,2732
,|2732,2733
AAO3|2734,2738
,|2738,2739
no|2740,2742
asterxis|2743,2751
<EOL>|2753,2754
SKIN|2754,2758
:|2758,2759
warm|2760,2764
and|2765,2768
well|2769,2773
perfused|2774,2782
,|2782,2783
no|2784,2786
excoriations|2787,2799
or|2800,2802
lesions|2803,2810
,|2810,2811
no|2812,2814
<EOL>|2815,2816
rashes|2816,2822
<EOL>|2822,2823
<EOL>|2823,2824
DISCHARGE|2824,2833
PHYSICAL|2834,2842
EXAM|2843,2847
<EOL>|2847,2848
=|2848,2849
=|2849,2850
=|2850,2851
=|2851,2852
=|2852,2853
=|2853,2854
=|2854,2855
=|2855,2856
=|2856,2857
=|2857,2858
=|2858,2859
=|2859,2860
=|2860,2861
=|2861,2862
=|2862,2863
=|2863,2864
=|2864,2865
=|2865,2866
=|2866,2867
=|2867,2868
=|2868,2869
=|2869,2870
=|2870,2871
<EOL>|2871,2872
Vitals|2872,2878
-|2879,2880
Tm|2881,2883
98.6|2884,2888
,|2888,2889
Tc|2890,2892
98.2|2893,2897
,|2897,2898
BP|2899,2901
82|2902,2904
-|2904,2905
98|2905,2907
/|2907,2908
42|2908,2910
-|2910,2911
68|2911,2913
,|2913,2914
HR|2915,2917
80|2918,2920
-|2920,2921
95|2921,2923
,|2923,2924
RR|2925,2927
_|2928,2929
_|2929,2930
_|2930,2931
,|2931,2932
<EOL>|2933,2934
O2|2934,2936
91|2937,2939
-|2939,2940
99|2940,2942
%|2942,2943
RA|2944,2946
.|2946,2947
<EOL>|2947,2948
GENERAL|2948,2955
:|2955,2956
NAD|2957,2960
,|2960,2961
lying|2962,2967
on|2968,2970
her|2971,2974
right|2975,2980
side|2981,2985
.|2985,2986
<EOL>|2986,2987
HEENT|2987,2992
:|2992,2993
AT|2994,2996
/|2996,2997
NC|2997,2999
,|2999,3000
EOMI|3001,3005
,|3005,3006
PERRL|3007,3012
,|3012,3013
anicteric|3014,3023
sclera|3024,3030
,|3030,3031
pink|3032,3036
conjunctiva|3037,3048
,|3048,3049
<EOL>|3050,3051
MMM|3051,3054
,|3054,3055
good|3056,3060
dentition|3061,3070
<EOL>|3072,3073
NECK|3073,3077
:|3077,3078
nontender|3079,3088
supple|3089,3095
neck|3096,3100
,|3100,3101
no|3102,3104
LAD|3105,3108
,|3108,3109
no|3110,3112
JVD|3113,3116
<EOL>|3118,3119
CARDIAC|3119,3126
:|3126,3127
RRR|3128,3131
,|3131,3132
S1|3133,3135
/|3135,3136
S2|3136,3138
,|3138,3139
no|3140,3142
murmurs|3143,3150
,|3150,3151
gallops|3152,3159
,|3159,3160
or|3161,3163
rubs|3164,3168
<EOL>|3170,3171
LUNG|3171,3175
:|3175,3176
CTAB|3177,3181
,|3181,3182
no|3183,3185
wheezes|3186,3193
,|3193,3194
rales|3195,3200
,|3200,3201
rhonchi|3202,3209
,|3209,3210
breathing|3211,3220
comfortably|3221,3232
<EOL>|3233,3234
without|3234,3241
use|3242,3245
of|3246,3248
accessory|3249,3258
muscles|3259,3266
<EOL>|3268,3269
ABDOMEN|3269,3276
:|3276,3277
soft|3278,3282
,|3282,3283
decreased|3284,3293
distension|3294,3304
,|3304,3305
not|3306,3309
tense|3310,3315
.|3315,3316
NABS|3317,3321
,|3321,3322
nontender|3323,3332
<EOL>|3334,3335
<EOL>|3335,3336
EXTREMITIES|3336,3347
:|3347,3348
no|3349,3351
cyanosis|3352,3360
,|3360,3361
clubbing|3362,3370
or|3371,3373
edema|3374,3379
,|3379,3380
moving|3381,3387
all|3388,3391
4|3392,3393
<EOL>|3394,3395
extremities|3395,3406
with|3407,3411
purpose|3412,3419
<EOL>|3419,3420
PULSES|3420,3426
:|3426,3427
2|3428,3429
+|3429,3430
DP|3431,3433
pulses|3434,3440
bilaterally|3441,3452
<EOL>|3454,3455
NEURO|3455,3460
:|3460,3461
CN|3462,3464
II|3465,3467
-|3467,3468
XII|3468,3471
intact|3472,3478
,|3478,3479
AAO3|3480,3484
,|3484,3485
no|3486,3488
asterxis|3489,3497
<EOL>|3499,3500
SKIN|3500,3504
:|3504,3505
warm|3506,3510
and|3511,3514
well|3515,3519
perfused|3520,3528
,|3528,3529
no|3530,3532
excoriations|3533,3545
or|3546,3548
lesions|3549,3556
,|3556,3557
no|3558,3560
<EOL>|3561,3562
rashes|3562,3568
<EOL>|3568,3569
<EOL>|3570,3571
Pertinent|3571,3580
Results|3581,3588
:|3588,3589
<EOL>|3589,3590
ADMISSION|3590,3599
LABS|3600,3604
<EOL>|3604,3605
=|3605,3606
=|3606,3607
=|3607,3608
=|3608,3609
=|3609,3610
=|3610,3611
=|3611,3612
=|3612,3613
=|3613,3614
=|3614,3615
=|3615,3616
=|3616,3617
=|3617,3618
=|3618,3619
<EOL>|3619,3620
_|3620,3621
_|3621,3622
_|3622,3623
09|3624,3626
:|3626,3627
20PM|3627,3631
BLOOD|3632,3637
WBC|3638,3641
-|3641,3642
8|3642,3643
.|3643,3644
2|3644,3645
#|3645,3646
RBC|3647,3650
-|3650,3651
3|3651,3652
.|3652,3653
48|3653,3655
*|3655,3656
Hgb|3657,3660
-|3660,3661
12.3|3661,3665
Hct|3666,3669
-|3669,3670
36.7|3670,3674
<EOL>|3675,3676
MCV|3676,3679
-|3679,3680
106|3680,3683
*|3683,3684
MCH|3685,3688
-|3688,3689
35|3689,3691
.|3691,3692
5|3692,3693
*|3693,3694
MCHC|3695,3699
-|3699,3700
33.6|3700,3704
RDW|3705,3708
-|3708,3709
16|3709,3711
.|3711,3712
5|3712,3713
*|3713,3714
Plt|3715,3718
_|3719,3720
_|3720,3721
_|3721,3722
<EOL>|3722,3723
_|3723,3724
_|3724,3725
_|3725,3726
09|3727,3729
:|3729,3730
28PM|3730,3734
BLOOD|3735,3740
_|3741,3742
_|3742,3743
_|3743,3744
PTT|3745,3748
-|3748,3749
31.8|3749,3753
_|3754,3755
_|3755,3756
_|3756,3757
<EOL>|3757,3758
_|3758,3759
_|3759,3760
_|3760,3761
09|3762,3764
:|3764,3765
20PM|3765,3769
BLOOD|3770,3775
Glucose|3776,3783
-|3783,3784
118|3784,3787
*|3787,3788
UreaN|3789,3794
-|3794,3795
33|3795,3797
*|3797,3798
Creat|3799,3804
-|3804,3805
0.6|3805,3808
Na|3809,3811
-|3811,3812
127|3812,3815
*|3815,3816
<EOL>|3817,3818
K|3818,3819
-|3819,3820
5|3820,3821
.|3821,3822
3|3822,3823
*|3823,3824
Cl|3825,3827
-|3827,3828
97|3828,3830
HCO3|3831,3835
-|3835,3836
24|3836,3838
AnGap|3839,3844
-|3844,3845
11|3845,3847
<EOL>|3847,3848
_|3848,3849
_|3849,3850
_|3850,3851
09|3852,3854
:|3854,3855
20PM|3855,3859
BLOOD|3860,3865
ALT|3866,3869
-|3869,3870
135|3870,3873
*|3873,3874
AST|3875,3878
-|3878,3879
244|3879,3882
*|3882,3883
AlkPhos|3884,3891
-|3891,3892
123|3892,3895
*|3895,3896
<EOL>|3897,3898
TotBili|3898,3905
-|3905,3906
1.3|3906,3909
<EOL>|3909,3910
_|3910,3911
_|3911,3912
_|3912,3913
09|3914,3916
:|3916,3917
20PM|3917,3921
BLOOD|3922,3927
Albumin|3928,3935
-|3935,3936
3.5|3936,3939
Calcium|3940,3947
-|3947,3948
8|3948,3949
.|3949,3950
3|3950,3951
*|3951,3952
Phos|3953,3957
-|3957,3958
3.3|3958,3961
Mg|3962,3964
-|3964,3965
2.3|3965,3968
<EOL>|3968,3969
_|3969,3970
_|3970,3971
_|3971,3972
09|3973,3975
:|3975,3976
27PM|3976,3980
BLOOD|3981,3986
Lactate|3987,3994
-|3994,3995
2|3995,3996
.|3996,3997
1|3997,3998
*|3998,3999
<EOL>|3999,4000
<EOL>|4000,4001
NOTABLE|4001,4008
LABS|4009,4013
<EOL>|4013,4014
=|4014,4015
=|4015,4016
=|4016,4017
=|4017,4018
=|4018,4019
=|4019,4020
=|4020,4021
=|4021,4022
=|4022,4023
=|4023,4024
=|4024,4025
=|4025,4026
<EOL>|4026,4027
_|4027,4028
_|4028,4029
_|4029,4030
12|4031,4033
:|4033,4034
30AM|4034,4038
ASCITES|4039,4046
WBC|4047,4050
-|4050,4051
220|4051,4054
*|4054,4055
_|4056,4057
_|4057,4058
_|4058,4059
Polys|4060,4065
-|4065,4066
17|4066,4068
*|4068,4069
<EOL>|4070,4071
Lymphs|4071,4077
-|4077,4078
48|4078,4080
*|4080,4081
Monos|4082,4087
-|4087,4088
19|4088,4090
*|4090,4091
Mesothe|4092,4099
-|4099,4100
2|4100,4101
*|4101,4102
Macroph|4103,4110
-|4110,4111
12|4111,4113
*|4113,4114
Other|4115,4120
-|4120,4121
2|4121,4122
*|4122,4123
<EOL>|4123,4124
_|4124,4125
_|4125,4126
_|4126,4127
12|4128,4130
:|4130,4131
30AM|4131,4135
ASCITES|4136,4143
TotPro|4144,4150
-|4150,4151
0.7|4151,4154
Glucose|4155,4162
-|4162,4163
129|4163,4166
<EOL>|4166,4167
<EOL>|4167,4168
MICROBIOLOGY|4168,4180
<EOL>|4180,4181
=|4181,4182
=|4182,4183
=|4183,4184
=|4184,4185
=|4185,4186
=|4186,4187
=|4187,4188
=|4188,4189
=|4189,4190
=|4190,4191
=|4191,4192
=|4192,4193
<EOL>|4193,4194
_|4194,4195
_|4195,4196
_|4196,4197
12|4198,4200
:|4200,4201
30|4201,4203
am|4204,4206
PERITONEAL|4207,4217
FLUID|4218,4223
<EOL>|4223,4224
<EOL>|4224,4225
GRAM|4228,4232
STAIN|4233,4238
(|4239,4240
Final|4240,4245
_|4246,4247
_|4247,4248
_|4248,4249
:|4249,4250
<EOL>|4251,4252
NO|4258,4260
POLYMORPHONUCLEAR|4261,4278
LEUKOCYTES|4279,4289
SEEN|4290,4294
.|4294,4295
<EOL>|4296,4297
NO|4303,4305
MICROORGANISMS|4306,4320
SEEN|4321,4325
.|4325,4326
<EOL>|4327,4328
<EOL>|4328,4329
FLUID|4332,4337
CULTURE|4338,4345
(|4346,4347
Final|4347,4352
_|4353,4354
_|4354,4355
_|4355,4356
:|4356,4357
NO|4361,4363
GROWTH|4364,4370
.|4370,4371
<EOL>|4372,4373
<EOL>|4373,4374
ANAEROBIC|4377,4386
CULTURE|4387,4394
(|4395,4396
Preliminary|4396,4407
)|4407,4408
:|4408,4409
NO|4413,4415
GROWTH|4416,4422
.|4422,4423
<EOL>|4423,4424
<EOL>|4424,4425
_|4425,4426
_|4426,4427
_|4427,4428
VRE|4429,4432
screen|4433,4439
:|4439,4440
No|4441,4443
VRE|4444,4447
isolated|4448,4456
.|4456,4457
<EOL>|4457,4458
<EOL>|4458,4459
IMAGING|4459,4466
/|4466,4467
STUDIES|4467,4474
<EOL>|4474,4475
=|4475,4476
=|4476,4477
=|4477,4478
=|4478,4479
=|4479,4480
=|4480,4481
=|4481,4482
=|4482,4483
=|4483,4484
=|4484,4485
=|4485,4486
=|4486,4487
=|4487,4488
=|4488,4489
=|4489,4490
<EOL>|4490,4491
CXR|4491,4494
_|4495,4496
_|4496,4497
_|4497,4498
<EOL>|4498,4499
No|4499,4501
acute|4502,4507
cardiopulmonary|4508,4523
process|4524,4531
.|4531,4532
<EOL>|4532,4533
<EOL>|4533,4534
RUQUS|4534,4539
_|4540,4541
_|4541,4542
_|4542,4543
<EOL>|4543,4544
Cirrhotic|4544,4553
,|4553,4554
mild|4555,4559
splenomegaly|4560,4572
and|4573,4576
ascites|4577,4584
.|4584,4585
A|4587,4588
solid|4589,4594
3cm|4595,4598
nodule|4599,4605
in|4606,4608
<EOL>|4609,4610
the|4610,4613
left|4614,4618
lobe|4619,4623
of|4624,4626
the|4627,4630
liver|4631,4636
is|4637,4639
stable|4640,4646
in|4647,4649
size|4650,4654
and|4655,4658
appearance|4659,4669
.|4669,4670
<EOL>|4671,4672
<EOL>|4672,4673
DISCHARGE|4673,4682
LABS|4683,4687
<EOL>|4687,4688
=|4688,4689
=|4689,4690
=|4690,4691
=|4691,4692
=|4692,4693
=|4693,4694
=|4694,4695
=|4695,4696
=|4696,4697
=|4697,4698
=|4698,4699
=|4699,4700
=|4700,4701
=|4701,4702
<EOL>|4702,4703
_|4703,4704
_|4704,4705
_|4705,4706
06|4707,4709
:|4709,4710
15AM|4710,4714
BLOOD|4715,4720
WBC|4721,4724
-|4724,4725
5.6|4725,4728
RBC|4729,4732
-|4732,4733
3|4733,4734
.|4734,4735
27|4735,4737
*|4737,4738
Hgb|4739,4742
-|4742,4743
11|4743,4745
.|4745,4746
6|4746,4747
*|4747,4748
Hct|4749,4752
-|4752,4753
33|4753,4755
.|4755,4756
5|4756,4757
*|4757,4758
<EOL>|4759,4760
MCV|4760,4763
-|4763,4764
103|4764,4767
*|4767,4768
MCH|4769,4772
-|4772,4773
35|4773,4775
.|4775,4776
5|4776,4777
*|4777,4778
MCHC|4779,4783
-|4783,4784
34.5|4784,4788
RDW|4789,4792
-|4792,4793
16|4793,4795
.|4795,4796
1|4796,4797
*|4797,4798
Plt|4799,4802
_|4803,4804
_|4804,4805
_|4805,4806
<EOL>|4806,4807
_|4807,4808
_|4808,4809
_|4809,4810
06|4811,4813
:|4813,4814
15AM|4814,4818
BLOOD|4819,4824
_|4825,4826
_|4826,4827
_|4827,4828
PTT|4829,4832
-|4832,4833
36.0|4833,4837
_|4838,4839
_|4839,4840
_|4840,4841
<EOL>|4841,4842
_|4842,4843
_|4843,4844
_|4844,4845
06|4846,4848
:|4848,4849
15AM|4849,4853
BLOOD|4854,4859
Glucose|4860,4867
-|4867,4868
87|4868,4870
UreaN|4871,4876
-|4876,4877
29|4877,4879
*|4879,4880
Creat|4881,4886
-|4886,4887
0.4|4887,4890
Na|4891,4893
-|4893,4894
123|4894,4897
*|4897,4898
<EOL>|4899,4900
K|4900,4901
-|4901,4902
5|4902,4903
.|4903,4904
4|4904,4905
*|4905,4906
Cl|4907,4909
-|4909,4910
93|4910,4912
*|4912,4913
HCO3|4914,4918
-|4918,4919
24|4919,4921
AnGap|4922,4927
-|4927,4928
11|4928,4930
<EOL>|4930,4931
_|4931,4932
_|4932,4933
_|4933,4934
06|4935,4937
:|4937,4938
15AM|4938,4942
BLOOD|4943,4948
ALT|4949,4952
-|4952,4953
112|4953,4956
*|4956,4957
AST|4958,4961
-|4961,4962
176|4962,4965
*|4965,4966
AlkPhos|4967,4974
-|4974,4975
101|4975,4978
<EOL>|4979,4980
TotBili|4980,4987
-|4987,4988
2|4988,4989
.|4989,4990
8|4990,4991
*|4991,4992
<EOL>|4992,4993
_|4993,4994
_|4994,4995
_|4995,4996
06|4997,4999
:|4999,5000
15AM|5000,5004
BLOOD|5005,5010
Albumin|5011,5018
-|5018,5019
3.5|5019,5022
Calcium|5023,5030
-|5030,5031
8.8|5031,5034
Phos|5035,5039
-|5039,5040
3.4|5040,5043
Mg|5044,5046
-|5046,5047
2.|5047,5049
_|5049,5050
_|5050,5051
_|5051,5052
w|5053,5054
/|5054,5055
HIV|5056,5059
on|5060,5062
HAART|5063,5068
,|5068,5069
COPD|5070,5074
on|5075,5077
3L|5078,5080
home|5081,5085
O2|5086,5088
,|5088,5089
HCV|5090,5093
cirrhosis|5094,5103
<EOL>|5104,5105
decompensated|5105,5118
(|5119,5120
ascites|5120,5127
requiring|5128,5137
biweekly|5138,5146
therapeutic|5147,5158
<EOL>|5159,5160
paracenteses|5160,5172
,|5172,5173
hepatic|5174,5181
encephalopathy|5182,5196
;|5196,5197
not|5198,5201
on|5202,5204
transplant|5205,5215
list|5216,5220
_|5221,5222
_|5222,5223
_|5223,5224
<EOL>|5225,5226
<EOL>|5227,5228
comorbidities|5228,5241
)|5241,5242
p|5243,5244
/|5244,5245
w|5245,5246
worsening|5247,5256
abd|5257,5260
girth|5261,5266
and|5267,5270
pain|5271,5275
.|5275,5276
<EOL>|5276,5277
<EOL>|5277,5278
#|5278,5279
Goals|5280,5285
of|5286,5288
care|5289,5293
:|5293,5294
The|5296,5299
patient|5300,5307
expressed|5308,5317
that|5318,5322
her|5323,5326
desire|5327,5333
to|5334,5336
"|5337,5338
let|5338,5341
<EOL>|5342,5343
go|5343,5345
"|5345,5346
and|5347,5350
be|5351,5353
at|5354,5356
peace|5357,5362
.|5362,5363
She|5364,5367
is|5368,5370
tired|5371,5376
of|5377,5379
"|5380,5381
fighting|5381,5389
"|5389,5390
her|5391,5394
end|5395,5398
stage|5399,5404
<EOL>|5405,5406
liver|5406,5411
disease|5412,5419
and|5420,5423
does|5424,5428
not|5429,5432
feel|5433,5437
that|5438,5442
she|5443,5446
has|5447,5450
a|5451,5452
good|5453,5457
quality|5458,5465
of|5466,5468
<EOL>|5469,5470
life|5470,5474
.|5474,5475
She|5476,5479
wished|5480,5486
to|5487,5489
meet|5490,5494
with|5495,5499
a|5500,5501
representative|5502,5516
from|5517,5521
hospice|5522,5529
,|5529,5530
<EOL>|5531,5532
which|5532,5537
we|5538,5540
were|5541,5545
able|5546,5550
to|5551,5553
arrange|5554,5561
,|5561,5562
and|5563,5566
she|5567,5570
decided|5571,5578
that|5579,5583
she|5584,5587
would|5588,5593
<EOL>|5594,5595
like|5595,5599
to|5600,5602
go|5603,5605
home|5606,5610
with|5611,5615
hospice|5616,5623
.|5623,5624
A|5625,5626
conversation|5627,5639
was|5640,5643
held|5644,5648
with|5649,5653
the|5654,5657
<EOL>|5658,5659
patient|5659,5666
regarding|5667,5676
code|5677,5681
status|5682,5688
.|5688,5689
She|5690,5693
noted|5694,5699
that|5700,5704
she|5705,5708
would|5709,5714
probably|5715,5723
<EOL>|5724,5725
be|5725,5727
DNR|5728,5731
/|5731,5732
DNI|5732,5735
,|5735,5736
but|5737,5740
would|5741,5746
like|5747,5751
to|5752,5754
discuss|5755,5762
it|5763,5765
with|5766,5770
her|5771,5774
son|5775,5778
(|5779,5780
HCP|5780,5783
)|5783,5784
.|5784,5785
<EOL>|5786,5787
Therefore|5787,5796
,|5796,5797
at|5798,5800
this|5801,5805
time|5806,5810
,|5810,5811
she|5812,5815
remains|5816,5823
full|5824,5828
code|5829,5833
.|5833,5834
We|5835,5837
also|5838,5842
<EOL>|5843,5844
discussed|5844,5853
the|5854,5857
possibility|5858,5869
of|5870,5872
her|5873,5876
getting|5877,5884
a|5885,5886
pleurex|5887,5894
catheter|5895,5903
<EOL>|5904,5905
placed|5905,5911
because|5912,5919
of|5920,5922
her|5923,5926
repeated|5927,5935
paracenteses|5936,5948
.|5948,5949
She|5950,5953
was|5954,5957
discharged|5958,5968
<EOL>|5969,5970
to|5970,5972
home|5973,5977
with|5978,5982
hospice|5983,5990
on|5991,5993
_|5994,5995
_|5995,5996
_|5996,5997
.|5997,5998
<EOL>|5998,5999
<EOL>|5999,6000
#|6000,6001
Decompensated|6002,6015
HCV|6016,6019
cirrhosis|6020,6029
with|6030,6034
ascites|6035,6042
:|6042,6043
The|6044,6047
patient|6048,6055
<EOL>|6056,6057
presented|6057,6066
with|6067,6071
worsening|6072,6081
ascites|6082,6089
.|6089,6090
Her|6091,6094
pain|6095,6099
was|6100,6103
initially|6104,6113
managed|6114,6121
<EOL>|6122,6123
with|6123,6127
tramadol|6128,6136
and|6137,6140
morphine|6141,6149
.|6149,6150
She|6151,6154
underwent|6155,6164
_|6165,6166
_|6166,6167
_|6167,6168
paracentesis|6169,6181
<EOL>|6182,6183
on|6183,6185
_|6186,6187
_|6187,6188
_|6188,6189
with|6190,6194
removal|6195,6202
of|6203,6205
3.5|6206,6209
L|6209,6210
and|6211,6214
she|6215,6218
received|6219,6227
albumin|6228,6235
.|6235,6236
Studies|6237,6244
<EOL>|6245,6246
on|6246,6248
the|6249,6252
fluid|6253,6258
were|6259,6263
negative|6264,6272
,|6272,6273
and|6274,6277
she|6278,6281
reported|6282,6290
a|6291,6292
significant|6293,6304
<EOL>|6305,6306
improvement|6306,6317
in|6318,6320
her|6321,6324
pain|6325,6329
.|6329,6330
<EOL>|6330,6331
<EOL>|6332,6333
#|6333,6334
Hyperkalemia|6335,6347
:|6347,6348
During|6349,6355
her|6356,6359
hospitalization|6360,6375
,|6375,6376
it|6377,6379
was|6380,6383
noted|6384,6389
that|6390,6394
<EOL>|6395,6396
she|6396,6399
had|6400,6403
hyperkalemia|6404,6416
5.3|6417,6420
-|6421,6422
>|6422,6423
5.9|6424,6427
-|6428,6429
>|6429,6430
6.9|6431,6434
without|6435,6442
EKG|6443,6446
changes|6447,6454
.|6454,6455
<EOL>|6456,6457
After|6457,6462
treatment|6463,6472
with|6473,6477
calcium|6478,6485
gluconate|6486,6495
2gm|6496,6499
x2|6500,6502
,|6502,6503
insulin|6504,6511
and|6512,6515
D50|6516,6519
x|6520,6521
<EOL>|6522,6523
2|6523,6524
,|6524,6525
and|6526,6529
kayexelate|6530,6540
,|6540,6541
her|6542,6545
K|6546,6547
downtrended|6548,6559
to|6560,6562
5.4|6563,6566
.|6566,6567
Her|6568,6571
K|6572,6573
has|6574,6577
been|6578,6582
<EOL>|6583,6584
persistently|6584,6596
elevated|6597,6605
in|6606,6608
the|6609,6612
past|6613,6617
and|6618,6621
should|6622,6628
continue|6629,6637
to|6638,6640
be|6641,6643
<EOL>|6644,6645
monitored|6645,6654
.|6654,6655
<EOL>|6655,6656
<EOL>|6656,6657
#|6657,6658
Hepatic|6659,6666
encephalopathy|6667,6681
:|6681,6682
The|6683,6686
patient|6687,6694
's|6694,6696
mental|6697,6703
status|6704,6710
was|6711,6714
A|6715,6716
+|6716,6717
Ox3|6717,6720
<EOL>|6721,6722
on|6722,6724
admission|6725,6734
.|6734,6735
She|6736,6739
was|6740,6743
continued|6744,6753
on|6754,6756
rifaximin|6757,6766
and|6767,6770
lactulose|6771,6780
<EOL>|6781,6782
in|6782,6784
-|6784,6785
house|6785,6790
and|6791,6794
at|6795,6797
discharge|6798,6807
.|6807,6808
<EOL>|6808,6809
<EOL>|6809,6810
CHRONIC|6810,6817
ISSUES|6818,6824
<EOL>|6824,6825
=|6825,6826
=|6826,6827
=|6827,6828
=|6828,6829
=|6829,6830
=|6830,6831
=|6831,6832
=|6832,6833
=|6833,6834
=|6834,6835
=|6835,6836
=|6836,6837
=|6837,6838
=|6838,6839
<EOL>|6839,6840
<EOL>|6840,6841
#|6841,6842
Hyponatremia|6843,6855
-|6856,6857
The|6858,6861
patient|6862,6869
has|6870,6873
a|6874,6875
history|6876,6883
of|6884,6886
asymptomatic|6887,6899
<EOL>|6900,6901
hyponatremia|6901,6913
.|6913,6914
It|6915,6917
is|6918,6920
most|6921,6925
likely|6926,6932
hypervolemic|6933,6945
hyponatremia|6946,6958
<EOL>|6959,6960
related|6960,6967
to|6968,6970
underlying|6971,6981
liver|6982,6987
disease|6988,6995
as|6996,6998
well|6999,7003
as|7004,7006
aldosterone|7007,7018
axis|7019,7023
<EOL>|7024,7025
dysfunction|7025,7036
related|7037,7044
to|7045,7047
liver|7048,7053
disease|7054,7061
.|7061,7062
She|7063,7066
remained|7067,7075
asymptomatic|7076,7088
<EOL>|7089,7090
through|7090,7097
her|7098,7101
hospitalization|7102,7117
.|7117,7118
Because|7119,7126
she|7127,7130
was|7131,7134
also|7135,7139
started|7140,7147
on|7148,7150
<EOL>|7151,7152
10mg|7152,7156
of|7157,7159
furosemide|7160,7170
to|7171,7173
help|7174,7178
prevent|7179,7186
fluid|7187,7192
re-accumulation|7193,7208
,|7208,7209
she|7210,7213
<EOL>|7214,7215
will|7215,7219
require|7220,7227
BMPs|7228,7232
twice|7233,7238
weekly|7239,7245
in|7246,7248
the|7249,7252
outpatient|7253,7263
setting|7264,7271
.|7271,7272
<EOL>|7272,7273
<EOL>|7273,7274
#|7274,7275
HIV|7276,7279
:|7279,7280
Emtricitabine|7281,7294
-|7294,7295
Tenofovir|7295,7304
(|7305,7306
Truvada|7306,7313
)|7313,7314
and|7315,7318
Raltegravir|7319,7330
were|7331,7335
<EOL>|7336,7337
continued|7337,7346
in|7347,7349
-|7349,7350
house|7350,7355
and|7356,7359
at|7360,7362
discharge|7363,7372
.|7372,7373
<EOL>|7375,7376
<EOL>|7376,7377
#|7377,7378
COPD|7379,7383
:|7383,7384
fluticasone|7385,7396
,|7396,7397
tiotropium|7398,7408
and|7409,7412
albuterol|7413,7422
were|7423,7427
continued|7428,7437
<EOL>|7438,7439
in|7439,7441
-|7441,7442
house|7442,7447
and|7448,7451
at|7452,7454
discharge|7455,7464
.|7464,7465
<EOL>|7465,7466
<EOL>|7466,7467
TRANSITIONAL|7467,7479
ISSUES|7480,7486
<EOL>|7486,7487
=|7487,7488
=|7488,7489
=|7489,7490
=|7490,7491
=|7491,7492
=|7492,7493
=|7493,7494
=|7494,7495
=|7495,7496
=|7496,7497
=|7497,7498
=|7498,7499
=|7499,7500
=|7500,7501
=|7501,7502
=|7502,7503
=|7503,7504
=|7504,7505
=|7505,7506
<EOL>|7506,7507
[|7507,7508
]|7509,7510
Follow|7511,7517
-|7517,7518
up|7518,7520
peritoneal|7521,7531
fluid|7532,7537
culture|7538,7545
<EOL>|7545,7546
[|7546,7547
]|7548,7549
New|7550,7553
/|7553,7554
changed|7554,7561
medications|7562,7573
:|7573,7574
Furosemide|7575,7585
10mg|7586,7590
daily|7591,7596
(|7597,7598
new|7598,7601
)|7601,7602
<EOL>|7602,7603
[|7603,7604
]|7605,7606
For|7607,7610
hyperkalemia|7611,7623
and|7624,7627
hyponatremia|7628,7640
,|7640,7641
the|7642,7645
patient|7646,7653
should|7654,7660
have|7661,7665
<EOL>|7666,7667
biweekly|7667,7675
BMPs|7676,7680
(|7681,7682
script|7682,7688
written|7689,7696
)|7696,7697
.|7697,7698
If|7699,7701
K|7702,7703
>|7704,7705
5.3|7706,7709
,|7709,7710
she|7711,7714
should|7715,7721
be|7722,7724
given|7725,7730
<EOL>|7731,7732
kayexelate|7732,7742
once|7743,7747
weekly|7748,7754
.|7754,7755
Lab|7756,7759
results|7760,7767
will|7768,7772
be|7773,7775
faxed|7776,7781
/|7781,7782
sent|7782,7786
to|7787,7789
Dr|7790,7792
.|7792,7793
<EOL>|7794,7795
_|7795,7796
_|7796,7797
_|7797,7798
.|7798,7799
<EOL>|7799,7800
[|7800,7801
]|7802,7803
Continue|7804,7812
conversation|7813,7825
regarding|7826,7835
pleurex|7836,7843
catheter|7844,7852
placement|7853,7862
<EOL>|7863,7864
and|7864,7867
code|7868,7872
status|7873,7879
.|7879,7880
<EOL>|7880,7881
[|7881,7882
]|7883,7884
She|7885,7888
will|7889,7893
continue|7894,7902
to|7903,7905
have|7906,7910
twice|7911,7916
weekly|7917,7923
paracenteses|7924,7936
<EOL>|7936,7937
<EOL>|7937,7938
#|7938,7939
Code|7940,7944
:|7944,7945
full|7946,7950
<EOL>|7952,7953
#|7953,7954
Emergency|7955,7964
Contact|7965,7972
:|7972,7973
_|7974,7975
_|7975,7976
_|7976,7977
_|7978,7979
_|7979,7980
_|7980,7981
<EOL>|7982,7983
<EOL>|7984,7985
_|7985,7986
_|7986,7987
_|7987,7988
on|7989,7991
Admission|7992,8001
:|8001,8002
<EOL>|8002,8003
The|8003,8006
Preadmission|8007,8019
Medication|8020,8030
list|8031,8035
is|8036,8038
accurate|8039,8047
and|8048,8051
complete|8052,8060
.|8060,8061
<EOL>|8061,8062
1|8062,8063
.|8063,8064
Calcium|8065,8072
Carbonate|8073,8082
500|8083,8086
mg|8087,8089
PO|8090,8092
BID|8093,8096
<EOL>|8097,8098
2.|8098,8100
Emtricitabine|8101,8114
-|8114,8115
Tenofovir|8115,8124
(|8125,8126
Truvada|8126,8133
)|8133,8134
1|8135,8136
TAB|8137,8140
PO|8141,8143
DAILY|8144,8149
<EOL>|8150,8151
3.|8151,8153
Fluticasone|8154,8165
Propionate|8166,8176
110mcg|8177,8183
1|8184,8185
PUFF|8186,8190
IH|8191,8193
BID|8194,8197
<EOL>|8198,8199
4.|8199,8201
Lactulose|8202,8211
30|8212,8214
mL|8215,8217
PO|8218,8220
TID|8221,8224
<EOL>|8225,8226
5.|8226,8228
Raltegravir|8229,8240
400|8241,8244
mg|8245,8247
PO|8248,8250
BID|8251,8254
<EOL>|8255,8256
6.|8256,8258
Rifaximin|8259,8268
550|8269,8272
mg|8273,8275
PO|8276,8278
BID|8279,8282
<EOL>|8283,8284
7.|8284,8286
TraMADOL|8287,8295
(|8296,8297
Ultram|8297,8303
)|8303,8304
_|8305,8306
_|8306,8307
_|8307,8308
mg|8309,8311
PO|8312,8314
Q6H|8315,8318
:|8318,8319
PRN|8319,8322
pain|8323,8327
<EOL>|8328,8329
8.|8329,8331
albuterol|8332,8341
sulfate|8342,8349
90|8350,8352
mcg|8353,8356
/|8356,8357
actuation|8357,8366
inhalation|8367,8377
Q6H|8378,8381
:|8381,8382
PRN|8382,8385
<EOL>|8386,8387
Wheezing|8387,8395
<EOL>|8396,8397
9.|8397,8399
Tiotropium|8400,8410
Bromide|8411,8418
1|8419,8420
CAP|8421,8424
IH|8425,8427
DAILY|8428,8433
<EOL>|8434,8435
<EOL>|8435,8436
<EOL>|8437,8438
Discharge|8438,8447
Medications|8448,8459
:|8459,8460
<EOL>|8460,8461
1.|8461,8463
albuterol|8464,8473
sulfate|8474,8481
90|8482,8484
mcg|8485,8488
/|8488,8489
actuation|8489,8498
inhalation|8499,8509
Q6H|8510,8513
:|8513,8514
PRN|8514,8517
<EOL>|8518,8519
Wheezing|8519,8527
<EOL>|8528,8529
2|8529,8530
.|8530,8531
Calcium|8532,8539
Carbonate|8540,8549
500|8550,8553
mg|8554,8556
PO|8557,8559
BID|8560,8563
<EOL>|8564,8565
3.|8565,8567
Emtricitabine|8568,8581
-|8581,8582
Tenofovir|8582,8591
(|8592,8593
Truvada|8593,8600
)|8600,8601
1|8602,8603
TAB|8604,8607
PO|8608,8610
DAILY|8611,8616
<EOL>|8617,8618
4.|8618,8620
Fluticasone|8621,8632
Propionate|8633,8643
110mcg|8644,8650
1|8651,8652
PUFF|8653,8657
IH|8658,8660
BID|8661,8664
<EOL>|8665,8666
5.|8666,8668
Lactulose|8669,8678
30|8679,8681
mL|8682,8684
PO|8685,8687
TID|8688,8691
<EOL>|8692,8693
6.|8693,8695
Raltegravir|8696,8707
400|8708,8711
mg|8712,8714
PO|8715,8717
BID|8718,8721
<EOL>|8722,8723
7.|8723,8725
Rifaximin|8726,8735
550|8736,8739
mg|8740,8742
PO|8743,8745
BID|8746,8749
<EOL>|8750,8751
8.|8751,8753
Tiotropium|8754,8764
Bromide|8765,8772
1|8773,8774
CAP|8775,8778
IH|8779,8781
DAILY|8782,8787
<EOL>|8788,8789
9.|8789,8791
TraMADOL|8792,8800
(|8801,8802
Ultram|8802,8808
)|8808,8809
_|8810,8811
_|8811,8812
_|8812,8813
mg|8814,8816
PO|8817,8819
Q6H|8820,8823
:|8823,8824
PRN|8824,8827
pain|8828,8832
<EOL>|8833,8834
10|8834,8836
.|8836,8837
Furosemide|8838,8848
10|8849,8851
mg|8852,8854
PO|8855,8857
DAILY|8858,8863
<EOL>|8864,8865
RX|8865,8867
*|8868,8869
furosemide|8869,8879
20|8880,8882
mg|8883,8885
0.5|8886,8889
(|8890,8891
One|8891,8894
half|8895,8899
)|8899,8900
tablet|8901,8907
(|8907,8908
s|8908,8909
)|8909,8910
by|8911,8913
mouth|8914,8919
Please|8920,8926
<EOL>|8927,8928
take|8928,8932
1|8933,8934
tablet|8935,8941
daily|8942,8947
.|8947,8948
Disp|8949,8953
#|8954,8955
*|8955,8956
15|8956,8958
Tablet|8959,8965
Refills|8966,8973
:|8973,8974
*|8974,8975
0|8975,8976
<EOL>|8976,8977
11.|8977,8980
Outpatient|8981,8991
Lab|8992,8995
Work|8996,9000
<EOL>|9000,9001
Please|9001,9007
obtain|9008,9014
biweekly|9015,9023
BMP|9024,9027
to|9028,9030
monitor|9031,9038
K|9039,9040
and|9041,9044
Na|9045,9047
.|9047,9048
Please|9049,9055
fax|9056,9059
<EOL>|9060,9061
results|9061,9068
to|9069,9071
Dr.|9072,9075
_|9076,9077
_|9077,9078
_|9078,9079
at|9080,9082
the|9083,9086
_|9087,9088
_|9088,9089
_|9089,9090
at|9091,9093
_|9094,9095
_|9095,9096
_|9096,9097
.|9097,9098
<EOL>|9098,9099
<EOL>|9099,9100
<EOL>|9101,9102
Discharge|9102,9111
Disposition|9112,9123
:|9123,9124
<EOL>|9124,9125
Home|9125,9129
With|9130,9134
Service|9135,9142
<EOL>|9142,9143
<EOL>|9144,9145
Facility|9145,9153
:|9153,9154
<EOL>|9154,9155
_|9155,9156
_|9156,9157
_|9157,9158
<EOL>|9158,9159
<EOL>|9160,9161
Discharge|9161,9170
Diagnosis|9171,9180
:|9180,9181
<EOL>|9181,9182
PRIMARY|9182,9189
DIAGNOSIS|9190,9199
<EOL>|9199,9200
=|9200,9201
=|9201,9202
=|9202,9203
=|9203,9204
=|9204,9205
=|9205,9206
=|9206,9207
=|9207,9208
=|9208,9209
=|9209,9210
=|9210,9211
=|9211,9212
=|9212,9213
=|9213,9214
=|9214,9215
=|9215,9216
=|9216,9217
<EOL>|9217,9218
-|9218,9219
Decompensated|9219,9232
HCV|9233,9236
cirrhosis|9237,9246
<EOL>|9246,9247
-|9247,9248
Hyperkalemia|9248,9260
<EOL>|9260,9261
<EOL>|9261,9262
SECONDARY|9262,9271
DIAGNOSES|9272,9281
<EOL>|9281,9282
=|9282,9283
=|9283,9284
=|9284,9285
=|9285,9286
=|9286,9287
=|9287,9288
=|9288,9289
=|9289,9290
=|9290,9291
=|9291,9292
=|9292,9293
=|9293,9294
=|9294,9295
=|9295,9296
=|9296,9297
=|9297,9298
=|9298,9299
=|9299,9300
=|9300,9301
<EOL>|9301,9302
-|9302,9303
HIV|9303,9306
<EOL>|9306,9307
-|9307,9308
COPD|9308,9312
<EOL>|9312,9313
-|9313,9314
Hyponatremia|9314,9326
<EOL>|9326,9327
<EOL>|9327,9328
<EOL>|9329,9330
Discharge|9330,9339
Condition|9340,9349
:|9349,9350
<EOL>|9350,9351
Mental|9351,9357
Status|9358,9364
:|9364,9365
Clear|9366,9371
and|9372,9375
coherent|9376,9384
.|9384,9385
<EOL>|9385,9386
Level|9386,9391
of|9392,9394
Consciousness|9395,9408
:|9408,9409
Alert|9410,9415
and|9416,9419
interactive|9420,9431
.|9431,9432
<EOL>|9432,9433
Activity|9433,9441
Status|9442,9448
:|9448,9449
Ambulatory|9450,9460
-|9461,9462
Independent|9463,9474
.|9474,9475
<EOL>|9475,9476
<EOL>|9476,9477
<EOL>|9478,9479
Discharge|9479,9488
Instructions|9489,9501
:|9501,9502
<EOL>|9502,9503
Dear|9503,9507
Ms.|9508,9511
_|9512,9513
_|9513,9514
_|9514,9515
,|9515,9516
<EOL>|9516,9517
<EOL>|9517,9518
It|9518,9520
was|9521,9524
a|9525,9526
pleasure|9527,9535
caring|9536,9542
for|9543,9546
you|9547,9550
during|9551,9557
your|9558,9562
stay|9563,9567
at|9568,9570
_|9571,9572
_|9572,9573
_|9573,9574
.|9574,9575
You|9576,9579
<EOL>|9580,9581
were|9581,9585
admitted|9586,9594
because|9595,9602
of|9603,9605
worsening|9606,9615
abdominal|9616,9625
pain|9626,9630
.|9630,9631
It|9632,9634
is|9635,9637
likely|9638,9644
<EOL>|9645,9646
that|9646,9650
this|9651,9655
pain|9656,9660
was|9661,9664
due|9665,9668
to|9669,9671
increasing|9672,9682
fluid|9683,9688
in|9689,9691
the|9692,9695
abdomen|9696,9703
from|9704,9708
<EOL>|9709,9710
your|9710,9714
cirrhosis|9715,9724
.|9724,9725
After|9726,9731
a|9732,9733
paracentesis|9734,9746
in|9747,9749
which|9750,9755
much|9756,9760
of|9761,9763
this|9764,9768
fluid|9769,9774
<EOL>|9775,9776
was|9776,9779
removed|9780,9787
,|9787,9788
your|9789,9793
pain|9794,9798
improved|9799,9807
significantly|9808,9821
.|9821,9822
You|9823,9826
were|9827,9831
noted|9832,9837
to|9838,9840
<EOL>|9841,9842
have|9842,9846
a|9847,9848
high|9849,9853
potassium|9854,9863
during|9864,9870
your|9871,9875
hospitalization|9876,9891
,|9891,9892
which|9893,9898
came|9899,9903
<EOL>|9904,9905
down|9905,9909
with|9910,9914
treatment|9915,9924
but|9925,9928
this|9929,9933
should|9934,9940
continue|9941,9949
to|9950,9952
be|9953,9955
followed|9956,9964
as|9965,9967
<EOL>|9968,9969
an|9969,9971
outpatient|9972,9982
.|9982,9983
You|9984,9987
also|9988,9992
emphasized|9993,10003
your|10004,10008
desire|10009,10015
to|10016,10018
speak|10019,10024
with|10025,10029
a|10030,10031
<EOL>|10032,10033
representative|10033,10047
from|10048,10052
hospice|10053,10060
.|10060,10061
Because|10062,10069
of|10070,10072
your|10073,10077
repeated|10078,10086
<EOL>|10087,10088
paracenteses|10088,10100
,|10100,10101
we|10102,10104
also|10105,10109
discussed|10110,10119
the|10120,10123
possibility|10124,10135
of|10136,10138
a|10139,10140
pleurex|10141,10148
<EOL>|10149,10150
catheter|10150,10158
placement|10159,10168
.|10168,10169
We|10170,10172
arranged|10173,10181
for|10182,10185
you|10186,10189
to|10190,10192
meet|10193,10197
with|10198,10202
hospice|10203,10210
<EOL>|10211,10212
coordinators|10212,10224
,|10224,10225
and|10226,10229
you|10230,10233
will|10234,10238
be|10239,10241
discharged|10242,10252
home|10253,10257
with|10258,10262
hospice|10263,10270
.|10270,10271
<EOL>|10271,10272
<EOL>|10272,10273
We|10273,10275
wish|10276,10280
you|10281,10284
all|10285,10288
the|10289,10292
best|10293,10297
!|10297,10298
<EOL>|10298,10299
<EOL>|10299,10300
Your|10300,10304
_|10305,10306
_|10306,10307
_|10307,10308
care|10309,10313
team|10314,10318
<EOL>|10318,10319
<EOL>|10320,10321
Followup|10321,10329
Instructions|10330,10342
:|10342,10343
<EOL>|10343,10344
_|10344,10345
_|10345,10346
_|10346,10347
<EOL>|10347,10348

