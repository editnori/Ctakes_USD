 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|32,36
No|37,39
:|39,40
_|43,44
_|44,45
_|45,46
<EOL>|46,47
<EOL>|48,49
Admission|49,58
Date|59,63
:|63,64
_|66,67
_|67,68
_|68,69
Discharge|83,92
Date|93,97
:|97,98
_|101,102
_|102,103
_|103,104
<EOL>|104,105
<EOL>|106,107
Date|107,111
of|112,114
Birth|115,120
:|120,121
_|123,124
_|124,125
_|125,126
Sex|139,142
:|142,143
F|146,147
<EOL>|147,148
<EOL>|149,150
Service|150,157
:|157,158
MEDICINE|159,167
<EOL>|167,168
<EOL>|169,170
Penicillins|182,193
/|194,195
Dilantin|196,204
Kapseal|205,212
/|213,214
Zofran|215,221
(|222,223
as|223,225
hydrochloride|226,239
)|239,240
<EOL>|240,241
<EOL>|242,243
Attending|243,252
:|252,253
_|254,255
_|255,256
_|256,257
.|257,258
<EOL>|258,259
<EOL>|260,261
Right|278,283
hip|284,287
pain|288,292
<EOL>|293,294
<EOL>|295,296
Major|296,301
Surgical|302,310
or|311,313
Invasive|314,322
Procedure|323,332
:|332,333
<EOL>|333,334
None|334,338
<EOL>|338,339
<EOL>|339,340
<EOL>|341,342
_|370,371
_|371,372
_|372,373
is|374,376
a|377,378
_|379,380
_|380,381
_|381,382
y|383,384
/|384,385
o|385,386
F|387,388
with|389,393
PMHx|394,398
CHF|399,402
,|402,403
Afib|404,408
not|409,412
on|413,415
<EOL>|416,417
anticoagulation|417,432
,|432,433
severe|434,440
advanced|441,449
Alzheimer|450,459
's|459,461
dementia|462,470
,|470,471
<EOL>|472,473
osteoporosis|473,485
,|485,486
HTN|487,490
,|490,491
who|492,495
presents|496,504
from|505,509
assisted|510,518
living|519,525
facility|526,534
<EOL>|535,536
with|536,540
R|541,542
hip|543,546
pain|547,551
.|551,552
<EOL>|552,553
<EOL>|553,554
The|554,557
patient|558,565
has|566,569
severe|570,576
dementia|577,585
,|585,586
with|587,591
short|592,597
term|598,602
memory|603,609
loss|610,614
so|615,617
<EOL>|618,619
is|619,621
unable|622,628
to|629,631
provide|632,639
history|640,647
.|647,648
Much|649,653
of|654,656
the|657,660
history|661,668
is|669,671
obtained|672,680
<EOL>|681,682
from|682,686
multiple|687,695
family|696,702
members|703,710
in|711,713
the|714,717
room|718,722
.|722,723
She|724,727
has|728,731
multiple|732,740
<EOL>|741,742
family|742,748
members|749,756
who|757,760
live|761,765
close|766,771
by|772,774
and|775,778
are|779,782
involved|783,791
intimately|792,802
in|803,805
<EOL>|806,807
her|807,810
care|811,815
.|815,816
They|817,821
were|822,826
called|827,833
from|834,838
the|839,842
assisted|843,851
living|852,858
facility|859,867
<EOL>|868,869
this|869,873
morning|874,881
when|882,886
the|887,890
patient|891,898
was|899,902
in|903,905
_|906,907
_|907,908
_|908,909
right|910,915
hip|916,919
pain|920,924
.|924,925
This|926,930
<EOL>|931,932
occurred|932,940
suddenly|941,949
.|949,950
No|951,953
trauma|954,960
.|960,961
No|962,964
reported|965,973
falls|974,979
.|979,980
She|981,984
was|985,988
not|989,992
<EOL>|993,994
complaining|994,1005
of|1006,1008
other|1009,1014
symptoms|1015,1023
.|1023,1024
She|1025,1028
was|1029,1032
brought|1033,1040
to|1041,1043
the|1044,1047
ED|1048,1050
.|1050,1051
<EOL>|1052,1053
<EOL>|1053,1054
Discussing|1054,1064
with|1065,1069
the|1070,1073
patient|1074,1081
,|1081,1082
she|1083,1086
moved|1087,1092
into|1093,1097
the|1098,1101
Assisted|1102,1110
living|1111,1117
<EOL>|1118,1119
facility|1119,1127
in|1128,1130
_|1131,1132
_|1132,1133
_|1133,1134
in|1135,1137
_|1138,1139
_|1139,1140
_|1140,1141
given|1142,1147
worsening|1148,1157
of|1158,1160
her|1161,1164
<EOL>|1165,1166
dementia|1166,1174
.|1174,1175
She|1176,1179
was|1180,1183
in|1184,1186
her|1187,1190
USOH|1191,1195
,|1195,1196
bowling|1197,1204
weekly|1205,1211
and|1212,1215
very|1216,1220
social|1221,1227
,|1227,1228
<EOL>|1229,1230
until|1230,1235
_|1236,1237
_|1237,1238
_|1238,1239
when|1240,1244
she|1245,1248
developed|1249,1258
acute|1259,1264
SOB|1265,1268
with|1269,1273
ambulation|1274,1284
<EOL>|1285,1286
prompting|1286,1295
admission|1296,1305
to|1306,1308
_|1309,1310
_|1310,1311
_|1311,1312
where|1313,1318
she|1319,1322
was|1323,1326
noted|1327,1332
<EOL>|1333,1334
to|1334,1336
be|1337,1339
in|1340,1342
Afib|1343,1347
.|1347,1348
She|1349,1352
had|1353,1356
a|1357,1358
week|1359,1363
long|1364,1368
hospital|1369,1377
stay|1378,1382
complicated|1383,1394
by|1395,1397
<EOL>|1398,1399
an|1399,1401
ICU|1402,1405
course|1406,1412
for|1413,1416
an|1417,1419
allergic|1420,1428
reaction|1429,1437
to|1438,1440
a|1441,1442
medication|1443,1453
(|1454,1455
family|1455,1461
<EOL>|1462,1463
thinks|1463,1469
Zofran|1470,1476
)|1476,1477
.|1477,1478
Since|1479,1484
returning|1485,1494
from|1495,1499
this|1500,1504
hospitalization|1505,1520
,|1520,1521
she|1522,1525
<EOL>|1526,1527
has|1527,1530
not|1531,1534
been|1535,1539
back|1540,1544
to|1545,1547
baseline|1548,1556
and|1557,1560
has|1561,1564
deteriorated|1565,1577
.|1577,1578
She|1579,1582
has|1583,1586
<EOL>|1587,1588
spent|1588,1593
much|1594,1598
of|1599,1601
her|1602,1605
time|1606,1610
wheelchair|1611,1621
bound|1622,1627
given|1628,1633
deconditioning|1634,1648
.|1648,1649
<EOL>|1650,1651
She|1651,1654
has|1655,1658
worsening|1659,1668
memory|1669,1675
function|1676,1684
,|1684,1685
now|1686,1689
with|1690,1694
severe|1695,1701
short|1702,1707
term|1708,1712
<EOL>|1713,1714
memory|1714,1720
loss|1721,1725
.|1725,1726
Decreased|1727,1736
appetite|1737,1745
and|1746,1749
PO|1750,1752
intake|1753,1759
.|1759,1760
She|1761,1764
was|1765,1768
recently|1769,1777
<EOL>|1778,1779
seen|1779,1783
in|1784,1786
_|1787,1788
_|1788,1789
_|1789,1790
clinic|1791,1797
by|1798,1800
Dr.|1801,1804
_|1805,1806
_|1806,1807
_|1807,1808
new|1809,1812
diagnosis|1813,1822
of|1823,1825
CHF|1826,1829
.|1829,1830
She|1831,1834
<EOL>|1835,1836
underwent|1836,1845
an|1846,1848
TTE|1849,1852
at|1853,1855
_|1856,1857
_|1857,1858
_|1858,1859
yesterday|1860,1869
_|1870,1871
_|1871,1872
_|1872,1873
to|1874,1876
evaluate|1877,1885
her|1886,1889
<EOL>|1890,1891
systolic|1891,1899
function|1900,1908
.|1908,1909
<EOL>|1910,1911
<EOL>|1912,1913
In|1913,1915
the|1916,1919
ED|1920,1922
,|1922,1923
initial|1924,1931
vitals|1932,1938
were|1939,1943
:|1943,1944
<EOL>|1945,1946
98.7|1946,1950
,|1950,1951
96|1952,1954
,|1954,1955
122|1956,1959
/|1959,1960
48|1960,1962
,|1962,1963
20|1964,1966
,|1966,1967
96|1968,1970
%|1970,1971
RA|1972,1974
.|1974,1975
<EOL>|1976,1977
<EOL>|1977,1978
Exam|1978,1982
was|1983,1986
significant|1987,1998
for|1999,2002
:|2002,2003
<EOL>|2004,2005
R|2005,2006
hip|2007,2010
TTP|2011,2014
greater|2015,2022
trochanter|2023,2033
,|2033,2034
neg|2035,2038
straight|2039,2047
leg|2048,2051
raise|2052,2057
.|2057,2058
_|2059,2060
_|2060,2061
_|2061,2062
<EOL>|2063,2064
pulses|2064,2070
2|2071,2072
+|2072,2073
<EOL>|2073,2074
LLE|2074,2077
2|2078,2079
+|2079,2080
edema|2081,2086
,|2086,2087
unknown|2088,2095
duration|2096,2104
<EOL>|2104,2105
Labs|2105,2109
were|2110,2114
significant|2115,2126
for|2127,2130
:|2131,2132
<EOL>|2133,2134
K|2134,2135
2.8|2136,2139
<EOL>|2140,2141
Cr|2141,2143
0.8|2144,2147
<EOL>|2147,2148
CBC|2148,2151
:|2151,2152
13.9|2153,2157
/|2157,2158
12.5|2158,2162
/|2162,2163
39|2163,2165
.|2165,2166
2|2166,2167
/|2167,2168
168|2168,2171
<EOL>|2171,2172
UA|2172,2174
:|2174,2175
WBC|2176,2179
22|2180,2182
,|2182,2183
moderate|2184,2192
leuks|2193,2198
,|2198,2199
negative|2200,2208
nitrites|2209,2217
<EOL>|2218,2219
<EOL>|2219,2220
Studies|2220,2227
:|2227,2228
<EOL>|2229,2230
Lower|2230,2235
extremity|2236,2245
ultrasound|2246,2256
:|2256,2257
1.|2258,2260
Deep|2261,2265
vein|2266,2270
thrombosis|2271,2281
of|2282,2284
the|2285,2288
left|2289,2293
<EOL>|2294,2295
common|2295,2301
femoral|2302,2309
vein|2310,2314
extending|2315,2324
into|2325,2329
at|2330,2332
least|2333,2338
the|2339,2342
popliteal|2343,2352
vein|2353,2357
.|2357,2358
<EOL>|2359,2360
Left|2360,2364
calf|2365,2369
veins|2370,2375
were|2376,2380
not|2381,2384
clearly|2385,2392
identified|2393,2403
and|2404,2407
possibly|2408,2416
also|2417,2421
<EOL>|2422,2423
occluded|2423,2431
.|2431,2432
<EOL>|2432,2433
2|2433,2434
.|2434,2435
No|2436,2438
DVT|2439,2442
in|2443,2445
the|2446,2449
right|2450,2455
lower|2456,2461
extremity|2462,2471
.|2471,2472
<EOL>|2472,2473
<EOL>|2473,2474
CXR|2474,2477
<EOL>|2477,2478
Bilateral|2478,2487
pleural|2488,2495
effusions|2496,2505
,|2505,2506
large|2507,2512
on|2513,2515
the|2516,2519
right|2520,2525
and|2526,2529
small|2530,2535
on|2536,2538
the|2539,2542
<EOL>|2543,2544
left|2544,2548
.|2548,2549
No|2550,2552
definite|2553,2561
focal|2562,2567
consolidation|2568,2581
identified|2582,2592
,|2592,2593
although|2594,2602
<EOL>|2603,2604
evaluation|2604,2614
is|2615,2617
limited|2618,2625
secondary|2626,2635
to|2636,2638
these|2639,2644
effusions|2645,2654
.|2654,2655
<EOL>|2656,2657
<EOL>|2657,2658
She|2658,2661
was|2662,2665
given|2666,2671
80|2672,2674
mEq|2675,2678
of|2679,2681
K|2682,2683
and|2684,2687
60mg|2688,2692
Enoxaparin|2693,2703
Sodium|2704,2710
.|2710,2711
<EOL>|2712,2713
<EOL>|2715,2716
Vitals|2716,2722
on|2723,2725
transfer|2726,2734
were|2735,2739
:|2739,2740
97.9|2741,2745
,|2745,2746
79|2747,2749
,|2749,2750
125|2751,2754
/|2754,2755
53|2755,2757
,|2757,2758
18|2759,2761
,|2761,2762
100|2763,2766
%|2766,2767
Nasal|2768,2773
<EOL>|2774,2775
Cannula|2775,2782
.|2782,2783
<EOL>|2784,2785
<EOL>|2786,2787
On|2787,2789
the|2790,2793
floor|2794,2799
,|2799,2800
she|2801,2804
is|2805,2807
resting|2808,2815
comfortably|2816,2827
in|2828,2830
bed|2831,2834
.|2834,2835
History|2836,2843
is|2844,2846
<EOL>|2847,2848
obtained|2848,2856
as|2857,2859
above|2860,2865
with|2866,2870
family|2871,2877
members|2878,2885
.|2885,2886
She|2887,2890
sleeps|2891,2897
with|2898,2902
2|2903,2904
pillows|2905,2912
<EOL>|2913,2914
at|2914,2916
home|2917,2921
and|2922,2925
has|2926,2929
DOE|2930,2933
.|2933,2934
She|2935,2938
has|2939,2942
not|2943,2946
had|2947,2950
a|2951,2952
bowel|2953,2958
movement|2959,2967
in|2968,2970
2|2971,2972
days|2973,2977
.|2977,2978
<EOL>|2979,2980
<EOL>|2980,2981
<EOL>|2981,2982
Review|2982,2988
of|2989,2991
systems|2992,2999
:|2999,3000
<EOL>|3002,3003
(|3003,3004
+|3004,3005
)|3005,3006
Per|3007,3010
HPI|3011,3014
<EOL>|3016,3017
(|3017,3018
-|3018,3019
)|3019,3020
Denies|3021,3027
fever|3028,3033
,|3033,3034
chills|3035,3041
,|3041,3042
night|3043,3048
sweats|3049,3055
.|3055,3056
denies|3057,3063
headache|3064,3072
,|3072,3073
sinus|3074,3079
<EOL>|3080,3081
tenderness|3081,3091
,|3091,3092
rhinorrhea|3093,3103
or|3104,3106
congestion|3107,3117
.|3117,3118
Denies|3119,3125
cough|3126,3131
.|3131,3132
Denies|3133,3139
<EOL>|3140,3141
nausea|3141,3147
,|3147,3148
vomiting|3149,3157
,|3157,3158
diarrhea|3159,3167
,|3167,3168
constipation|3169,3181
or|3182,3184
abdominal|3185,3194
pain|3195,3199
.|3199,3200
No|3201,3203
<EOL>|3204,3205
dysuria|3205,3212
.|3212,3213
Denies|3214,3220
arthralgias|3221,3232
or|3233,3235
myalgias|3236,3244
.|3244,3245
<EOL>|3247,3248
<EOL>|3248,3249
<EOL>|3250,3251
Hypertension|3273,3285
<EOL>|3285,3286
Dementia|3286,3294
<EOL>|3294,3295
Osteoporosis|3295,3307
<EOL>|3307,3308
Irritable|3308,3317
bowel|3318,3323
syndrome|3324,3332
<EOL>|3332,3333
Macrocytosis|3333,3345
of|3346,3348
unclear|3349,3356
etiology|3357,3365
<EOL>|3365,3366
Left|3366,3370
ear|3371,3374
hearing|3375,3382
loss|3383,3387
<EOL>|3387,3388
Status|3388,3394
post|3395,3399
hysterectomy|3400,3412
<EOL>|3412,3413
Status|3413,3419
post|3420,3424
appendectomy|3425,3437
<EOL>|3437,3438
Status|3438,3444
post|3445,3449
ovarian|3450,3457
cyst|3458,3462
removal|3463,3470
<EOL>|3470,3471
Cataract|3471,3479
surgery|3480,3487
<EOL>|3487,3488
Glaucoma|3488,3496
<EOL>|3496,3497
<EOL>|3498,3499
:|3513,3514
<EOL>|3514,3515
_|3515,3516
_|3516,3517
_|3517,3518
<EOL>|3518,3519
:|3533,3534
<EOL>|3534,3535
Not|3535,3538
relevant|3539,3547
to|3548,3550
the|3551,3554
current|3555,3562
admission|3563,3572
.|3572,3573
<EOL>|3573,3574
<EOL>|3575,3576
ADMISSION|3591,3600
EXAM|3601,3605
<EOL>|3606,3607
=|3607,3608
=|3608,3609
=|3609,3610
=|3610,3611
=|3611,3612
=|3612,3613
=|3613,3614
=|3614,3615
=|3615,3616
=|3616,3617
=|3617,3618
=|3618,3619
=|3619,3620
=|3620,3621
<EOL>|3621,3622
Vital|3622,3627
Signs|3628,3633
:|3633,3634
98.3|3635,3639
,|3639,3640
107|3641,3644
/|3644,3645
43|3645,3647
,|3647,3648
72|3649,3651
,|3651,3652
16|3653,3655
,|3655,3656
99|3657,3659
2L|3660,3662
NC|3663,3665
<EOL>|3667,3668
General|3668,3675
:|3675,3676
AOx1|3677,3681
,|3681,3682
pleasant|3683,3691
,|3691,3692
smiling|3693,3700
,|3700,3701
at|3702,3704
baseline|3705,3713
per|3714,3717
family|3718,3724
members|3725,3732
<EOL>|3733,3734
at|3734,3736
bedside|3737,3744
<EOL>|3745,3746
_|3746,3747
_|3747,3748
_|3748,3749
:|3749,3750
Sclera|3751,3757
anicteric|3758,3767
,|3767,3768
MMM|3769,3772
,|3772,3773
oropharynx|3774,3784
clear|3785,3790
,|3790,3791
EOMI|3792,3796
,|3796,3797
PERRL|3798,3803
,|3803,3804
<EOL>|3805,3806
neck|3806,3810
supple|3811,3817
,|3817,3818
JVP|3819,3822
not|3823,3826
elevated|3827,3835
,|3835,3836
no|3837,3839
LAD|3840,3843
<EOL>|3845,3846
CV|3846,3848
:|3848,3849
Regular|3850,3857
rate|3858,3862
and|3863,3866
rhythm|3867,3873
,|3873,3874
normal|3875,3881
S1|3882,3884
+|3885,3886
S2|3887,3889
,|3889,3890
soft|3891,3895
_|3896,3897
_|3897,3898
_|3898,3899
systolic|3900,3908
<EOL>|3909,3910
murmur|3910,3916
.|3916,3917
<EOL>|3920,3921
Lungs|3921,3926
:|3926,3927
Moderate|3928,3936
inspiratory|3937,3948
effort|3949,3955
,|3955,3956
decreased|3957,3966
breath|3967,3973
sounds|3974,3980
<EOL>|3981,3982
bilaterally|3982,3993
at|3994,3996
bases|3997,4002
L|4003,4004
>|4004,4005
R.|4005,4007
No|4008,4010
wheezes|4011,4018
,|4018,4019
rales|4020,4025
,|4025,4026
rhonchi|4027,4034
<EOL>|4036,4037
Abdomen|4037,4044
:|4044,4045
Soft|4046,4050
,|4050,4051
non-tender|4052,4062
,|4062,4063
non-distended|4064,4077
,|4077,4078
bowel|4079,4084
sounds|4085,4091
present|4092,4099
,|4099,4100
<EOL>|4101,4102
no|4102,4104
organomegaly|4105,4117
,|4117,4118
no|4119,4121
rebound|4122,4129
or|4130,4132
guarding|4133,4141
<EOL>|4143,4144
GU|4144,4146
:|4146,4147
No|4148,4150
foley|4151,4156
<EOL>|4158,4159
Ext|4159,4162
:|4162,4163
Warm|4164,4168
,|4168,4169
well|4170,4174
perfused|4175,4183
,|4183,4184
2|4185,4186
+|4186,4187
pulses|4188,4194
,|4194,4195
L|4196,4197
>|4197,4198
R|4198,4199
lower|4200,4205
extremity|4206,4215
<EOL>|4216,4217
swelling|4217,4225
with|4226,4230
left|4231,4235
leg|4236,4239
erythematous|4240,4252
and|4253,4256
tender|4257,4263
to|4264,4266
palpation|4267,4276
,|4276,4277
2|4278,4279
+|4279,4280
<EOL>|4281,4282
pitting|4282,4289
edema|4290,4295
tender|4296,4302
,|4302,4303
right|4304,4309
lower|4310,4315
extremity|4316,4325
with|4326,4330
e|4331,4332
/|4332,4333
o|4333,4334
chronic|4335,4342
<EOL>|4343,4344
venous|4344,4350
stasis|4351,4357
changes|4358,4365
,|4365,4366
1|4367,4368
+|4368,4369
pitting|4370,4377
edema|4378,4383
non|4384,4387
tender|4388,4394
.|4394,4395
<EOL>|4397,4398
Neuro|4398,4403
:|4403,4404
AOx1|4405,4409
,|4409,4410
strength|4411,4419
_|4420,4421
_|4421,4422
_|4422,4423
upper|4424,4429
and|4430,4433
lower|4434,4439
exteremities|4440,4452
,|4452,4453
all|4454,4457
<EOL>|4458,4459
facial|4459,4465
movements|4466,4475
in|4476,4478
tact|4479,4483
,|4483,4484
sensation|4485,4494
grossly|4495,4502
in|4503,4505
tact|4506,4510
,|4510,4511
gait|4512,4516
<EOL>|4517,4518
deferred|4518,4526
.|4526,4527
<EOL>|4529,4530
<EOL>|4531,4532
DISCHARGE|4532,4541
EXAM|4542,4546
<EOL>|4547,4548
=|4548,4549
=|4549,4550
=|4550,4551
=|4551,4552
=|4552,4553
=|4553,4554
=|4554,4555
=|4555,4556
=|4556,4557
=|4557,4558
=|4558,4559
=|4559,4560
=|4560,4561
=|4561,4562
<EOL>|4562,4563
Vitals|4563,4569
:|4569,4570
T|4571,4572
:|4572,4573
97.9|4573,4577
,|4577,4578
144|4579,4582
/|4582,4583
59|4583,4585
,|4585,4586
72|4587,4589
,|4589,4590
20|4591,4593
,|4593,4594
93|4595,4597
RA|4598,4600
<EOL>|4601,4602
<EOL>|4602,4603
General|4603,4610
:|4610,4611
AOx1|4612,4616
,|4616,4617
pleasant|4618,4626
,|4626,4627
smiling|4628,4635
,|4635,4636
at|4637,4639
baseline|4640,4648
per|4649,4652
family|4653,4659
members|4660,4667
<EOL>|4668,4669
at|4669,4671
bedside|4672,4679
<EOL>|4680,4681
_|4681,4682
_|4682,4683
_|4683,4684
:|4684,4685
Sclera|4686,4692
anicteric|4693,4702
,|4702,4703
MMM|4704,4707
<EOL>|4709,4710
CV|4710,4712
:|4712,4713
Irregularly|4714,4725
irregular|4726,4735
,|4735,4736
normal|4737,4743
S1|4744,4746
+|4747,4748
S2|4749,4751
,|4751,4752
soft|4753,4757
_|4758,4759
_|4759,4760
_|4760,4761
systolic|4762,4770
<EOL>|4771,4772
murmur|4772,4778
.|4778,4779
<EOL>|4782,4783
Lungs|4783,4788
:|4788,4789
Moderate|4790,4798
inspiratory|4799,4810
effort|4811,4817
,|4817,4818
decreased|4819,4828
breath|4829,4835
sounds|4836,4842
<EOL>|4843,4844
bilateral|4844,4853
bases|4854,4859
<EOL>|4860,4861
Ext|4861,4864
:|4864,4865
Warm|4866,4870
,|4870,4871
well|4872,4876
perfused|4877,4885
,|4885,4886
2|4887,4888
+|4888,4889
pulses|4890,4896
,|4896,4897
L|4898,4899
>|4899,4900
R|4900,4901
lower|4902,4907
extremity|4908,4917
<EOL>|4918,4919
swelling|4919,4927
with|4928,4932
left|4933,4937
leg|4938,4941
erythematous|4942,4954
and|4955,4958
minimal|4959,4966
tender|4967,4973
to|4974,4976
<EOL>|4977,4978
palpation|4978,4987
,|4987,4988
2|4989,4990
+|4990,4991
pitting|4992,4999
edema|5000,5005
tender|5006,5012
,|5012,5013
right|5014,5019
lower|5020,5025
extremity|5026,5035
with|5036,5040
<EOL>|5041,5042
e|5042,5043
/|5043,5044
o|5044,5045
chronic|5046,5053
venous|5054,5060
stasis|5061,5067
changes|5068,5075
,|5075,5076
1|5077,5078
+|5078,5079
pitting|5080,5087
edema|5088,5093
non|5094,5097
tender|5098,5104
.|5104,5105
<EOL>|5107,5108
<EOL>|5108,5109
Neuro|5109,5114
:|5114,5115
AOx1|5116,5120
<EOL>|5122,5123
<EOL>|5123,5124
<EOL>|5125,5126
Pertinent|5126,5135
Results|5136,5143
:|5143,5144
<EOL>|5144,5145
ADMISSION|5145,5154
LABS|5155,5159
<EOL>|5159,5160
=|5160,5161
=|5161,5162
=|5162,5163
=|5163,5164
=|5164,5165
=|5165,5166
=|5166,5167
=|5167,5168
=|5168,5169
=|5169,5170
=|5170,5171
=|5171,5172
=|5172,5173
=|5173,5174
<EOL>|5174,5175
_|5175,5176
_|5176,5177
_|5177,5178
11|5179,5181
:|5181,5182
35AM|5182,5186
URINE|5187,5192
RBC|5194,5197
-|5197,5198
2|5198,5199
WBC|5200,5203
-|5203,5204
22|5204,5206
*|5206,5207
BACTERIA|5208,5216
-|5216,5217
NONE|5217,5221
YEAST|5222,5227
-|5227,5228
NONE|5228,5232
<EOL>|5233,5234
EPI|5234,5237
-|5237,5238
<|5238,5239
1|5239,5240
TRANS|5241,5246
EPI|5247,5250
-|5250,5251
<|5251,5252
1|5252,5253
<EOL>|5253,5254
_|5254,5255
_|5255,5256
_|5256,5257
11|5258,5260
:|5260,5261
35AM|5261,5265
URINE|5266,5271
BLOOD|5273,5278
-|5278,5279
NEG|5279,5282
NITRITE|5283,5290
-|5290,5291
NEG|5291,5294
PROTEIN|5295,5302
-|5302,5303
NEG|5303,5306
<EOL>|5307,5308
GLUCOSE|5308,5315
-|5315,5316
NEG|5316,5319
KETONE|5320,5326
-|5326,5327
NEG|5327,5330
BILIRUBIN|5331,5340
-|5340,5341
NEG|5341,5344
UROBILNGN|5345,5354
-|5354,5355
NEG|5355,5358
PH|5359,5361
-|5361,5362
5.5|5362,5365
<EOL>|5366,5367
LEUK|5367,5371
-|5371,5372
MOD|5372,5375
<EOL>|5375,5376
_|5376,5377
_|5377,5378
_|5378,5379
12|5380,5382
:|5382,5383
00PM|5383,5387
PLT|5390,5393
COUNT|5394,5399
-|5399,5400
168|5400,5403
<EOL>|5403,5404
_|5404,5405
_|5405,5406
_|5406,5407
12|5408,5410
:|5410,5411
00PM|5411,5415
NEUTS|5418,5423
-|5423,5424
81|5424,5426
.|5426,5427
1|5427,5428
*|5428,5429
LYMPHS|5430,5436
-|5436,5437
10|5437,5439
.|5439,5440
8|5440,5441
*|5441,5442
MONOS|5443,5448
-|5448,5449
6.7|5449,5452
EOS|5453,5456
-|5456,5457
0|5457,5458
.|5458,5459
1|5459,5460
*|5460,5461
<EOL>|5462,5463
BASOS|5463,5468
-|5468,5469
0.2|5469,5472
IM|5473,5475
_|5476,5477
_|5477,5478
_|5478,5479
AbsNeut|5480,5487
-|5487,5488
11|5488,5490
.|5490,5491
29|5491,5493
*|5493,5494
AbsLymp|5495,5502
-|5502,5503
1|5503,5504
.|5504,5505
51|5505,5507
AbsMono|5508,5515
-|5515,5516
0|5516,5517
.|5517,5518
94|5518,5520
*|5520,5521
<EOL>|5522,5523
AbsEos|5523,5529
-|5529,5530
0|5530,5531
.|5531,5532
02|5532,5534
*|5534,5535
AbsBaso|5536,5543
-|5543,5544
0|5544,5545
.|5545,5546
03|5546,5548
<EOL>|5548,5549
_|5549,5550
_|5550,5551
_|5551,5552
12|5553,5555
:|5555,5556
00PM|5556,5560
WBC|5563,5566
-|5566,5567
13|5567,5569
.|5569,5570
9|5570,5571
*|5571,5572
RBC|5573,5576
-|5576,5577
3|5577,5578
.|5578,5579
78|5579,5581
*|5581,5582
HGB|5583,5586
-|5586,5587
12.5|5587,5591
HCT|5592,5595
-|5595,5596
39.2|5596,5600
<EOL>|5601,5602
MCV|5602,5605
-|5605,5606
104|5606,5609
*|5609,5610
MCH|5611,5614
-|5614,5615
33|5615,5617
.|5617,5618
1|5618,5619
*|5619,5620
MCHC|5621,5625
-|5625,5626
31|5626,5628
.|5628,5629
9|5629,5630
*|5630,5631
RDW|5632,5635
-|5635,5636
13.6|5636,5640
RDWSD|5641,5646
-|5646,5647
51|5647,5649
.|5649,5650
9|5650,5651
*|5651,5652
<EOL>|5652,5653
_|5653,5654
_|5654,5655
_|5655,5656
12|5657,5659
:|5659,5660
00PM|5660,5664
CALCIUM|5667,5674
-|5674,5675
7|5675,5676
.|5676,5677
8|5677,5678
*|5678,5679
PHOSPHATE|5680,5689
-|5689,5690
3.7|5690,5693
MAGNESIUM|5694,5703
-|5703,5704
1.6|5704,5707
<EOL>|5707,5708
_|5708,5709
_|5709,5710
_|5710,5711
12|5712,5714
:|5714,5715
00PM|5715,5719
cTropnT|5722,5729
-|5729,5730
0|5730,5731
.|5731,5732
03|5732,5734
*|5734,5735
proBNP|5736,5742
-|5742,5743
8428|5743,5747
*|5747,5748
<EOL>|5748,5749
_|5749,5750
_|5750,5751
_|5751,5752
12|5753,5755
:|5755,5756
00PM|5756,5760
GLUCOSE|5763,5770
-|5770,5771
118|5771,5774
*|5774,5775
UREA|5776,5780
N|5781,5782
-|5782,5783
26|5783,5785
*|5785,5786
CREAT|5787,5792
-|5792,5793
0.8|5793,5796
SODIUM|5797,5803
-|5803,5804
144|5804,5807
<EOL>|5808,5809
POTASSIUM|5809,5818
-|5818,5819
2|5819,5820
.|5820,5821
8|5821,5822
*|5822,5823
CHLORIDE|5824,5832
-|5832,5833
95|5833,5835
*|5835,5836
TOTAL|5837,5842
CO2|5843,5846
-|5846,5847
38|5847,5849
*|5849,5850
ANION|5851,5856
GAP|5857,5860
-|5860,5861
14|5861,5863
<EOL>|5863,5864
<EOL>|5864,5865
STUDIES|5865,5872
<EOL>|5872,5873
=|5873,5874
=|5874,5875
=|5875,5876
=|5876,5877
=|5877,5878
=|5878,5879
=|5879,5880
<EOL>|5880,5881
<EOL>|5881,5882
CXR|5882,5885
<EOL>|5886,5887
Bilateral|5887,5896
pleural|5897,5904
effusions|5905,5914
,|5914,5915
large|5916,5921
on|5922,5924
the|5925,5928
right|5929,5934
and|5935,5938
small|5939,5944
on|5945,5947
the|5948,5951
<EOL>|5952,5953
left|5953,5957
.|5957,5958
No|5960,5962
<EOL>|5963,5964
definite|5964,5972
focal|5973,5978
consolidation|5979,5992
identified|5993,6003
,|6003,6004
although|6005,6013
evaluation|6014,6024
is|6025,6027
<EOL>|6028,6029
limited|6029,6036
<EOL>|6037,6038
secondary|6038,6047
to|6048,6050
these|6051,6056
effusions|6057,6066
.|6066,6067
<EOL>|6068,6069
<EOL>|6069,6070
Pelvis|6070,6076
Xray|6077,6081
<EOL>|6082,6083
There|6083,6088
is|6089,6091
no|6092,6094
acute|6095,6100
fracture|6101,6109
or|6110,6112
dislocation|6113,6124
.|6124,6125
No|6127,6129
focal|6130,6135
lytic|6136,6141
or|6142,6144
<EOL>|6145,6146
sclerotic|6146,6155
<EOL>|6156,6157
osseous|6157,6164
lesion|6165,6171
is|6172,6174
seen|6175,6179
.|6179,6180
There|6182,6187
is|6188,6190
no|6191,6193
radiopaque|6194,6204
foreign|6205,6212
body|6213,6217
.|6217,6218
<EOL>|6220,6221
Vascular|6221,6229
<EOL>|6230,6231
calcifications|6231,6245
are|6246,6249
noted|6250,6255
.|6255,6256
The|6258,6261
visualized|6262,6272
bowel|6273,6278
gas|6279,6282
pattern|6283,6290
is|6291,6293
<EOL>|6294,6295
nonobstructive|6295,6309
.|6309,6310
<EOL>|6311,6312
<EOL>|6314,6315
IMPRESSION|6315,6325
:|6325,6326
No|6328,6330
acute|6331,6336
fracture|6337,6345
or|6346,6348
dislocation|6349,6360
.|6360,6361
<EOL>|6362,6363
<EOL>|6363,6364
Lower|6364,6369
extremity|6370,6379
ultrasound|6380,6390
<EOL>|6391,6392
1.|6392,6394
Deep|6395,6399
vein|6400,6404
thrombosis|6405,6415
of|6416,6418
the|6419,6422
left|6423,6427
common|6428,6434
femoral|6435,6442
vein|6443,6447
<EOL>|6448,6449
extending|6449,6458
into|6459,6463
at|6464,6466
<EOL>|6467,6468
least|6468,6473
the|6474,6477
popliteal|6478,6487
vein|6488,6492
.|6492,6493
Left|6495,6499
calf|6500,6504
veins|6505,6510
were|6511,6515
not|6516,6519
clearly|6520,6527
<EOL>|6528,6529
identified|6529,6539
,|6539,6540
<EOL>|6541,6542
possibly|6542,6550
also|6551,6555
occluded|6556,6564
.|6564,6565
<EOL>|6566,6567
2|6567,6568
.|6568,6569
No|6571,6573
right|6574,6579
DVT|6580,6583
.|6583,6584
<EOL>|6585,6586
<EOL>|6586,6587
LAST|6587,6591
LABS|6592,6596
BEFORE|6597,6603
DISCHARGE|6604,6613
<EOL>|6614,6615
=|6615,6616
=|6616,6617
=|6617,6618
=|6618,6619
=|6619,6620
=|6620,6621
=|6621,6622
=|6622,6623
=|6623,6624
=|6624,6625
=|6625,6626
=|6626,6627
=|6627,6628
=|6628,6629
=|6629,6630
=|6630,6631
=|6631,6632
=|6632,6633
=|6633,6634
=|6634,6635
=|6635,6636
=|6636,6637
=|6637,6638
=|6638,6639
=|6639,6640
=|6640,6641
=|6641,6642
=|6642,6643
=|6643,6644
=|6644,6645
=|6645,6646
<EOL>|6646,6647
_|6647,6648
_|6648,6649
_|6649,6650
06|6651,6653
:|6653,6654
55AM|6654,6658
BLOOD|6659,6664
WBC|6665,6668
-|6668,6669
14|6669,6671
.|6671,6672
9|6672,6673
*|6673,6674
RBC|6675,6678
-|6678,6679
3|6679,6680
.|6680,6681
51|6681,6683
*|6683,6684
Hgb|6685,6688
-|6688,6689
11.5|6689,6693
Hct|6694,6697
-|6697,6698
36.8|6698,6702
<EOL>|6703,6704
MCV|6704,6707
-|6707,6708
105|6708,6711
*|6711,6712
MCH|6713,6716
-|6716,6717
32|6717,6719
.|6719,6720
8|6720,6721
*|6721,6722
MCHC|6723,6727
-|6727,6728
31|6728,6730
.|6730,6731
3|6731,6732
*|6732,6733
RDW|6734,6737
-|6737,6738
13.8|6738,6742
RDWSD|6743,6748
-|6748,6749
53|6749,6751
.|6751,6752
1|6752,6753
*|6753,6754
Plt|6755,6758
_|6759,6760
_|6760,6761
_|6761,6762
<EOL>|6762,6763
_|6763,6764
_|6764,6765
_|6765,6766
06|6767,6769
:|6769,6770
55AM|6770,6774
BLOOD|6775,6780
Glucose|6781,6788
-|6788,6789
109|6789,6792
*|6792,6793
UreaN|6794,6799
-|6799,6800
32|6800,6802
*|6802,6803
Creat|6804,6809
-|6809,6810
0.9|6810,6813
Na|6814,6816
-|6816,6817
144|6817,6820
<EOL>|6821,6822
K|6822,6823
-|6823,6824
3.7|6824,6827
Cl|6828,6830
-|6830,6831
96|6831,6833
HCO3|6834,6838
-|6838,6839
37|6839,6841
*|6841,6842
AnGap|6843,6848
-|6848,6849
15|6849,6851
<EOL>|6851,6852
_|6852,6853
_|6853,6854
_|6854,6855
06|6856,6858
:|6858,6859
55AM|6859,6863
BLOOD|6864,6869
Albumin|6870,6877
-|6877,6878
2|6878,6879
.|6879,6880
5|6880,6881
*|6881,6882
Calcium|6883,6890
-|6890,6891
8|6891,6892
.|6892,6893
0|6893,6894
*|6894,6895
Phos|6896,6900
-|6900,6901
3.2|6901,6904
<EOL>|6905,6906
Mg|6906,6908
-|6908,6909
1|6909,6910
.|6910,6911
5|6911,6912
*|6912,6913
<EOL>|6913,6914
<EOL>|6915,6916
_|6939,6940
_|6940,6941
_|6941,6942
is|6943,6945
a|6946,6947
_|6948,6949
_|6949,6950
_|6950,6951
y|6952,6953
/|6953,6954
o|6954,6955
F|6956,6957
with|6958,6962
PMHx|6963,6967
CHF|6968,6971
,|6971,6972
Afib|6973,6977
not|6978,6981
on|6982,6984
<EOL>|6985,6986
anticoagulation|6986,7001
,|7001,7002
severe|7003,7009
advanced|7010,7018
Alzheimer|7019,7028
's|7028,7030
dementia|7031,7039
,|7039,7040
<EOL>|7041,7042
osteoporosis|7042,7054
,|7054,7055
HTN|7056,7059
,|7059,7060
who|7061,7064
presents|7065,7073
from|7074,7078
assisted|7079,7087
living|7088,7094
facility|7095,7103
<EOL>|7104,7105
with|7105,7109
R|7110,7111
hip|7112,7115
pain|7116,7120
,|7120,7121
found|7122,7127
to|7128,7130
have|7131,7135
DVT|7136,7139
left|7140,7144
common|7145,7151
femoral|7152,7159
vein|7160,7164
with|7165,7169
<EOL>|7170,7171
volume|7171,7177
overload|7178,7186
.|7186,7187
During|7188,7194
a|7195,7196
meeting|7197,7204
with|7205,7209
patient|7210,7217
and|7218,7221
her|7222,7225
family|7226,7232
,|7232,7233
<EOL>|7234,7235
decision|7235,7243
was|7244,7247
made|7248,7252
to|7253,7255
transition|7256,7266
care|7267,7271
to|7272,7274
comfort|7275,7282
-|7282,7283
directed|7283,7291
<EOL>|7292,7293
measures|7293,7301
only|7302,7306
and|7307,7310
to|7311,7313
pursue|7314,7320
hospice|7321,7328
services|7329,7337
on|7338,7340
discharge|7341,7350
.|7350,7351
<EOL>|7352,7353
<EOL>|7353,7354
ACTIVE|7354,7360
ISSUES|7361,7367
<EOL>|7368,7369
=|7369,7370
=|7370,7371
=|7371,7372
=|7372,7373
=|7373,7374
=|7374,7375
=|7375,7376
=|7376,7377
=|7377,7378
=|7378,7379
=|7379,7380
=|7380,7381
=|7381,7382
<EOL>|7382,7383
#|7383,7384
CMO|7385,7388
.|7388,7389
The|7390,7393
team|7394,7398
had|7399,7402
a|7403,7404
family|7405,7411
meeting|7412,7419
on|7420,7422
_|7423,7424
_|7424,7425
_|7425,7426
and|7427,7430
decision|7431,7439
was|7440,7443
<EOL>|7444,7445
made|7445,7449
to|7450,7452
transition|7453,7463
care|7464,7468
to|7469,7471
CMO|7472,7475
and|7476,7479
pursue|7480,7486
24|7487,7489
hour|7490,7494
hospice|7495,7502
<EOL>|7503,7504
services|7504,7512
on|7513,7515
discharge|7516,7525
.|7525,7526
Family|7527,7533
did|7534,7537
not|7538,7541
want|7542,7546
to|7547,7549
pursue|7550,7556
active|7557,7563
<EOL>|7564,7565
treatments|7565,7575
such|7576,7580
as|7581,7583
Lasix|7584,7589
,|7589,7590
which|7591,7596
would|7597,7602
make|7603,7607
her|7608,7611
uncomfortable|7612,7625
<EOL>|7626,7627
given|7627,7632
incontinence|7633,7645
or|7646,7648
shots|7649,7654
such|7655,7659
as|7660,7662
lovenox|7663,7670
for|7671,7674
treatment|7675,7684
of|7685,7687
<EOL>|7688,7689
DVT|7689,7692
.|7692,7693
Home|7694,7698
medications|7699,7710
metoprolol|7711,7721
,|7721,7722
donepezil|7723,7732
and|7733,7736
Memantine|7737,7746
were|7747,7751
<EOL>|7752,7753
continued|7753,7762
for|7763,7766
comfort|7767,7774
.|7774,7775
She|7776,7779
was|7780,7783
discharged|7784,7794
to|7795,7797
an|7798,7800
_|7801,7802
_|7802,7803
_|7803,7804
<EOL>|7805,7806
_|7806,7807
_|7807,7808
_|7808,7809
facility|7810,7818
.|7818,7819
<EOL>|7820,7821
<EOL>|7821,7822
OTHER|7822,7827
HOSPITAL|7828,7836
ISSUES|7837,7843
<EOL>|7844,7845
=|7845,7846
=|7846,7847
=|7847,7848
=|7848,7849
=|7849,7850
=|7850,7851
=|7851,7852
=|7852,7853
=|7853,7854
=|7854,7855
=|7855,7856
=|7856,7857
=|7857,7858
=|7858,7859
=|7859,7860
=|7860,7861
=|7861,7862
=|7862,7863
=|7863,7864
=|7864,7865
=|7865,7866
<EOL>|7866,7867
<EOL>|7867,7868
#|7868,7869
DVT|7870,7873
.|7873,7874
Deep|7875,7879
vein|7880,7884
thrombosis|7885,7895
of|7896,7898
the|7899,7902
left|7903,7907
common|7908,7914
femoral|7915,7922
vein|7923,7927
<EOL>|7928,7929
extending|7929,7938
into|7939,7943
at|7944,7946
least|7947,7952
the|7953,7956
popliteal|7957,7966
vein|7967,7971
diagnosed|7972,7981
on|7982,7984
<EOL>|7985,7986
ultrasound|7986,7996
on|7997,7999
admission|8000,8009
.|8009,8010
This|8011,8015
was|8016,8019
likely|8020,8026
acquired|8027,8035
in|8036,8038
the|8039,8042
setting|8043,8050
<EOL>|8051,8052
of|8052,8054
immobility|8055,8065
,|8065,8066
as|8067,8069
the|8070,8073
patient|8074,8081
had|8082,8085
been|8086,8090
restricted|8091,8101
to|8102,8104
her|8105,8108
<EOL>|8109,8110
wheelchair|8110,8120
at|8121,8123
her|8124,8127
assisted|8128,8136
living|8137,8143
for|8144,8147
greater|8148,8155
than|8156,8160
1|8161,8162
month|8163,8168
due|8169,8172
<EOL>|8173,8174
to|8174,8176
deconditioning|8177,8191
.|8191,8192
She|8193,8196
was|8197,8200
initially|8201,8210
started|8211,8218
on|8219,8221
Lovenox|8222,8229
for|8230,8233
<EOL>|8234,8235
treatment|8235,8244
but|8245,8248
this|8249,8253
was|8254,8257
discontinued|8258,8270
in|8271,8273
the|8274,8277
setting|8278,8285
of|8286,8288
transition|8289,8299
<EOL>|8300,8301
to|8301,8303
care|8304,8308
to|8309,8311
CMO|8312,8315
as|8316,8318
above|8319,8324
.|8324,8325
<EOL>|8326,8327
<EOL>|8327,8328
#|8328,8329
Acute|8330,8335
CHF|8336,8339
.|8339,8340
Patient|8341,8348
was|8349,8352
volume|8353,8359
overloaded|8360,8370
on|8371,8373
presentation|8374,8386
with|8387,8391
<EOL>|8392,8393
pleural|8393,8400
effusions|8401,8410
.|8410,8411
She|8412,8415
was|8416,8419
diuresed|8420,8428
with|8429,8433
IV|8434,8436
Lasix|8437,8442
.|8442,8443
Home|8444,8448
<EOL>|8449,8450
metoprolol|8450,8460
was|8461,8464
continued|8465,8474
at|8475,8477
a|8478,8479
decreased|8480,8489
dose|8490,8494
.|8494,8495
In|8496,8498
the|8499,8502
setting|8503,8510
of|8511,8513
<EOL>|8514,8515
transition|8515,8525
to|8526,8528
care|8529,8533
to|8534,8536
CMO|8537,8540
,|8540,8541
Lasix|8542,8547
was|8548,8551
discontinued|8552,8564
.|8564,8565
She|8566,8569
was|8570,8573
<EOL>|8574,8575
continued|8575,8584
on|8585,8587
metoprolol|8588,8598
for|8599,8602
comfort|8603,8610
.|8610,8611
She|8612,8615
remained|8616,8624
on|8625,8627
room|8628,8632
air|8633,8636
<EOL>|8637,8638
without|8638,8645
respiratory|8646,8657
distress|8658,8666
.|8666,8667
<EOL>|8669,8670
<EOL>|8670,8671
#|8671,8672
Afib|8673,8677
.|8677,8678
She|8679,8682
presented|8683,8692
in|8693,8695
sinus|8696,8701
rhythm|8702,8708
,|8708,8709
rate|8710,8714
controlled|8715,8725
on|8726,8728
<EOL>|8729,8730
metoprolol|8730,8740
.|8740,8741
Metoprolol|8742,8752
was|8753,8756
continued|8757,8766
at|8767,8769
a|8770,8771
decreased|8772,8781
dose|8782,8786
for|8787,8790
<EOL>|8791,8792
comfort|8792,8799
.|8799,8800
<EOL>|8801,8802
<EOL>|8802,8803
#|8803,8804
Hip|8805,8808
pain|8809,8813
.|8813,8814
The|8815,8818
right|8819,8824
hip|8825,8828
pain|8829,8833
that|8834,8838
she|8839,8842
presented|8843,8852
with|8853,8857
was|8858,8861
<EOL>|8862,8863
resolved|8863,8871
by|8872,8874
the|8875,8878
time|8879,8883
of|8884,8886
admission|8887,8896
.|8896,8897
Pelvic|8898,8904
xray|8905,8909
was|8910,8913
without|8914,8921
<EOL>|8922,8923
fracture|8923,8931
.|8931,8932
She|8933,8936
was|8937,8940
treated|8941,8948
with|8949,8953
Tylenol|8954,8961
scheduled|8962,8971
for|8972,8975
pain|8976,8980
<EOL>|8981,8982
control|8982,8989
.|8989,8990
<EOL>|8991,8992
<EOL>|8992,8993
#|8993,8994
Al|8995,8997
_|8997,8998
_|8998,8999
_|8999,9000
Dementia|9001,9009
.|9009,9010
She|9011,9014
was|9015,9018
AOx1|9019,9023
at|9024,9026
her|9027,9030
baseline|9031,9039
per|9040,9043
family|9044,9050
<EOL>|9051,9052
members|9052,9059
.|9059,9060
She|9061,9064
was|9065,9068
continued|9069,9078
on|9079,9081
Aricept|9082,9089
/|9089,9090
Namenda|9090,9097
.|9097,9098
<EOL>|9100,9101
<EOL>|9101,9102
TRANSITIONAL|9102,9114
ISSUES|9115,9121
<EOL>|9122,9123
=|9123,9124
=|9124,9125
=|9125,9126
=|9126,9127
=|9127,9128
=|9128,9129
=|9129,9130
=|9130,9131
=|9131,9132
=|9132,9133
=|9133,9134
=|9134,9135
=|9135,9136
=|9136,9137
=|9137,9138
=|9138,9139
=|9139,9140
=|9140,9141
=|9141,9142
<EOL>|9142,9143
<EOL>|9143,9144
-|9144,9145
_|9146,9147
_|9147,9148
_|9148,9149
facility|9150,9158
to|9159,9161
continue|9162,9170
writing|9171,9178
orders|9179,9185
for|9186,9189
<EOL>|9190,9191
pain|9191,9195
/|9195,9196
anxiety|9196,9203
/|9203,9204
secretions|9204,9214
and|9215,9218
other|9219,9224
symptoms|9225,9233
.|9233,9234
<EOL>|9235,9236
-|9236,9237
Continued|9238,9247
metoprolol|9248,9258
succinate|9259,9268
and|9269,9272
Memantine|9273,9282
and|9283,9286
donepezil|9287,9296
on|9297,9299
<EOL>|9300,9301
discharge|9301,9310
for|9311,9314
comfort|9315,9322
.|9322,9323
Continuation|9324,9336
of|9337,9339
these|9340,9345
medications|9346,9357
can|9358,9361
be|9362,9364
<EOL>|9365,9366
further|9366,9373
decided|9374,9381
at|9382,9384
inpatient|9385,9394
hospice|9395,9402
.|9402,9403
<EOL>|9404,9405
-|9405,9406
MOLST|9407,9412
form|9413,9417
:|9417,9418
DNR|9419,9422
/|9422,9423
DNI|9423,9426
,|9426,9427
do|9428,9430
not|9431,9434
re-hospitalize|9435,9449
<EOL>|9450,9451
<EOL>|9451,9452
#|9452,9453
CODE|9454,9458
:|9458,9459
DNR|9460,9463
/|9463,9464
DNI|9464,9467
,|9467,9468
CMO|9469,9472
<EOL>|9473,9474
#|9474,9475
CONTACT|9476,9483
:|9483,9484
HCP|9485,9488
_|9489,9490
_|9490,9491
_|9491,9492
(|9493,9494
daughter|9494,9502
)|9502,9503
_|9504,9505
_|9505,9506
_|9506,9507
Primary|9508,9515
,|9515,9516
<EOL>|9517,9518
secondary|9518,9527
_|9528,9529
_|9529,9530
_|9530,9531
(|9532,9533
son|9533,9536
)|9536,9537
_|9538,9539
_|9539,9540
_|9540,9541
<EOL>|9541,9542
<EOL>|9543,9544
Medications|9544,9555
on|9556,9558
Admission|9559,9568
:|9568,9569
<EOL>|9569,9570
The|9570,9573
Preadmission|9574,9586
Medication|9587,9597
list|9598,9602
is|9603,9605
accurate|9606,9614
and|9615,9618
complete|9619,9627
.|9627,9628
<EOL>|9628,9629
1.|9629,9631
Metoprolol|9632,9642
Succinate|9643,9652
XL|9653,9655
150|9656,9659
mg|9660,9662
PO|9663,9665
BID|9666,9669
<EOL>|9670,9671
2.|9671,9673
Torsemide|9674,9683
40|9684,9686
mg|9687,9689
PO|9690,9692
DAILY|9693,9698
<EOL>|9699,9700
3.|9700,9702
Aspirin|9703,9710
81|9711,9713
mg|9714,9716
PO|9717,9719
DAILY|9720,9725
<EOL>|9726,9727
4.|9727,9729
Donepezil|9730,9739
10|9740,9742
mg|9743,9745
PO|9746,9748
QHS|9749,9752
<EOL>|9753,9754
5.|9754,9756
raloxifene|9757,9767
60|9768,9770
mg|9771,9773
oral|9774,9778
DAILY|9779,9784
<EOL>|9785,9786
6.|9786,9788
Multivitamins|9789,9802
1|9803,9804
TAB|9805,9808
PO|9809,9811
DAILY|9812,9817
<EOL>|9818,9819
7.|9819,9821
Namenda|9822,9829
XR|9830,9832
(|9833,9834
MEMAntine|9834,9843
)|9843,9844
21|9845,9847
mg|9848,9850
oral|9851,9855
DAILY|9856,9861
<EOL>|9862,9863
8.|9863,9865
Ascorbic|9866,9874
Acid|9875,9879
_|9880,9881
_|9881,9882
_|9882,9883
mg|9884,9886
PO|9887,9889
DAILY|9890,9895
<EOL>|9896,9897
9.|9897,9899
Calcium|9900,9907
Carbonate|9908,9917
1500|9918,9922
mg|9923,9925
PO|9926,9928
DAILY|9929,9934
<EOL>|9935,9936
10|9936,9938
.|9938,9939
Vitamin|9940,9947
D|9948,9949
1000|9950,9954
UNIT|9955,9959
PO|9960,9962
DAILY|9963,9968
<EOL>|9969,9970
11.|9970,9973
Fish|9974,9978
Oil|9979,9982
(|9983,9984
Omega|9984,9989
3|9990,9991
)|9991,9992
1000|9993,9997
mg|9998,10000
PO|10001,10003
DAILY|10004,10009
<EOL>|10010,10011
<EOL>|10011,10012
<EOL>|10013,10014
Discharge|10014,10023
Medications|10024,10035
:|10035,10036
<EOL>|10036,10037
1.|10037,10039
Donepezil|10040,10049
10|10050,10052
mg|10053,10055
PO|10056,10058
QHS|10059,10062
<EOL>|10063,10064
2.|10064,10066
Metoprolol|10067,10077
Succinate|10078,10087
XL|10088,10090
200|10091,10094
mg|10095,10097
PO|10098,10100
DAILY|10101,10106
<EOL>|10107,10108
3.|10108,10110
Namenda|10111,10118
XR|10119,10121
(|10122,10123
MEMAntine|10123,10132
)|10132,10133
21|10134,10136
mg|10137,10139
oral|10140,10144
DAILY|10145,10150
<EOL>|10151,10152
4.|10152,10154
Acetaminophen|10155,10168
1000|10169,10173
mg|10174,10176
PO|10177,10179
TID|10180,10183
<EOL>|10184,10185
5.|10185,10187
Glycopyrrolate|10188,10202
0.1|10203,10206
mg|10207,10209
IV|10210,10212
Q6H|10213,10216
:|10216,10217
PRN|10217,10220
excess|10221,10227
secretions|10228,10238
<EOL>|10239,10240
6.|10240,10242
Hyoscyamine|10243,10254
0.125|10255,10260
mg|10261,10263
SL|10264,10266
QID|10267,10270
:|10270,10271
PRN|10271,10274
excess|10275,10281
secretions|10282,10292
<EOL>|10294,10295
<EOL>|10295,10296
<EOL>|10297,10298
Discharge|10298,10307
Disposition|10308,10319
:|10319,10320
<EOL>|10320,10321
Extended|10321,10329
Care|10330,10334
<EOL>|10334,10335
<EOL>|10336,10337
Facility|10337,10345
:|10345,10346
<EOL>|10346,10347
_|10347,10348
_|10348,10349
_|10349,10350
<EOL>|10350,10351
<EOL>|10352,10353
Discharge|10353,10362
Diagnosis|10363,10372
:|10372,10373
<EOL>|10373,10374
-|10394,10395
-|10395,10396
-|10396,10397
-|10397,10398
-|10398,10399
-|10399,10400
-|10400,10401
-|10401,10402
-|10402,10403
-|10403,10404
-|10404,10405
-|10405,10406
-|10406,10407
-|10407,10408
-|10408,10409
<EOL>|10410,10411
Deep|10411,10415
Vein|10416,10420
Thrombosis|10421,10431
<EOL>|10433,10434
<EOL>|10435,10436
Secondary|10436,10445
Diagnosis|10446,10455
<EOL>|10457,10458
-|10458,10459
-|10459,10460
-|10460,10461
-|10461,10462
-|10462,10463
-|10463,10464
-|10464,10465
-|10465,10466
-|10466,10467
-|10467,10468
-|10468,10469
-|10469,10470
-|10470,10471
-|10471,10472
-|10472,10473
-|10473,10474
-|10474,10475
-|10475,10476
<EOL>|10477,10478
Congestive|10478,10488
heart|10489,10494
failure|10495,10502
<EOL>|10503,10504
Atrial|10504,10510
fibrillation|10511,10523
<EOL>|10525,10526
Constipation|10526,10538
<EOL>|10540,10541
Malnutrition|10541,10553
<EOL>|10555,10556
Hypertension|10556,10568
<EOL>|10570,10571
Alzheimer|10571,10580
's|10580,10582
dementia|10583,10591
<EOL>|10593,10594
<EOL>|10594,10595
<EOL>|10596,10597
Mental|10618,10624
Status|10625,10631
:|10631,10632
Confused|10633,10641
-|10642,10643
always|10644,10650
.|10650,10651
<EOL>|10651,10652
Level|10652,10657
of|10658,10660
Consciousness|10661,10674
:|10674,10675
Alert|10676,10681
and|10682,10685
interactive|10686,10697
.|10697,10698
<EOL>|10698,10699
Activity|10699,10707
Status|10708,10714
:|10714,10715
Out|10716,10719
of|10720,10722
Bed|10723,10726
with|10727,10731
assistance|10732,10742
to|10743,10745
chair|10746,10751
or|10752,10754
<EOL>|10755,10756
wheelchair|10756,10766
.|10766,10767
<EOL>|10767,10768
<EOL>|10768,10769
<EOL>|10770,10771
Dear|10795,10799
_|10800,10801
_|10801,10802
_|10802,10803
,|10803,10804
<EOL>|10805,10806
<EOL>|10806,10807
It|10807,10809
was|10810,10813
a|10814,10815
pleasure|10816,10824
taking|10825,10831
care|10832,10836
of|10837,10839
you|10840,10843
during|10844,10850
your|10851,10855
<EOL>|10856,10857
hospitalization|10857,10872
.|10872,10873
Briefly|10874,10881
,|10881,10882
you|10883,10886
were|10887,10891
hospitalized|10892,10904
with|10905,10909
right|10910,10915
hip|10916,10919
<EOL>|10920,10921
pain|10921,10925
.|10925,10926
We|10927,10929
did|10930,10933
Xrays|10934,10939
of|10940,10942
your|10943,10947
hip|10948,10951
which|10952,10957
did|10958,10961
not|10962,10965
show|10966,10970
any|10971,10974
fractures|10975,10984
.|10984,10985
<EOL>|10986,10987
We|10987,10989
also|10990,10994
found|10995,11000
a|11001,11002
blood|11003,11008
clot|11009,11013
in|11014,11016
your|11017,11021
left|11022,11026
leg|11027,11030
and|11031,11034
noticed|11035,11042
that|11043,11047
<EOL>|11048,11049
your|11049,11053
heart|11054,11059
was|11060,11063
n't|11063,11066
pumping|11067,11074
very|11075,11079
efficiently|11080,11091
.|11091,11092
We|11093,11095
talked|11096,11102
with|11103,11107
you|11108,11111
<EOL>|11112,11113
and|11113,11116
your|11117,11121
family|11122,11128
,|11128,11129
who|11130,11133
shared|11134,11140
with|11141,11145
us|11146,11148
many|11149,11153
of|11154,11156
your|11157,11161
wishes|11162,11168
about|11169,11174
<EOL>|11175,11176
being|11176,11181
hospitalized|11182,11194
and|11195,11198
the|11199,11202
type|11203,11207
of|11208,11210
care|11211,11215
you|11216,11219
would|11220,11225
like|11226,11230
to|11231,11233
<EOL>|11234,11235
receive|11235,11242
.|11242,11243
We|11244,11246
decided|11247,11254
to|11255,11257
focus|11258,11263
on|11264,11266
your|11267,11271
comfort|11272,11279
.|11279,11280
Because|11281,11288
of|11289,11291
this|11292,11296
,|11296,11297
<EOL>|11298,11299
you|11299,11302
are|11303,11306
being|11307,11312
discharged|11313,11323
to|11324,11326
_|11327,11328
_|11328,11329
_|11329,11330
for|11331,11334
hospice|11335,11342
care|11343,11347
.|11347,11348
<EOL>|11351,11352
<EOL>|11352,11353
We|11353,11355
wish|11356,11360
you|11361,11364
and|11365,11368
your|11369,11373
family|11374,11380
the|11381,11384
_|11385,11386
_|11386,11387
_|11387,11388
,|11388,11389
<EOL>|11390,11391
<EOL>|11391,11392
Your|11392,11396
_|11397,11398
_|11398,11399
_|11399,11400
Treatment|11401,11410
Team|11411,11415
<EOL>|11416,11417
<EOL>|11418,11419
Followup|11419,11427
Instructions|11428,11440
:|11440,11441
<EOL>|11441,11442
_|11442,11443
_|11443,11444
_|11444,11445
<EOL>|11445,11446

