 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|50,59|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|50,59|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|50,64|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|84,93|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|84,93|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|84,93|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|84,93|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|84,93|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|84,98|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|116,121|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|116,121|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|116,121|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|140,143|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|140,143|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|140,143|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|140,143|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|140,143|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|151,158|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|151,158|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|160,168|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Drug|Organic Chemical|Allergies|183,191|false|false|false|C0086787|Percocet|Percocet
Drug|Pharmacologic Substance|Allergies|183,191|false|false|false|C0086787|Percocet|Percocet
Event|Event|Allergies|194,203|false|false|false|||Attending
Finding|Functional Concept|Allergies|194,203|false|false|false|C1999232|Attending (action)|Attending
Anatomy|Body Location or Region|Chief Complaint|229,238|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|Chief Complaint|229,247|false|false|false|C0235318|Fullness abdominal|abdominal fullness
Event|Event|Chief Complaint|239,247|false|false|false|||fullness
Event|Event|Chief Complaint|252,262|false|false|false|||discomfort
Finding|Sign or Symptom|Chief Complaint|252,262|false|false|false|C2364135|Discomfort|discomfort
Finding|Classification|Chief Complaint|265,270|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|271,279|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|271,279|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|283,301|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|292,301|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|292,301|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|292,301|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|292,301|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|292,301|false|false|false|C0184661|Interventional procedure|Procedure
Drug|Indicator, Reagent, or Diagnostic Aid|Chief Complaint|307,317|false|false|false|C0358514|Diagnostic agents|diagnostic
Event|Event|Chief Complaint|307,317|false|false|false|||diagnostic
Finding|Functional Concept|Chief Complaint|307,317|false|false|false|C0348026;C1547424|Diagnostic;Location Service Code - Diagnostic|diagnostic
Finding|Intellectual Product|Chief Complaint|307,317|false|false|false|C0348026;C1547424|Diagnostic;Location Service Code - Diagnostic|diagnostic
Procedure|Diagnostic Procedure|Chief Complaint|307,317|false|false|false|C0011900;C0430533|Diagnosis;Diagnostic dental procedure|diagnostic
Event|Event|Chief Complaint|318,330|false|false|false|||paracentesis
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|318,330|false|false|false|C0034115|Paracentesis|paracentesis
Drug|Organic Chemical|Chief Complaint|335,346|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Drug|Pharmacologic Substance|Chief Complaint|335,346|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Event|Event|Chief Complaint|335,346|false|false|false|||therapeutic
Finding|Functional Concept|Chief Complaint|335,346|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Finding|Intellectual Product|Chief Complaint|335,346|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|335,346|false|false|false|C0087111|Therapeutic procedure|therapeutic
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|335,359|false|false|false|C2057774|Therapeutic abdominal paracentesis|therapeutic paracentesis
Event|Event|Chief Complaint|347,359|false|false|false|||paracentesis
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|347,359|false|false|false|C0034115|Paracentesis|paracentesis
Disorder|Disease or Syndrome|History of Present Illness|400,403|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Disorder|Virus|History of Present Illness|400,403|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Drug|Immunologic Factor|History of Present Illness|400,403|false|false|false|C0086413|HIV Vaccine|HIV
Drug|Pharmacologic Substance|History of Present Illness|400,403|false|false|false|C0086413|HIV Vaccine|HIV
Event|Event|History of Present Illness|400,403|false|false|false|||HIV
Event|Event|History of Present Illness|407,412|false|false|false|||HAART
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|407,412|false|false|false|C0887947|Antiretroviral Therapy, Highly Active|HAART
Disorder|Disease or Syndrome|History of Present Illness|414,418|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|History of Present Illness|414,418|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|History of Present Illness|414,418|false|false|false|||COPD
Finding|Gene or Genome|History of Present Illness|414,418|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|History of Present Illness|420,423|false|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|HCV
Disorder|Virus|History of Present Illness|420,423|false|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|HCV
Event|Event|History of Present Illness|420,423|false|false|false|||HCV
Disorder|Disease or Syndrome|History of Present Illness|424,433|false|false|false|C0023890;C1623038|Cirrhosis;Liver Cirrhosis|cirrhosis
Event|Event|History of Present Illness|424,433|false|false|false|||cirrhosis
Event|Event|History of Present Illness|434,445|false|false|false|||complicated
Disorder|Disease or Syndrome|History of Present Illness|450,457|false|false|false|C0003962|Ascites|ascites
Event|Event|History of Present Illness|450,457|false|false|false|||ascites
Finding|Pathologic Function|History of Present Illness|450,457|false|false|false|C5441966|Peritoneal Effusion|ascites
Event|Event|History of Present Illness|465,473|false|false|false|||admitted
Anatomy|Body Location or Region|History of Present Illness|479,488|false|false|false|C0000726|Abdomen|abdominal
Finding|Finding|History of Present Illness|479,499|false|false|false|C0000731|Abdomen distended|abdominal distention
Finding|Finding|History of Present Illness|479,508|false|false|false|C2749840|Abdominal distention and pain|abdominal distention and pain
Event|Event|History of Present Illness|489,499|false|false|false|||distention
Finding|Finding|History of Present Illness|489,499|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Finding|Pathologic Function|History of Present Illness|489,499|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Attribute|Clinical Attribute|History of Present Illness|504,508|false|false|false|C2598155||pain
Event|Event|History of Present Illness|504,508|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|504,508|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|504,508|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|519,527|false|false|false|||admitted
Event|Event|History of Present Illness|548,556|false|false|false|||symptoms
Finding|Functional Concept|History of Present Illness|548,556|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|History of Present Illness|548,556|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Drug|Substance|History of Present Illness|578,583|true|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|History of Present Illness|578,583|true|false|false|||fluid
Finding|Intellectual Product|History of Present Illness|578,583|true|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|History of Present Illness|584,591|true|false|false|||removed
Attribute|Clinical Attribute|History of Present Illness|596,599|true|false|false|C0871470|Systolic Pressure|SBP
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|596,599|true|false|false|C0085805|Androgen Binding Protein|SBP
Drug|Biologically Active Substance|History of Present Illness|596,599|true|false|false|C0085805|Androgen Binding Protein|SBP
Event|Event|History of Present Illness|596,599|true|false|false|||SBP
Finding|Gene or Genome|History of Present Illness|596,599|true|false|false|C1705296;C3274833|CCHCR1 wt Allele;SHBG wt Allele|SBP
Procedure|Diagnostic Procedure|History of Present Illness|596,599|true|false|false|C1306620|Systolic blood pressure measurement|SBP
Finding|Gene or Genome|History of Present Illness|612,615|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|History of Present Illness|621,625|false|false|false|||felt
Event|Event|History of Present Illness|626,632|false|false|false|||better
Finding|Idea or Concept|History of Present Illness|626,632|false|false|false|C1550462|Observation Interpretation - better|better
Event|Event|History of Present Illness|640,649|false|false|false|||discharge
Finding|Body Substance|History of Present Illness|640,649|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|History of Present Illness|640,649|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|History of Present Illness|640,649|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|History of Present Illness|640,649|false|false|false|C0030685|Patient Discharge|discharge
Anatomy|Body Location or Region|History of Present Illness|655,662|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|History of Present Illness|655,662|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Event|Event|History of Present Illness|655,662|false|false|false|||abdomen
Finding|Finding|History of Present Illness|655,662|false|false|false|C0941288|Abdomen problem|abdomen
Event|Event|History of Present Illness|667,673|false|false|false|||become
Event|Event|History of Present Illness|688,697|false|false|false|||distended
Finding|Finding|History of Present Illness|688,697|false|false|false|C0700124|Dilated|distended
Attribute|Clinical Attribute|History of Present Illness|703,707|false|false|false|C2598155||pain
Event|Event|History of Present Illness|703,707|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|703,707|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|703,707|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|714,719|false|false|false|||feels
Event|Event|History of Present Illness|720,727|false|false|false|||similar
Event|Event|History of Present Illness|738,746|false|false|false|||episodes
Disorder|Disease or Syndrome|History of Present Illness|750,757|false|false|false|C0003962|Ascites|ascites
Event|Event|History of Present Illness|750,757|false|false|false|||ascites
Finding|Pathologic Function|History of Present Illness|750,757|false|false|false|C5441966|Peritoneal Effusion|ascites
Drug|Pharmacologic Substance|History of Present Illness|765,774|false|false|false|C0012798|Diuretics|diuretics
Event|Event|History of Present Illness|765,774|false|false|false|||diuretics
Event|Event|History of Present Illness|789,798|false|false|false|||decreased
Event|Event|History of Present Illness|813,822|false|false|false|||worsening
Finding|Idea or Concept|History of Present Illness|813,822|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Disorder|Disease or Syndrome|History of Present Illness|824,836|false|false|false|C0020625|Hyponatremia|hyponatremia
Event|Event|History of Present Illness|824,836|false|false|false|||hyponatremia
Event|Event|History of Present Illness|845,857|false|false|false|||hyperkalemia
Finding|Finding|History of Present Illness|845,857|false|false|false|C0020461;C5700154|Hyperkalemia;Serum potassium level above reference range|hyperkalemia
Finding|Body Substance|History of Present Illness|863,870|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|863,870|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|863,870|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|History of Present Illness|871,877|false|false|false|||states
Event|Event|History of Present Illness|892,901|false|false|false|||compliant
Finding|Individual Behavior|History of Present Illness|892,901|false|false|false|C1321605|Compliance behavior|compliant
Disorder|Disease or Syndrome|History of Present Illness|911,914|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Disorder|Virus|History of Present Illness|911,914|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Drug|Immunologic Factor|History of Present Illness|911,914|false|false|false|C0086413|HIV Vaccine|HIV
Drug|Pharmacologic Substance|History of Present Illness|911,914|false|false|false|C0086413|HIV Vaccine|HIV
Event|Event|History of Present Illness|911,914|false|false|false|||HIV
Drug|Pharmacologic Substance|History of Present Illness|919,927|false|false|false|C0012798;C5399719|Diuretic [APC];Diuretics|diuretic
Attribute|Clinical Attribute|History of Present Illness|928,939|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|History of Present Illness|928,939|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|History of Present Illness|928,939|false|false|false|||medications
Finding|Intellectual Product|History of Present Illness|928,939|false|false|false|C4284232|Medications|medications
Event|Event|History of Present Illness|951,957|true|false|false|||filled
Drug|Organic Chemical|History of Present Illness|966,975|true|false|false|C0022957|lactulose|lactulose
Drug|Pharmacologic Substance|History of Present Illness|966,975|true|false|false|C0022957|lactulose|lactulose
Attribute|Clinical Attribute|History of Present Illness|976,988|true|false|false|C5886759|Prescription (attribute)|prescription
Event|Event|History of Present Illness|976,988|true|false|false|||prescription
Finding|Intellectual Product|History of Present Illness|976,988|true|false|false|C1521941|prescription document|prescription
Procedure|Health Care Activity|History of Present Illness|976,988|true|false|false|C0033080|Prescription (procedure)|prescription
Event|Event|History of Present Illness|994,1000|false|false|false|||states
Disorder|Disease or Syndrome|History of Present Illness|1018,1021|false|false|false|C0006430|Burning Mouth Syndrome|BMs
Event|Event|History of Present Illness|1018,1021|false|false|false|||BMs
Finding|Finding|History of Present Illness|1028,1035|false|false|false|C4534363|At home|at home
Event|Event|History of Present Illness|1031,1035|false|false|false|||home
Finding|Idea or Concept|History of Present Illness|1031,1035|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|History of Present Illness|1031,1035|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|History of Present Illness|1031,1035|false|false|false|C1553498|home health encounter|home
Finding|Functional Concept|History of Present Illness|1054,1060|false|false|false|C0234621|Visual|visual
Finding|Sign or Symptom|History of Present Illness|1054,1075|false|false|false|C0233763|Hallucinations, Visual|visual hallucinations
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|1061,1075|false|false|false|C0018524|Hallucinations|hallucinations
Event|Event|History of Present Illness|1061,1075|false|false|false|||hallucinations
Event|Event|History of Present Illness|1081,1094|false|false|false|||forgetfulness
Finding|Sign or Symptom|History of Present Illness|1081,1094|false|false|false|C0542476|Forgetful|forgetfulness
Event|Event|History of Present Illness|1100,1108|false|false|false|||appetite
Finding|Organism Function|History of Present Illness|1100,1108|false|false|false|C0003618|Desire for food|appetite
Event|Event|History of Present Illness|1118,1122|false|false|false|||poor
Finding|Intellectual Product|History of Present Illness|1118,1122|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Finding|Idea or Concept|History of Present Illness|1137,1144|false|false|false|C1555582|Initial (abbreviation)|initial
Event|Event|History of Present Illness|1145,1151|false|false|false|||vitals
Anatomy|Cell Component|History of Present Illness|1183,1186|false|false|false|C2263086|Nuclear cap binding complex location|CBC
Procedure|Laboratory Procedure|History of Present Illness|1183,1186|false|false|false|C0009555|Complete Blood Count|CBC
Drug|Biomedical or Dental Material|History of Present Illness|1193,1201|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|History of Present Illness|1193,1201|false|false|false|||baseline
Finding|Idea or Concept|History of Present Illness|1193,1201|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Attribute|Clinical Attribute|History of Present Illness|1203,1206|false|false|false|C0368980|Coagulation tissue factor induced.INR|INR
Event|Event|History of Present Illness|1203,1206|false|false|false|||INR
Procedure|Laboratory Procedure|History of Present Illness|1203,1206|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1203,1206|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Anatomy|Body Space or Junction|History of Present Illness|1228,1231|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|History of Present Illness|1228,1231|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1228,1231|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|History of Present Illness|1228,1231|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|History of Present Illness|1228,1231|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|History of Present Illness|1228,1231|false|false|false|||AST
Finding|Gene or Genome|History of Present Illness|1228,1231|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Disorder|Neoplastic Process|History of Present Illness|1236,1239|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1236,1239|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|History of Present Illness|1236,1239|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|History of Present Illness|1236,1239|false|false|false|||ALT
Finding|Gene or Genome|History of Present Illness|1236,1239|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|History of Present Illness|1236,1239|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|History of Present Illness|1236,1239|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1236,1239|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Finding|Idea or Concept|History of Present Illness|1247,1252|false|false|false|C1552828|Table Frame - above|above
Drug|Biomedical or Dental Material|History of Present Illness|1254,1262|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|History of Present Illness|1254,1262|false|false|false|||baseline
Finding|Idea or Concept|History of Present Illness|1254,1262|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1279,1286|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Drug|Biologically Active Substance|History of Present Illness|1279,1286|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Drug|Pharmacologic Substance|History of Present Illness|1279,1286|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Event|Event|History of Present Illness|1279,1286|false|false|false|||albumin
Finding|Gene or Genome|History of Present Illness|1279,1286|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|albumin
Finding|Physiologic Function|History of Present Illness|1279,1286|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|albumin
Procedure|Laboratory Procedure|History of Present Illness|1279,1286|false|false|false|C0201838|Albumin measurement|albumin
Drug|Indicator, Reagent, or Diagnostic Aid|History of Present Illness|1292,1302|false|false|false|C0358514|Diagnostic agents|Diagnostic
Event|Event|History of Present Illness|1292,1302|false|false|false|||Diagnostic
Finding|Functional Concept|History of Present Illness|1292,1302|false|false|false|C0348026;C1547424|Diagnostic;Location Service Code - Diagnostic|Diagnostic
Finding|Intellectual Product|History of Present Illness|1292,1302|false|false|false|C0348026;C1547424|Diagnostic;Location Service Code - Diagnostic|Diagnostic
Procedure|Diagnostic Procedure|History of Present Illness|1292,1302|false|false|false|C0011900;C0430533|Diagnosis;Diagnostic dental procedure|Diagnostic
Event|Event|History of Present Illness|1303,1307|false|false|false|||para
Finding|Finding|History of Present Illness|1303,1307|false|false|false|C0030563|Parity|para
Anatomy|Cell|History of Present Illness|1318,1321|false|false|false|C0023516|Leukocytes|WBC
Event|Event|History of Present Illness|1326,1329|false|false|false|||PMN
Finding|Cell Function|History of Present Illness|1326,1329|false|false|false|C2612881;C2825189|Premarket Device Notification;piecemeal microautophagy of the nucleus|PMN
Finding|Intellectual Product|History of Present Illness|1326,1329|false|false|false|C2612881;C2825189|Premarket Device Notification;piecemeal microautophagy of the nucleus|PMN
Finding|Physiologic Function|History of Present Illness|1331,1344|false|false|false|C4553020|Total protein metabolic function|total protein
Lab|Laboratory or Test Result|History of Present Illness|1331,1344|false|false|false|C1261360|Total protein result|total protein
Procedure|Laboratory Procedure|History of Present Illness|1331,1344|false|false|false|C0555903|Total protein measurement|total protein
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1337,1344|false|false|false|C0033684|Proteins|protein
Drug|Biologically Active Substance|History of Present Illness|1337,1344|false|false|false|C0033684|Proteins|protein
Event|Event|History of Present Illness|1337,1344|false|false|false|||protein
Finding|Conceptual Entity|History of Present Illness|1337,1344|false|false|false|C1521746|Protein Info|protein
Procedure|Laboratory Procedure|History of Present Illness|1337,1344|false|false|false|C0202202|Protein measurement|protein
Event|Event|History of Present Illness|1350,1352|false|false|false|||UA
Anatomy|Cell|History of Present Illness|1370,1373|false|false|false|C0023516|Leukocytes|WBC
Disorder|Disease or Syndrome|History of Present Illness|1375,1378|false|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|mod
Finding|Finding|History of Present Illness|1386,1389|false|false|false|C5848551|Neg - answer|neg
Event|Event|History of Present Illness|1400,1412|false|false|false|||contaminated
Finding|Finding|History of Present Illness|1400,1412|false|false|false|C0205279;C1548222;C1548791;C2349974|Bed Status - Contaminated;Contaminated;Contamination;Specimen Condition - Contaminated|contaminated
Finding|Functional Concept|History of Present Illness|1400,1412|false|false|false|C0205279;C1548222;C1548791;C2349974|Bed Status - Contaminated;Contaminated;Contamination;Specimen Condition - Contaminated|contaminated
Finding|Idea or Concept|History of Present Illness|1400,1412|false|false|false|C0205279;C1548222;C1548791;C2349974|Bed Status - Contaminated;Contaminated;Contamination;Specimen Condition - Contaminated|contaminated
Disorder|Disease or Syndrome|History of Present Illness|1420,1423|false|false|false|C0267963|Exocrine pancreatic insufficiency|epi
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1420,1423|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|epi
Drug|Biologically Active Substance|History of Present Illness|1420,1423|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|epi
Drug|Hormone|History of Present Illness|1420,1423|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|epi
Drug|Organic Chemical|History of Present Illness|1420,1423|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|epi
Drug|Pharmacologic Substance|History of Present Illness|1420,1423|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|epi
Event|Event|History of Present Illness|1420,1423|false|false|false|||epi
Finding|Gene or Genome|History of Present Illness|1420,1423|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|epi
Finding|Intellectual Product|History of Present Illness|1420,1423|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|epi
Procedure|Diagnostic Procedure|History of Present Illness|1420,1423|false|false|false|C0162734;C3641909|Echo-Planar Imaging;Electronic Portal Imaging|epi
Event|Event|History of Present Illness|1425,1428|false|false|false|||CXR
Procedure|Diagnostic Procedure|History of Present Illness|1425,1428|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|History of Present Illness|1429,1434|false|false|false|||clear
Finding|Idea or Concept|History of Present Illness|1429,1434|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Location or Region|History of Present Illness|1436,1439|true|false|false|C0230177|Structure of right upper quadrant of abdomen|RUQ
Event|Event|History of Present Illness|1455,1463|true|false|false|||thrombus
Finding|Pathologic Function|History of Present Illness|1455,1463|true|false|false|C0087086;C0302148|Blood Clot;Thrombus|thrombus
Finding|Finding|History of Present Illness|1465,1473|true|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|History of Present Illness|1465,1473|true|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Disorder|Disease or Syndrome|History of Present Illness|1474,1481|true|false|false|C0003962|Ascites|ascites
Event|Event|History of Present Illness|1474,1481|true|false|false|||ascites
Finding|Pathologic Function|History of Present Illness|1474,1481|true|false|false|C5441966|Peritoneal Effusion|ascites
Drug|Organic Chemical|History of Present Illness|1497,1508|false|false|false|C0061851|ondansetron|ondansetron
Drug|Pharmacologic Substance|History of Present Illness|1497,1508|false|false|false|C0061851|ondansetron|ondansetron
Event|Event|History of Present Illness|1497,1508|false|false|false|||ondansetron
Drug|Organic Chemical|History of Present Illness|1521,1529|false|false|false|C0026549|morphine|morphine
Drug|Pharmacologic Substance|History of Present Illness|1521,1529|false|false|false|C0026549|morphine|morphine
Event|Event|History of Present Illness|1521,1529|false|false|false|||morphine
Anatomy|Anatomical Structure|History of Present Illness|1562,1567|false|false|false|C3714591|Floor (anatomic)|floor
Event|Event|History of Present Illness|1576,1583|false|false|false|||feeling
Event|Event|History of Present Illness|1584,1592|false|false|false|||improved
Finding|Finding|History of Present Illness|1584,1592|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Finding|Intellectual Product|History of Present Illness|1584,1592|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Disorder|Disease or Syndrome|History of Present Illness|1597,1602|false|false|false|C1410088|Still|still
Anatomy|Body Location or Region|History of Present Illness|1607,1616|false|false|false|C0000726|Abdomen|abdominal
Event|Event|History of Present Illness|1618,1628|false|false|false|||distention
Finding|Finding|History of Present Illness|1618,1628|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Finding|Pathologic Function|History of Present Illness|1618,1628|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Event|Event|History of Present Illness|1633,1643|false|false|false|||discomfort
Finding|Sign or Symptom|History of Present Illness|1633,1643|false|false|false|C2364135|Discomfort|discomfort
Anatomy|Body Space or Junction|History of Present Illness|1647,1650|false|false|false|C0262327|rostral sulcus|ROS
Drug|Biologically Active Substance|History of Present Illness|1647,1650|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Element, Ion, or Isotope|History of Present Illness|1647,1650|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Organic Chemical|History of Present Illness|1647,1650|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Pharmacologic Substance|History of Present Illness|1647,1650|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Event|Event|History of Present Illness|1647,1650|false|false|false|||ROS
Finding|Gene or Genome|History of Present Illness|1647,1650|false|false|false|C0812281;C1709820|ROS1 gene;ROS1 wt Allele|ROS
Procedure|Health Care Activity|History of Present Illness|1647,1650|false|false|false|C0489633|Review of systems (procedure)|ROS
Anatomy|Body Location or Region|History of Present Illness|1653,1662|false|false|false|C0000726|Abdomen|Abdominal
Finding|Finding|History of Present Illness|1653,1673|false|false|false|C0000731|Abdomen distended|Abdominal distention
Finding|Finding|History of Present Illness|1653,1682|false|false|false|C2749840|Abdominal distention and pain|Abdominal distention and pain
Event|Event|History of Present Illness|1663,1673|false|false|false|||distention
Finding|Finding|History of Present Illness|1663,1673|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Finding|Pathologic Function|History of Present Illness|1663,1673|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Attribute|Clinical Attribute|History of Present Illness|1678,1682|false|false|false|C2598155||pain
Event|Event|History of Present Illness|1678,1682|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|1678,1682|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1678,1682|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|History of Present Illness|1693,1699|true|false|false|C4554530|Bloody|bloody
Finding|Sign or Symptom|History of Present Illness|1693,1706|true|false|false|C1321898|Blood in stool|bloody stools
Attribute|Clinical Attribute|History of Present Illness|1700,1706|true|false|false|C0489144||stools
Event|Event|History of Present Illness|1700,1706|true|false|false|||stools
Finding|Body Substance|History of Present Illness|1700,1706|true|false|false|C0015733|Feces|stools
Attribute|Clinical Attribute|History of Present Illness|1716,1720|true|false|false|C2598155||pain
Event|Event|History of Present Illness|1716,1720|true|false|false|||pain
Finding|Functional Concept|History of Present Illness|1716,1720|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1716,1720|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|1724,1732|true|false|false|||swelling
Finding|Finding|History of Present Illness|1724,1732|true|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|History of Present Illness|1724,1732|true|false|false|C0013604;C0038999|Edema;Swelling|swelling
Event|Event|History of Present Illness|1737,1743|true|false|false|||fevers
Finding|Sign or Symptom|History of Present Illness|1737,1743|true|false|false|C0015967|Fever|fevers
Event|Event|History of Present Illness|1747,1753|true|false|false|||chills
Finding|Sign or Symptom|History of Present Illness|1747,1753|true|false|false|C0085593|Chills|chills
Event|Event|History of Present Illness|1755,1761|false|false|false|||Denies
Anatomy|Body Location or Region|History of Present Illness|1762,1767|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|1762,1767|true|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|1762,1772|true|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|1762,1772|true|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|1768,1772|true|false|false|C2598155||pain
Event|Event|History of Present Illness|1768,1772|true|false|false|||pain
Finding|Functional Concept|History of Present Illness|1768,1772|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1768,1772|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|History of Present Illness|1775,1781|true|false|false|C4255480||nausea
Event|Event|History of Present Illness|1775,1781|true|false|false|||nausea
Finding|Sign or Symptom|History of Present Illness|1775,1781|true|false|false|C0027497|Nausea|nausea
Event|Event|History of Present Illness|1783,1791|true|false|false|||vomiting
Finding|Sign or Symptom|History of Present Illness|1783,1791|true|false|false|C0042963|Vomiting|vomiting
Event|Event|History of Present Illness|1796,1803|true|false|false|||dysuria
Finding|Sign or Symptom|History of Present Illness|1796,1803|true|false|false|C0013428|Dysuria|dysuria
Event|Event|History of Present Illness|1807,1816|true|false|false|||frequency
Finding|Intellectual Product|History of Present Illness|1807,1816|true|false|false|C3898838;C4321352|Frequency;How Often|frequency
Disorder|Disease or Syndrome|Past Medical History|1846,1849|true|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|HCV
Disorder|Virus|Past Medical History|1846,1849|true|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|HCV
Event|Event|Past Medical History|1846,1849|true|false|false|||HCV
Disorder|Disease or Syndrome|Past Medical History|1850,1859|true|false|false|C0023890;C1623038|Cirrhosis;Liver Cirrhosis|Cirrhosis
Event|Event|Past Medical History|1850,1859|true|false|false|||Cirrhosis
Event|Event|Past Medical History|1868,1875|true|false|false|||history
Finding|Conceptual Entity|Past Medical History|1868,1875|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Past Medical History|1868,1875|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Past Medical History|1868,1875|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Past Medical History|1868,1878|true|false|false|C0262926|Medical History|history of
Finding|Finding|Past Medical History|1879,1887|true|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Finding|Idea or Concept|Past Medical History|1879,1887|true|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Finding|Finding|Past Medical History|1879,1898|true|false|false|C0476427|Abnormal cervical smear|abnormal Pap smears
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1888,1891|true|false|false|C3496568|pars anterior of the paramedian lobule|Pap
Drug|Amino Acid, Peptide, or Protein|Past Medical History|1888,1891|true|false|false|C0760170;C1740167|ACPP protein, human;alpha 2-plasmin inhibitor-plasmin complex|Pap
Drug|Enzyme|Past Medical History|1888,1891|true|false|false|C0760170;C1740167|ACPP protein, human;alpha 2-plasmin inhibitor-plasmin complex|Pap
Drug|Immunologic Factor|Past Medical History|1888,1891|true|false|false|C0760170;C1740167|ACPP protein, human;alpha 2-plasmin inhibitor-plasmin complex|Pap
Finding|Finding|Past Medical History|1888,1891|true|false|false|C0428642;C1367456;C1413944;C1413945;C1418410;C1422804;C1423108;C1424700;C1538823;C1705529;C1705530;C1705531;C1863340;C2266415;C3538851;C3889402|ACP3 gene;ACP3 wt Allele;ASAP1 gene;ASAP1 wt Allele;ASAP2 gene;MRPS30 gene;PAPOLA gene;PAPOLA wt Allele;PDAP1 gene;PITUITARY ADENOMA PREDISPOSITION;Pulmonary artery pressure;REG3A gene;REG3A wt Allele;TUSC2 gene;TUSC2 wt Allele|Pap
Finding|Gene or Genome|Past Medical History|1888,1891|true|false|false|C0428642;C1367456;C1413944;C1413945;C1418410;C1422804;C1423108;C1424700;C1538823;C1705529;C1705530;C1705531;C1863340;C2266415;C3538851;C3889402|ACP3 gene;ACP3 wt Allele;ASAP1 gene;ASAP1 wt Allele;ASAP2 gene;MRPS30 gene;PAPOLA gene;PAPOLA wt Allele;PDAP1 gene;PITUITARY ADENOMA PREDISPOSITION;Pulmonary artery pressure;REG3A gene;REG3A wt Allele;TUSC2 gene;TUSC2 wt Allele|Pap
Finding|Molecular Function|Past Medical History|1888,1891|true|false|false|C0428642;C1367456;C1413944;C1413945;C1418410;C1422804;C1423108;C1424700;C1538823;C1705529;C1705530;C1705531;C1863340;C2266415;C3538851;C3889402|ACP3 gene;ACP3 wt Allele;ASAP1 gene;ASAP1 wt Allele;ASAP2 gene;MRPS30 gene;PAPOLA gene;PAPOLA wt Allele;PDAP1 gene;PITUITARY ADENOMA PREDISPOSITION;Pulmonary artery pressure;REG3A gene;REG3A wt Allele;TUSC2 gene;TUSC2 wt Allele|Pap
Procedure|Laboratory Procedure|Past Medical History|1888,1898|true|false|false|C0079104|Pap smear|Pap smears
Event|Event|Past Medical History|1892,1898|true|false|false|||smears
Procedure|Diagnostic Procedure|Past Medical History|1892,1898|true|false|false|C0444186|Smear test|smears
Event|Event|Past Medical History|1913,1926|false|false|false|||calcification
Finding|Organ or Tissue Function|Past Medical History|1913,1926|false|false|false|C0006660;C0006663;C1533591|Calcification;Calcinosis;Physiologic calcification|calcification
Finding|Pathologic Function|Past Medical History|1913,1926|false|false|false|C0006660;C0006663;C1533591|Calcification;Calcinosis;Physiologic calcification|calcification
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1934,1940|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|Past Medical History|1934,1940|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Event|Event|Past Medical History|1934,1940|false|false|false|||breast
Finding|Finding|Past Medical History|1934,1940|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1934,1940|false|false|false|C0191838|Procedures on breast|breast
Event|Event|Past Medical History|1952,1959|true|false|false|||removed
Finding|Body Substance|Past Medical History|1981,1988|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Past Medical History|1981,1988|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Past Medical History|1981,1988|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Past Medical History|2001,2007|true|false|false|||benign
Disorder|Disease or Syndrome|Past Medical History|2018,2021|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Disorder|Virus|Past Medical History|2018,2021|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Drug|Immunologic Factor|Past Medical History|2018,2021|false|false|false|C0086413|HIV Vaccine|HIV
Drug|Pharmacologic Substance|Past Medical History|2018,2021|false|false|false|C0086413|HIV Vaccine|HIV
Disorder|Disease or Syndrome|Past Medical History|2018,2029|false|false|false|C0019693|HIV Infections|HIV disease
Disorder|Disease or Syndrome|Past Medical History|2022,2029|false|false|false|C0012634|Disease|disease
Event|Event|Past Medical History|2022,2029|false|false|false|||disease
Event|Event|Past Medical History|2044,2052|false|false|false|||followed
Disorder|Disease or Syndrome|Past Medical History|2080,2084|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Past Medical History|2080,2084|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Past Medical History|2080,2084|false|false|false|||COPD
Finding|Gene or Genome|Past Medical History|2080,2084|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Finding|Past Medical History|2090,2102|false|false|false|C0332119|Past history of|Past history
Finding|Finding|Past Medical History|2090,2105|false|false|false|C0332119|Past history of|Past history of
Event|Event|Past Medical History|2095,2102|false|false|false|||history
Finding|Conceptual Entity|Past Medical History|2095,2102|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Past Medical History|2095,2102|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Past Medical History|2095,2102|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Past Medical History|2095,2105|false|false|false|C0262926|Medical History|history of
Event|Event|Past Medical History|2106,2113|false|false|false|||smoking
Finding|Individual Behavior|Past Medical History|2106,2113|false|false|false|C0037369;C0453996;C1548578|Location characteristic ID - Smoking;Smoking;Tobacco smoking behavior|smoking
Finding|Intellectual Product|Past Medical History|2106,2113|false|false|false|C0037369;C0453996;C1548578|Location characteristic ID - Smoking;Smoking;Tobacco smoking behavior|smoking
Anatomy|Body System|Past Medical History|2135,2139|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|Past Medical History|2135,2139|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|Past Medical History|2135,2139|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Finding|Body Substance|Past Medical History|2135,2139|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|Past Medical History|2135,2139|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Disorder|Disease or Syndrome|Past Medical History|2135,2146|false|false|false|C0037284|Skin lesion|skin lesion
Event|Event|Past Medical History|2140,2146|false|false|false|||lesion
Finding|Finding|Past Medical History|2140,2146|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|Past Medical History|2140,2146|false|false|false|C0221198;C1546698|Lesion|lesion
Event|Event|Past Medical History|2158,2166|false|false|false|||biopsied
Event|Event|Past Medical History|2171,2177|false|false|false|||showed
Anatomy|Body System|Past Medical History|2180,2184|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|Past Medical History|2180,2184|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|Past Medical History|2180,2184|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Finding|Body Substance|Past Medical History|2180,2184|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|Past Medical History|2180,2184|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Disorder|Neoplastic Process|Past Medical History|2180,2191|false|false|false|C0007114|Malignant neoplasm of skin|skin cancer
Disorder|Neoplastic Process|Past Medical History|2185,2191|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Past Medical History|2185,2191|false|false|false|||cancer
Finding|Body Substance|Past Medical History|2196,2203|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Past Medical History|2196,2203|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Past Medical History|2196,2203|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Past Medical History|2196,2210|false|false|false|C0747307|Patient-Reported|patient report
Attribute|Clinical Attribute|Past Medical History|2204,2210|false|false|false|C4255046||report
Event|Event|Past Medical History|2204,2210|false|false|false|||report
Finding|Intellectual Product|Past Medical History|2204,2210|false|false|false|C0684224|Report (document)|report
Procedure|Health Care Activity|Past Medical History|2204,2210|false|false|false|C0700287|Reporting|report
Event|Event|Past Medical History|2218,2227|false|false|false|||scheduled
Drug|Organic Chemical|Past Medical History|2234,2242|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Past Medical History|2234,2242|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Past Medical History|2234,2242|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|Past Medical History|2234,2242|false|false|false|||complete
Finding|Functional Concept|Past Medical History|2234,2242|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Past Medical History|2234,2242|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Event|Activity|Past Medical History|2245,2252|false|false|false|C1883720|Removing (action)|removal
Event|Event|Past Medical History|2245,2252|false|false|false|||removal
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2245,2252|false|false|false|C0015252;C0185115;C0728940|Excision;Extraction;removal technique|removal
Anatomy|Body System|Past Medical History|2260,2264|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|Past Medical History|2260,2264|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|Past Medical History|2260,2264|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Finding|Body Substance|Past Medical History|2260,2264|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|Past Medical History|2260,2264|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Disorder|Disease or Syndrome|Past Medical History|2260,2271|false|false|false|C0037284|Skin lesion|skin lesion
Event|Event|Past Medical History|2265,2271|false|false|false|||lesion
Finding|Finding|Past Medical History|2265,2271|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|Past Medical History|2265,2271|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Idea or Concept|Past Medical History|2287,2291|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|Past Medical History|2287,2291|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|Past Medical History|2319,2325|false|false|false|||lesion
Finding|Finding|Past Medical History|2319,2325|false|true|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|Past Medical History|2319,2325|false|true|false|C0221198;C1546698|Lesion|lesion
Anatomy|Body Location or Region|Past Medical History|2333,2341|false|false|false|C0016540|Forehead|forehead
Event|Event|Past Medical History|2356,2369|false|false|false|||discoloration
Finding|Finding|Past Medical History|2356,2369|false|false|false|C0332572|Abnormal color|discoloration
Event|Event|Past Medical History|2378,2386|true|false|false|||biopsied
Event|Event|Past Medical History|2390,2397|false|false|false|||exclude
Disorder|Neoplastic Process|Past Medical History|2425,2432|false|false|false|C1261473;C4551686|Malignant neoplasm of soft tissue;Sarcoma|sarcoma
Event|Event|Past Medical History|2425,2432|false|false|false|||sarcoma
Event|Event|Past Medical History|2438,2445|false|false|false|||results
Event|Event|Past Medical History|2449,2456|false|false|false|||pending
Finding|Idea or Concept|Past Medical History|2449,2456|false|false|false|C1691786;C1704475|Pending - Allergy Clinical Status;Pending - referral status|pending
Finding|Finding|Past Medical History|2471,2481|false|false|false|C5961011|Hypoechoic|hypoechoic
Event|Event|Past Medical History|2482,2488|false|false|false|||lesion
Finding|Finding|Past Medical History|2482,2488|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|Past Medical History|2482,2488|false|false|false|C0221198;C1546698|Lesion|lesion
Event|Event|Past Medical History|2496,2506|false|false|false|||ultrasound
Finding|Functional Concept|Past Medical History|2496,2506|false|false|false|C0220934|Ultrasonic|ultrasound
Phenomenon|Natural Phenomenon or Process|Past Medical History|2496,2506|false|false|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|ultrasound
Procedure|Diagnostic Procedure|Past Medical History|2496,2506|false|false|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|ultrasound
Event|Event|Past Medical History|2529,2538|false|false|false|||monitored
Event|Event|Past Medical History|2545,2548|false|false|false|||MRI
Finding|Gene or Genome|Past Medical History|2545,2548|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|Past Medical History|2545,2548|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|Past Medical History|2545,2548|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Event|Event|Past Medical History|2556,2563|false|false|false|||History
Finding|Conceptual Entity|Past Medical History|2556,2563|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|Past Medical History|2556,2563|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|Past Medical History|2556,2563|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|Past Medical History|2556,2566|false|false|false|C0262926|Medical History|History of
Disorder|Congenital Abnormality|Past Medical History|2567,2576|false|false|false|C0334044|Dysplasia|dysplasia
Event|Event|Past Medical History|2567,2576|false|false|false|||dysplasia
Disorder|Neoplastic Process|Past Medical History|2567,2584|false|false|false|C0347129|Dysplasia of anus|dysplasia of anus
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2580,2584|false|false|false|C0003461|Anus|anus
Disorder|Disease or Syndrome|Past Medical History|2580,2584|false|false|false|C0003462|Anus Diseases|anus
Event|Event|Past Medical History|2580,2584|false|false|false|||anus
Procedure|Health Care Activity|Past Medical History|2580,2584|false|false|false|C0870072|Procedure on anus|anus
Disorder|Mental or Behavioral Dysfunction|Past Medical History|2599,2625|false|false|false|C0005586;C1839839;C1852197;C1970943;C1970945;C2700438;C2700439;C2700440|Bipolar Disorder;MAJOR AFFECTIVE DISORDER 1;MAJOR AFFECTIVE DISORDER 2;MAJOR AFFECTIVE DISORDER 4;MAJOR AFFECTIVE DISORDER 6;MAJOR AFFECTIVE DISORDER 7;MAJOR AFFECTIVE DISORDER 8;MAJOR AFFECTIVE DISORDER 9|Bipolar affective disorder
Disorder|Mental or Behavioral Dysfunction|Past Medical History|2599,2648|false|false|false|C0338875|Bipolar affective disorder, currently manic, mild|Bipolar affective disorder, currently manic, mild
Disorder|Mental or Behavioral Dysfunction|Past Medical History|2607,2625|false|false|false|C0525045|Mood Disorders|affective disorder
Disorder|Disease or Syndrome|Past Medical History|2617,2625|false|false|false|C0012634|Disease|disorder
Event|Event|Past Medical History|2617,2625|false|false|false|||disorder
Disorder|Mental or Behavioral Dysfunction|Past Medical History|2637,2642|false|false|false|C0338831|Manic|manic
Event|Event|Past Medical History|2637,2642|false|false|false|||manic
Finding|Finding|Past Medical History|2637,2642|false|false|false|C0564408|Manic mood|manic
Event|Event|Past Medical History|2644,2648|false|false|false|||mild
Finding|Intellectual Product|Past Medical History|2644,2648|false|false|false|C1547225|Mild Severity of Illness Code|mild
Disorder|Disease or Syndrome|Past Medical History|2654,2658|false|false|false|C0038436;C0878676|6-pyruvoyl-tetrahydropterin synthase deficiency;Post-Traumatic Stress Disorder|PTSD
Disorder|Mental or Behavioral Dysfunction|Past Medical History|2654,2658|false|false|false|C0038436;C0878676|6-pyruvoyl-tetrahydropterin synthase deficiency;Post-Traumatic Stress Disorder|PTSD
Event|Event|Past Medical History|2654,2658|false|false|false|||PTSD
Event|Event|Past Medical History|2667,2674|false|false|false|||History
Finding|Conceptual Entity|Past Medical History|2667,2674|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|Past Medical History|2667,2674|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|Past Medical History|2667,2674|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|Past Medical History|2667,2677|false|false|false|C0262926|Medical History|History of
Disorder|Injury or Poisoning|Past Medical History|2678,2685|true|false|false|C0274659|Poisoning by cocaine|cocaine
Drug|Biomedical or Dental Material|Past Medical History|2678,2685|true|false|false|C0009170|cocaine|cocaine
Drug|Hazardous or Poisonous Substance|Past Medical History|2678,2685|true|false|false|C0009170|cocaine|cocaine
Drug|Organic Chemical|Past Medical History|2678,2685|true|false|false|C0009170|cocaine|cocaine
Drug|Pharmacologic Substance|Past Medical History|2678,2685|true|false|false|C0009170|cocaine|cocaine
Event|Event|Past Medical History|2678,2685|false|false|false|||cocaine
Procedure|Laboratory Procedure|Past Medical History|2678,2685|true|false|false|C0202362|Cocaine measurement|cocaine
Disorder|Injury or Poisoning|Past Medical History|2690,2696|true|false|false|C0161541|Poisoning by heroin|heroin
Drug|Hazardous or Poisonous Substance|Past Medical History|2690,2696|true|false|false|C0011892|heroin|heroin
Drug|Organic Chemical|Past Medical History|2690,2696|true|false|false|C0011892|heroin|heroin
Drug|Pharmacologic Substance|Past Medical History|2690,2696|true|false|false|C0011892|heroin|heroin
Event|Event|Past Medical History|2690,2696|false|false|false|||heroin
Event|Event|Past Medical History|2697,2700|false|false|false|||use
Finding|Functional Concept|Past Medical History|2697,2700|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|Past Medical History|2697,2700|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Event|Event|Family Medical History|2789,2796|true|false|false|||talking
Finding|Conceptual Entity|Family Medical History|2832,2839|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|brother
Finding|Idea or Concept|Family Medical History|2832,2839|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|brother
Event|Event|Family Medical History|2856,2861|false|false|false|||touch
Finding|Mental Process|Family Medical History|2856,2861|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Finding|Organ or Tissue Function|Family Medical History|2856,2861|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2856,2861|false|false|false|C0152054|Therapeutic Touch|touch
Event|Event|Family Medical History|2872,2877|false|false|false|||lives
Event|Event|Family Medical History|2897,2902|true|false|false|||aware
Finding|Mental Process|Family Medical History|2897,2902|true|false|false|C0004448|Awareness|aware
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2922,2927|true|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Family Medical History|2922,2927|true|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Family Medical History|2922,2927|true|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Family Medical History|2922,2927|true|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Family Medical History|2922,2927|true|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Family Medical History|2922,2927|true|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|Family Medical History|2922,2927|true|false|false|||liver
Finding|Finding|Family Medical History|2922,2927|true|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Family Medical History|2922,2927|true|false|false|C0872387|Procedures on liver|liver
Disorder|Disease or Syndrome|Family Medical History|2929,2936|true|false|false|C0012634|Disease|disease
Event|Event|Family Medical History|2929,2936|true|false|false|||disease
Drug|Amino Acid, Peptide, or Protein|Family Medical History|2940,2950|false|false|false|C3812393|ErbB Receptors|her family
Drug|Enzyme|Family Medical History|2940,2950|false|false|false|C3812393|ErbB Receptors|her family
Finding|Receptor|Family Medical History|2940,2950|false|false|false|C3812393|ErbB Receptors|her family
Finding|Classification|Family Medical History|2944,2950|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Family Medical History|2944,2950|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Family Medical History|2944,2950|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Family Medical History|2944,2950|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Procedure|Health Care Activity|General Exam|2971,2980|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|General Exam|2981,2989|false|false|false|||PHYSICAL
Finding|Finding|General Exam|2981,2989|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|General Exam|2981,2989|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|General Exam|2981,2989|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|General Exam|2981,2994|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|General Exam|2981,2994|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Event|Event|General Exam|2990,2994|false|false|false|||EXAM
Finding|Functional Concept|General Exam|2990,2994|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|2990,2994|false|false|false|C0582103|Medical Examination|EXAM
Event|Event|General Exam|3035,3042|false|false|false|||GENERAL
Finding|Classification|General Exam|3035,3042|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|General Exam|3035,3042|false|false|false|C3812897|General medical service|GENERAL
Disorder|Disease or Syndrome|General Exam|3049,3064|true|false|false|C0008715|Chronically Ill|chronically ill
Finding|Finding|General Exam|3049,3064|true|false|false|C2051413|Patient appears chronically ill|chronically ill
Finding|Sign or Symptom|General Exam|3061,3064|true|false|false|C0231218|Malaise|ill
Finding|Intellectual Product|General Exam|3087,3092|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|General Exam|3094,3102|true|false|false|||distress
Finding|Finding|General Exam|3094,3102|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|General Exam|3094,3102|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|General Exam|3105,3110|true|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|General Exam|3112,3118|true|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|General Exam|3112,3118|true|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|General Exam|3112,3118|true|false|false|||Sclera
Procedure|Health Care Activity|General Exam|3112,3118|true|false|false|C2228481|examination of sclera|Sclera
Event|Event|General Exam|3119,3128|true|false|false|||anicteric
Finding|Finding|General Exam|3119,3128|true|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|General Exam|3130,3133|true|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|General Exam|3130,3133|true|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Space or Junction|General Exam|3138,3142|true|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|General Exam|3138,3142|true|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|General Exam|3138,3142|true|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|General Exam|3138,3142|true|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|General Exam|3143,3150|true|false|false|||lesions
Finding|Finding|General Exam|3143,3150|true|false|false|C0221198|Lesion|lesions
Anatomy|Body Part, Organ, or Organ Component|General Exam|3153,3158|true|false|false|C0018787;C4037974|Chest>Heart;Heart|HEART
Disorder|Neoplastic Process|General Exam|3153,3158|true|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|HEART
Event|Event|General Exam|3153,3158|true|false|false|||HEART
Finding|Sign or Symptom|General Exam|3153,3158|true|false|false|C0795691|HEART PROBLEM|HEART
Event|Event|General Exam|3160,3163|true|false|false|||RRR
Event|Event|General Exam|3182,3189|true|false|false|||murmurs
Finding|Finding|General Exam|3182,3189|true|false|false|C0018808|Heart murmur|murmurs
Anatomy|Body Part, Organ, or Organ Component|General Exam|3192,3197|true|false|false|C0024109|Lung|LUNGS
Event|Event|General Exam|3199,3204|true|false|false|||Clear
Finding|Idea or Concept|General Exam|3199,3204|true|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|General Exam|3209,3216|true|false|false|||wheezes
Finding|Sign or Symptom|General Exam|3209,3216|true|false|false|C0043144|Wheezing|wheezes
Event|Event|General Exam|3218,3223|true|false|false|||rales
Finding|Finding|General Exam|3218,3223|true|false|false|C0034642;C0240859|Basilar Rales;Rales|rales
Event|Event|General Exam|3228,3235|true|false|false|||rhonchi
Finding|Finding|General Exam|3228,3235|true|false|false|C0035508|Rhonchi|rhonchi
Anatomy|Body Location or Region|General Exam|3238,3241|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|ABD
Disorder|Cell or Molecular Dysfunction|General Exam|3238,3241|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|ABD
Event|Event|General Exam|3238,3241|false|false|false|||ABD
Finding|Idea or Concept|General Exam|3243,3254|false|false|false|C0750502|Significant|Significant
Event|Event|General Exam|3255,3265|false|false|false|||distention
Finding|Finding|General Exam|3255,3265|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Finding|Pathologic Function|General Exam|3255,3265|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Anatomy|Body Part, Organ, or Organ Component|General Exam|3279,3284|false|false|false|C0042449|Veins|veins
Procedure|Therapeutic or Preventive Procedure|General Exam|3279,3284|false|false|false|C0398102|Procedure on vein|veins
Anatomy|Body Location or Region|General Exam|3294,3300|false|false|false|C0230171|Flank (surface region)|flanks
Event|Event|General Exam|3303,3312|false|false|false|||nontender
Event|Event|General Exam|3316,3325|false|false|false|||palpation
Procedure|Diagnostic Procedure|General Exam|3316,3325|false|false|false|C0030247|Palpation|palpation
Event|Event|General Exam|3327,3337|false|false|false|||tympanitic
Event|Event|General Exam|3341,3351|false|false|false|||percussion
Procedure|Diagnostic Procedure|General Exam|3341,3351|false|false|false|C0030987;C1880282|Dental Percussion;Percussion|percussion
Anatomy|Body Part, Organ, or Organ Component|General Exam|3360,3365|false|false|false|C0021853|Intestines|bowel
Phenomenon|Natural Phenomenon or Process|General Exam|3367,3373|false|false|false|C0037709||sounds
Disorder|Congenital Abnormality|General Exam|3376,3379|false|false|false|C0015306|Hereditary Multiple Exostoses|EXT
Event|Event|General Exam|3376,3379|false|false|false|||EXT
Finding|Gene or Genome|General Exam|3376,3379|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|EXT
Attribute|Clinical Attribute|General Exam|3388,3393|true|false|false|C1717255||edema
Event|Event|General Exam|3388,3393|true|false|false|||edema
Finding|Pathologic Function|General Exam|3388,3393|true|false|false|C0013604|Edema|edema
Drug|Food|General Exam|3409,3415|false|false|false|C5890763||pulses
Event|Event|General Exam|3409,3415|false|false|false|||pulses
Finding|Physiologic Function|General Exam|3409,3415|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|3409,3415|false|false|false|C0034107|Pulse taking|pulses
Attribute|Clinical Attribute|General Exam|3425,3430|true|false|false|C5890168||alert
Drug|Organic Chemical|General Exam|3425,3430|true|false|false|C0718338|Alert brand of caffeine|alert
Drug|Pharmacologic Substance|General Exam|3425,3430|true|false|false|C0718338|Alert brand of caffeine|alert
Event|Event|General Exam|3425,3430|true|false|false|||alert
Finding|Finding|General Exam|3425,3430|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Functional Concept|General Exam|3425,3430|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Intellectual Product|General Exam|3425,3430|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Event|Event|General Exam|3435,3443|true|false|false|||oriented
Finding|Finding|General Exam|3435,3443|true|false|false|C1961028|Oriented to place|oriented
Disorder|Mental or Behavioral Dysfunction|General Exam|3449,3457|true|false|false|C0009676|Confusion|confused
Event|Event|General Exam|3449,3457|true|false|false|||confused
Finding|Finding|General Exam|3449,3457|true|false|false|C0683369;C1547301|Clouded consciousness;Precaution Code - Confused|confused
Finding|Intellectual Product|General Exam|3449,3457|true|false|false|C0683369;C1547301|Clouded consciousness;Precaution Code - Confused|confused
Event|Event|General Exam|3462,3471|true|false|false|||asterixis
Finding|Sign or Symptom|General Exam|3462,3471|true|false|false|C0232766|Asterixis|asterixis
Finding|Body Substance|General Exam|3473,3482|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|3473,3482|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|3473,3482|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|3473,3482|true|false|false|C0030685|Patient Discharge|DISCHARGE
Attribute|Clinical Attribute|General Exam|3508,3511|false|false|false|C0871470|Systolic Pressure|SBP
Drug|Amino Acid, Peptide, or Protein|General Exam|3508,3511|false|false|false|C0085805|Androgen Binding Protein|SBP
Drug|Biologically Active Substance|General Exam|3508,3511|false|false|false|C0085805|Androgen Binding Protein|SBP
Event|Event|General Exam|3508,3511|false|false|false|||SBP
Finding|Gene or Genome|General Exam|3508,3511|false|false|false|C1705296;C3274833|CCHCR1 wt Allele;SHBG wt Allele|SBP
Procedure|Diagnostic Procedure|General Exam|3508,3511|false|false|false|C1306620|Systolic blood pressure measurement|SBP
Event|Event|General Exam|3539,3540|false|false|false|||/
Event|Event|General Exam|3560,3567|false|false|false|||GENERAL
Finding|Classification|General Exam|3560,3567|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|General Exam|3560,3567|false|false|false|C3812897|General medical service|GENERAL
Disorder|Disease or Syndrome|General Exam|3574,3589|true|false|false|C0008715|Chronically Ill|chronically ill
Finding|Finding|General Exam|3574,3589|true|false|false|C2051413|Patient appears chronically ill|chronically ill
Finding|Sign or Symptom|General Exam|3586,3589|true|false|false|C0231218|Malaise|ill
Finding|Intellectual Product|General Exam|3612,3617|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|General Exam|3619,3627|true|false|false|||distress
Finding|Finding|General Exam|3619,3627|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|General Exam|3619,3627|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|General Exam|3630,3635|true|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|General Exam|3637,3643|true|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|General Exam|3637,3643|true|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|General Exam|3637,3643|true|false|false|||Sclera
Procedure|Health Care Activity|General Exam|3637,3643|true|false|false|C2228481|examination of sclera|Sclera
Event|Event|General Exam|3644,3653|true|false|false|||anicteric
Finding|Finding|General Exam|3644,3653|true|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|General Exam|3655,3658|true|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|General Exam|3655,3658|true|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Space or Junction|General Exam|3663,3667|true|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|General Exam|3663,3667|true|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|General Exam|3663,3667|true|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|General Exam|3663,3667|true|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|General Exam|3668,3675|true|false|false|||lesions
Finding|Finding|General Exam|3668,3675|true|false|false|C0221198|Lesion|lesions
Anatomy|Body Part, Organ, or Organ Component|General Exam|3678,3683|true|false|false|C0018787;C4037974|Chest>Heart;Heart|HEART
Disorder|Neoplastic Process|General Exam|3678,3683|true|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|HEART
Event|Event|General Exam|3678,3683|true|false|false|||HEART
Finding|Sign or Symptom|General Exam|3678,3683|true|false|false|C0795691|HEART PROBLEM|HEART
Event|Event|General Exam|3685,3688|true|false|false|||RRR
Event|Event|General Exam|3707,3714|true|false|false|||murmurs
Finding|Finding|General Exam|3707,3714|true|false|false|C0018808|Heart murmur|murmurs
Anatomy|Body Part, Organ, or Organ Component|General Exam|3717,3722|true|false|false|C0024109|Lung|LUNGS
Event|Event|General Exam|3724,3729|true|false|false|||Clear
Finding|Idea or Concept|General Exam|3724,3729|true|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|General Exam|3734,3741|true|false|false|||wheezes
Finding|Sign or Symptom|General Exam|3734,3741|true|false|false|C0043144|Wheezing|wheezes
Event|Event|General Exam|3743,3748|true|false|false|||rales
Finding|Finding|General Exam|3743,3748|true|false|false|C0034642;C0240859|Basilar Rales;Rales|rales
Event|Event|General Exam|3753,3760|true|false|false|||rhonchi
Finding|Finding|General Exam|3753,3760|true|false|false|C0035508|Rhonchi|rhonchi
Anatomy|Body Location or Region|General Exam|3763,3766|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|ABD
Disorder|Cell or Molecular Dysfunction|General Exam|3763,3766|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|ABD
Event|Event|General Exam|3763,3766|false|false|false|||ABD
Finding|Idea or Concept|General Exam|3768,3779|false|false|false|C0750502|Significant|Significant
Event|Event|General Exam|3780,3790|false|false|false|||distention
Finding|Finding|General Exam|3780,3790|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Finding|Pathologic Function|General Exam|3780,3790|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Anatomy|Body Part, Organ, or Organ Component|General Exam|3804,3809|false|false|false|C0042449|Veins|veins
Procedure|Therapeutic or Preventive Procedure|General Exam|3804,3809|false|false|false|C0398102|Procedure on vein|veins
Anatomy|Body Location or Region|General Exam|3819,3825|false|false|false|C0230171|Flank (surface region)|flanks
Event|Event|General Exam|3828,3837|false|false|false|||nontender
Event|Event|General Exam|3841,3850|false|false|false|||palpation
Procedure|Diagnostic Procedure|General Exam|3841,3850|false|false|false|C0030247|Palpation|palpation
Event|Event|General Exam|3852,3862|false|false|false|||tympanitic
Event|Event|General Exam|3866,3876|false|false|false|||percussion
Procedure|Diagnostic Procedure|General Exam|3866,3876|false|false|false|C0030987;C1880282|Dental Percussion;Percussion|percussion
Anatomy|Body Part, Organ, or Organ Component|General Exam|3885,3890|false|false|false|C0021853|Intestines|bowel
Phenomenon|Natural Phenomenon or Process|General Exam|3892,3898|false|false|false|C0037709||sounds
Disorder|Congenital Abnormality|General Exam|3901,3904|false|false|false|C0015306|Hereditary Multiple Exostoses|EXT
Event|Event|General Exam|3901,3904|false|false|false|||EXT
Finding|Gene or Genome|General Exam|3901,3904|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|EXT
Attribute|Clinical Attribute|General Exam|3913,3918|true|false|false|C1717255||edema
Event|Event|General Exam|3913,3918|true|false|false|||edema
Finding|Pathologic Function|General Exam|3913,3918|true|false|false|C0013604|Edema|edema
Drug|Food|General Exam|3934,3940|false|false|false|C5890763||pulses
Event|Event|General Exam|3934,3940|false|false|false|||pulses
Finding|Physiologic Function|General Exam|3934,3940|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|3934,3940|false|false|false|C0034107|Pulse taking|pulses
Attribute|Clinical Attribute|General Exam|3950,3955|true|false|false|C5890168||alert
Drug|Organic Chemical|General Exam|3950,3955|true|false|false|C0718338|Alert brand of caffeine|alert
Drug|Pharmacologic Substance|General Exam|3950,3955|true|false|false|C0718338|Alert brand of caffeine|alert
Event|Event|General Exam|3950,3955|true|false|false|||alert
Finding|Finding|General Exam|3950,3955|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Functional Concept|General Exam|3950,3955|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Intellectual Product|General Exam|3950,3955|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Event|Event|General Exam|3960,3968|true|false|false|||oriented
Finding|Finding|General Exam|3960,3968|true|false|false|C1961028|Oriented to place|oriented
Disorder|Mental or Behavioral Dysfunction|General Exam|3974,3982|true|false|false|C0009676|Confusion|confused
Event|Event|General Exam|3974,3982|true|false|false|||confused
Finding|Finding|General Exam|3974,3982|true|false|false|C0683369;C1547301|Clouded consciousness;Precaution Code - Confused|confused
Finding|Intellectual Product|General Exam|3974,3982|true|false|false|C0683369;C1547301|Clouded consciousness;Precaution Code - Confused|confused
Event|Event|General Exam|3987,3996|true|false|false|||asterixis
Finding|Sign or Symptom|General Exam|3987,3996|true|false|false|C0232766|Asterixis|asterixis
Event|Event|General Exam|4018,4022|false|false|false|||LABS
Lab|Laboratory or Test Result|General Exam|4018,4022|false|false|false|C0587081|Laboratory test finding|LABS
Procedure|Health Care Activity|General Exam|4026,4035|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Disorder|Disease or Syndrome|General Exam|4049,4054|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4049,4054|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4049,4054|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|4064,4067|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|4084,4089|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4084,4089|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4084,4089|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|General Exam|4111,4116|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4111,4116|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4111,4116|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|General Exam|4138,4143|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4138,4143|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4138,4143|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|General Exam|4165,4170|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4165,4170|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4165,4170|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|General Exam|4187,4192|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4187,4192|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4187,4192|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Event|General Exam|4198,4202|false|false|false|||LABS
Lab|Laboratory or Test Result|General Exam|4198,4202|false|false|false|C0587081|Laboratory test finding|LABS
Finding|Body Substance|General Exam|4206,4215|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|4206,4215|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|4206,4215|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|4206,4215|false|false|false|C0030685|Patient Discharge|DISCHARGE
Disorder|Disease or Syndrome|General Exam|4229,4234|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4229,4234|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4229,4234|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|4244,4247|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|4264,4269|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4264,4269|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4264,4269|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|General Exam|4290,4295|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4290,4295|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4290,4295|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|General Exam|4317,4322|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4317,4322|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4317,4322|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|General Exam|4344,4349|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4344,4349|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4344,4349|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Event|General Exam|4355,4360|false|false|false|||MICRO
Finding|Conceptual Entity|General Exam|4355,4360|false|false|false|C3811161;C4049106|Micro (prefix);Microbiology - Laboratory Class|MICRO
Finding|Intellectual Product|General Exam|4355,4360|false|false|false|C3811161;C4049106|Micro (prefix);Microbiology - Laboratory Class|MICRO
Procedure|Laboratory Procedure|General Exam|4355,4360|false|false|false|C0085672|Microbiology procedure|MICRO
Finding|Body Substance|General Exam|4375,4380|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|4375,4380|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|4375,4380|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Event|Event|General Exam|4386,4392|false|false|false|||Source
Finding|Finding|General Exam|4386,4392|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|Source
Finding|Functional Concept|General Exam|4386,4392|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|Source
Finding|Intellectual Product|General Exam|4386,4392|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|Source
Finding|Idea or Concept|General Exam|4431,4436|false|false|false|C1546485|Diagnosis Type - Final|FINAL
Finding|Intellectual Product|General Exam|4431,4443|false|false|false|C0460114|Final report|FINAL REPORT
Attribute|Clinical Attribute|General Exam|4437,4443|false|false|false|C4255046||REPORT
Event|Event|General Exam|4437,4443|false|false|false|||REPORT
Finding|Intellectual Product|General Exam|4437,4443|false|false|false|C0684224|Report (document)|REPORT
Procedure|Health Care Activity|General Exam|4437,4443|false|false|false|C0700287|Reporting|REPORT
Finding|Body Substance|General Exam|4452,4457|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|4452,4457|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|4452,4457|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Procedure|Laboratory Procedure|General Exam|4452,4465|false|false|false|C0430404|Urine culture|URINE CULTURE
Drug|Biomedical or Dental Material|General Exam|4458,4465|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|General Exam|4458,4465|false|false|false|||CULTURE
Finding|Functional Concept|General Exam|4458,4465|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|General Exam|4458,4465|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|General Exam|4458,4465|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|General Exam|4467,4472|false|false|false|||Final
Finding|Idea or Concept|General Exam|4467,4472|false|false|false|C1546485|Diagnosis Type - Final|Final
Event|Event|General Exam|4485,4490|false|false|false|||MIXED
Anatomy|Cell|General Exam|4514,4520|false|false|false|C1947989|Colony (cells or organisms)|COLONY
Event|Event|General Exam|4529,4539|false|false|false|||CONSISTENT
Finding|Idea or Concept|General Exam|4529,4539|false|false|false|C0332290|Consistent with|CONSISTENT
Anatomy|Body System|General Exam|4546,4550|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|General Exam|4546,4550|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|General Exam|4546,4550|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|General Exam|4546,4550|false|false|false|||SKIN
Finding|Body Substance|General Exam|4546,4550|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|General Exam|4546,4550|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Event|Event|General Exam|4560,4561|false|false|false|||/
Anatomy|Body Part, Organ, or Organ Component|General Exam|4564,4571|false|false|false|C0017420;C0559522|Genital system;Genitalia|GENITAL
Anatomy|Body System|General Exam|4564,4571|false|false|false|C0017420;C0559522|Genital system;Genitalia|GENITAL
Finding|Body Substance|General Exam|4564,4571|false|false|false|C1546649;C1550642|Specimen Type - Genital|GENITAL
Finding|Intellectual Product|General Exam|4564,4571|false|false|false|C1546649;C1550642|Specimen Type - Genital|GENITAL
Event|Event|General Exam|4572,4585|false|false|false|||CONTAMINATION
Finding|Idea or Concept|General Exam|4572,4585|false|false|false|C2349974|Contamination|CONTAMINATION
Phenomenon|Human-caused Phenomenon or Process|General Exam|4572,4585|false|false|false|C0259846|adulteration|CONTAMINATION
Anatomy|Body Location or Region|General Exam|4601,4611|false|false|false|C0031153;C0442034|Peritoneum;peritoneal|PERITONEAL
Anatomy|Tissue|General Exam|4601,4611|false|false|false|C0031153;C0442034|Peritoneum;peritoneal|PERITONEAL
Finding|Body Substance|General Exam|4601,4617|false|false|false|C0003964|Peritoneal fluid (substance)|PERITONEAL FLUID
Procedure|Laboratory Procedure|General Exam|4601,4617|false|false|false|C2053903|Peritoneal fluid analysis|PERITONEAL FLUID
Drug|Substance|General Exam|4612,4617|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|FLUID
Event|Event|General Exam|4612,4617|false|false|false|||FLUID
Finding|Intellectual Product|General Exam|4612,4617|false|false|false|C1546638|Fluid Specimen Code|FLUID
Finding|Body Substance|General Exam|4612,4633|false|false|false|C0003964|Peritoneal fluid (substance)|FLUID      PERITONEAL
Anatomy|Body Location or Region|General Exam|4623,4633|false|false|false|C0031153;C0442034|Peritoneum;peritoneal|PERITONEAL
Anatomy|Tissue|General Exam|4623,4633|false|false|false|C0031153;C0442034|Peritoneum;peritoneal|PERITONEAL
Finding|Body Substance|General Exam|4623,4639|false|false|false|C0003964|Peritoneal fluid (substance)|PERITONEAL FLUID
Procedure|Laboratory Procedure|General Exam|4623,4639|false|false|false|C2053903|Peritoneal fluid analysis|PERITONEAL FLUID
Drug|Substance|General Exam|4634,4639|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|FLUID
Event|Event|General Exam|4634,4639|false|false|false|||FLUID
Finding|Intellectual Product|General Exam|4634,4639|false|false|false|C1546638|Fluid Specimen Code|FLUID
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|4646,4656|false|false|false|C0061856|Gram's stain|GRAM STAIN
Drug|Organic Chemical|General Exam|4646,4656|false|false|false|C0061856|Gram's stain|GRAM STAIN
Procedure|Laboratory Procedure|General Exam|4646,4656|false|false|false|C0200966|Bacterial stain, routine|GRAM STAIN
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|4651,4656|false|false|false|C0038128|Stains|STAIN
Event|Event|General Exam|4651,4656|false|false|false|||STAIN
Procedure|Laboratory Procedure|General Exam|4651,4656|false|false|false|C0487602|Staining method|STAIN
Finding|Idea or Concept|General Exam|4658,4663|false|false|false|C1546485|Diagnosis Type - Final|Final
Event|Event|General Exam|4696,4701|false|false|false|||FIELD
Finding|Conceptual Entity|General Exam|4696,4701|false|false|false|C1521738;C2346620;C2349184|Field;Force Field;Knowledge Field|FIELD
Procedure|Health Care Activity|General Exam|4696,4701|false|false|false|C1553496|field - patient encounter|FIELD
Event|Event|General Exam|4706,4723|false|false|false|||POLYMORPHONUCLEAR
Anatomy|Cell|General Exam|4725,4735|false|false|false|C0023516|Leukocytes|LEUKOCYTES
Event|Event|General Exam|4725,4735|false|false|false|||LEUKOCYTES
Finding|Body Substance|General Exam|4725,4735|false|false|false|C1547962;C1550647|Specimen Type - Leukocytes|LEUKOCYTES
Finding|Intellectual Product|General Exam|4725,4735|false|false|false|C1547962;C1550647|Specimen Type - Leukocytes|LEUKOCYTES
Finding|Finding|General Exam|4747,4766|true|false|false|C2924473|Microorganisms seen|MICROORGANISMS SEEN
Event|Event|General Exam|4762,4766|true|false|false|||SEEN
Event|Activity|General Exam|4798,4803|false|false|false|C1947932|Smear - instruction imperative|smear
Event|Event|General Exam|4798,4803|false|false|false|||smear
Finding|Functional Concept|General Exam|4798,4803|false|false|false|C3872789|Smearing technique|smear
Procedure|Diagnostic Procedure|General Exam|4798,4803|false|false|false|C0444186|Smear test|smear
Event|Event|General Exam|4821,4827|false|false|false|||method
Finding|Functional Concept|General Exam|4821,4827|false|false|false|C0025663;C0449851;C2828387|Method, LOINC Axis 6;Methods;Techniques|method
Finding|Intellectual Product|General Exam|4821,4827|false|false|false|C0025663;C0449851;C2828387|Method, LOINC Axis 6;Methods;Techniques|method
Event|Event|General Exam|4852,4862|false|false|false|||hematology
Finding|Intellectual Product|General Exam|4852,4862|false|false|false|C1547985|Diagnostic Service Section ID - Hematology|hematology
Procedure|Laboratory Procedure|General Exam|4852,4862|false|false|false|C0018941;C0200627;C2183233|Hematologic Tests;Hematology procedure;diagnostic service sources hematology (procedure)|hematology
Anatomy|Cell|General Exam|4882,4898|false|false|false|C0023516|Leukocytes|white blood cell
Lab|Laboratory or Test Result|General Exam|4882,4904|false|false|false|C0427512||white blood cell count
Procedure|Laboratory Procedure|General Exam|4882,4904|false|false|false|C0023508|White Blood Cell Count procedure|white blood cell count
Disorder|Disease or Syndrome|General Exam|4888,4893|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|General Exam|4888,4893|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Anatomy|Cell|General Exam|4888,4898|false|false|false|C0005773|Blood Cells|blood cell
Procedure|Laboratory Procedure|General Exam|4888,4904|false|false|false|C0005771;C0009555|Blood Cell Count;Complete Blood Count|blood cell count
Anatomy|Cell|General Exam|4894,4898|false|false|false|C0007634|Cells|cell
Finding|Gene or Genome|General Exam|4894,4898|false|false|false|C1413336;C1413337|CEL gene;CELP gene|cell
Procedure|Laboratory Procedure|General Exam|4894,4904|false|false|false|C0007584|Cell Count|cell count
Event|Event|General Exam|4899,4904|false|false|false|||count
Drug|Substance|General Exam|4912,4917|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|FLUID
Event|Event|General Exam|4912,4917|false|false|false|||FLUID
Finding|Intellectual Product|General Exam|4912,4917|false|false|false|C1546638|Fluid Specimen Code|FLUID
Drug|Biomedical or Dental Material|General Exam|4918,4925|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|General Exam|4918,4925|false|false|false|||CULTURE
Finding|Functional Concept|General Exam|4918,4925|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|General Exam|4918,4925|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|General Exam|4918,4925|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|General Exam|4927,4932|false|false|false|||Final
Finding|Idea or Concept|General Exam|4927,4932|false|false|false|C1546485|Diagnosis Type - Final|Final
Event|Event|General Exam|4944,4950|true|false|false|||GROWTH
Finding|Finding|General Exam|4944,4950|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organ or Tissue Function|General Exam|4944,4950|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organism Function|General Exam|4944,4950|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Physiologic Function|General Exam|4944,4950|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Phenomenon|Phenomenon or Process|General Exam|4944,4950|true|false|false|C2911660|Growth action|GROWTH
Procedure|Laboratory Procedure|General Exam|4957,4974|false|false|false|C1273935|Anaerobic microbial culture|ANAEROBIC CULTURE
Drug|Biomedical or Dental Material|General Exam|4967,4974|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|General Exam|4967,4974|false|false|false|||CULTURE
Finding|Functional Concept|General Exam|4967,4974|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|General Exam|4967,4974|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|General Exam|4967,4974|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|General Exam|4996,5002|true|false|false|||GROWTH
Finding|Finding|General Exam|4996,5002|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organ or Tissue Function|General Exam|4996,5002|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organism Function|General Exam|4996,5002|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Physiologic Function|General Exam|4996,5002|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Phenomenon|Phenomenon or Process|General Exam|4996,5002|true|false|false|C2911660|Growth action|GROWTH
Anatomy|Body Location or Region|General Exam|5017,5027|false|false|false|C0031153;C0442034|Peritoneum;peritoneal|PERITONEAL
Anatomy|Tissue|General Exam|5017,5027|false|false|false|C0031153;C0442034|Peritoneum;peritoneal|PERITONEAL
Finding|Body Substance|General Exam|5017,5033|false|false|false|C0003964|Peritoneal fluid (substance)|PERITONEAL FLUID
Procedure|Laboratory Procedure|General Exam|5017,5033|false|false|false|C2053903|Peritoneal fluid analysis|PERITONEAL FLUID
Drug|Substance|General Exam|5028,5033|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|FLUID
Event|Event|General Exam|5028,5033|false|false|false|||FLUID
Finding|Intellectual Product|General Exam|5028,5033|false|false|false|C1546638|Fluid Specimen Code|FLUID
Finding|Body Substance|General Exam|5028,5049|false|false|false|C0003964|Peritoneal fluid (substance)|FLUID      PERITONEAL
Anatomy|Body Location or Region|General Exam|5039,5049|false|false|false|C0031153;C0442034|Peritoneum;peritoneal|PERITONEAL
Anatomy|Tissue|General Exam|5039,5049|false|false|false|C0031153;C0442034|Peritoneum;peritoneal|PERITONEAL
Finding|Body Substance|General Exam|5039,5055|false|false|false|C0003964|Peritoneal fluid (substance)|PERITONEAL FLUID
Procedure|Laboratory Procedure|General Exam|5039,5055|false|false|false|C2053903|Peritoneal fluid analysis|PERITONEAL FLUID
Drug|Substance|General Exam|5050,5055|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|FLUID
Event|Event|General Exam|5050,5055|false|false|false|||FLUID
Finding|Intellectual Product|General Exam|5050,5055|false|false|false|C1546638|Fluid Specimen Code|FLUID
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|5062,5072|false|false|false|C0061856|Gram's stain|GRAM STAIN
Drug|Organic Chemical|General Exam|5062,5072|false|false|false|C0061856|Gram's stain|GRAM STAIN
Procedure|Laboratory Procedure|General Exam|5062,5072|false|false|false|C0200966|Bacterial stain, routine|GRAM STAIN
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|5067,5072|false|false|false|C0038128|Stains|STAIN
Event|Event|General Exam|5067,5072|false|false|false|||STAIN
Procedure|Laboratory Procedure|General Exam|5067,5072|false|false|false|C0487602|Staining method|STAIN
Finding|Idea or Concept|General Exam|5074,5079|false|false|false|C1546485|Diagnosis Type - Final|Final
Event|Event|General Exam|5112,5117|false|false|false|||FIELD
Finding|Conceptual Entity|General Exam|5112,5117|false|false|false|C1521738;C2346620;C2349184|Field;Force Field;Knowledge Field|FIELD
Procedure|Health Care Activity|General Exam|5112,5117|false|false|false|C1553496|field - patient encounter|FIELD
Event|Event|General Exam|5122,5139|false|false|false|||POLYMORPHONUCLEAR
Anatomy|Cell|General Exam|5141,5151|false|false|false|C0023516|Leukocytes|LEUKOCYTES
Event|Event|General Exam|5141,5151|false|false|false|||LEUKOCYTES
Finding|Body Substance|General Exam|5141,5151|false|false|false|C1547962;C1550647|Specimen Type - Leukocytes|LEUKOCYTES
Finding|Intellectual Product|General Exam|5141,5151|false|false|false|C1547962;C1550647|Specimen Type - Leukocytes|LEUKOCYTES
Finding|Finding|General Exam|5163,5182|true|false|false|C2924473|Microorganisms seen|MICROORGANISMS SEEN
Event|Event|General Exam|5178,5182|true|false|false|||SEEN
Event|Activity|General Exam|5214,5219|false|false|false|C1947932|Smear - instruction imperative|smear
Event|Event|General Exam|5214,5219|false|false|false|||smear
Finding|Functional Concept|General Exam|5214,5219|false|false|false|C3872789|Smearing technique|smear
Procedure|Diagnostic Procedure|General Exam|5214,5219|false|false|false|C0444186|Smear test|smear
Event|Event|General Exam|5237,5243|false|false|false|||method
Finding|Functional Concept|General Exam|5237,5243|false|false|false|C0025663;C0449851;C2828387|Method, LOINC Axis 6;Methods;Techniques|method
Finding|Intellectual Product|General Exam|5237,5243|false|false|false|C0025663;C0449851;C2828387|Method, LOINC Axis 6;Methods;Techniques|method
Event|Event|General Exam|5268,5278|false|false|false|||hematology
Finding|Intellectual Product|General Exam|5268,5278|false|false|false|C1547985|Diagnostic Service Section ID - Hematology|hematology
Procedure|Laboratory Procedure|General Exam|5268,5278|false|false|false|C0018941;C0200627;C2183233|Hematologic Tests;Hematology procedure;diagnostic service sources hematology (procedure)|hematology
Anatomy|Cell|General Exam|5298,5314|false|false|false|C0023516|Leukocytes|white blood cell
Lab|Laboratory or Test Result|General Exam|5298,5320|false|false|false|C0427512||white blood cell count
Procedure|Laboratory Procedure|General Exam|5298,5320|false|false|false|C0023508|White Blood Cell Count procedure|white blood cell count
Disorder|Disease or Syndrome|General Exam|5304,5309|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|General Exam|5304,5309|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Anatomy|Cell|General Exam|5304,5314|false|false|false|C0005773|Blood Cells|blood cell
Procedure|Laboratory Procedure|General Exam|5304,5320|false|false|false|C0005771;C0009555|Blood Cell Count;Complete Blood Count|blood cell count
Anatomy|Cell|General Exam|5310,5314|false|false|false|C0007634|Cells|cell
Finding|Gene or Genome|General Exam|5310,5314|false|false|false|C1413336;C1413337|CEL gene;CELP gene|cell
Procedure|Laboratory Procedure|General Exam|5310,5320|false|false|false|C0007584|Cell Count|cell count
Event|Event|General Exam|5315,5320|false|false|false|||count
Drug|Substance|General Exam|5328,5333|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|FLUID
Event|Event|General Exam|5328,5333|false|false|false|||FLUID
Finding|Intellectual Product|General Exam|5328,5333|false|false|false|C1546638|Fluid Specimen Code|FLUID
Drug|Biomedical or Dental Material|General Exam|5334,5341|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|General Exam|5334,5341|false|false|false|||CULTURE
Finding|Functional Concept|General Exam|5334,5341|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|General Exam|5334,5341|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|General Exam|5334,5341|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|General Exam|5343,5348|false|false|false|||Final
Finding|Idea or Concept|General Exam|5343,5348|false|false|false|C1546485|Diagnosis Type - Final|Final
Event|Event|General Exam|5360,5366|true|false|false|||GROWTH
Finding|Finding|General Exam|5360,5366|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organ or Tissue Function|General Exam|5360,5366|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organism Function|General Exam|5360,5366|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Physiologic Function|General Exam|5360,5366|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Phenomenon|Phenomenon or Process|General Exam|5360,5366|true|false|false|C2911660|Growth action|GROWTH
Procedure|Laboratory Procedure|General Exam|5373,5390|false|false|false|C1273935|Anaerobic microbial culture|ANAEROBIC CULTURE
Drug|Biomedical or Dental Material|General Exam|5383,5390|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|General Exam|5383,5390|false|false|false|||CULTURE
Finding|Functional Concept|General Exam|5383,5390|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|General Exam|5383,5390|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|General Exam|5383,5390|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|General Exam|5412,5418|true|false|false|||GROWTH
Finding|Finding|General Exam|5412,5418|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organ or Tissue Function|General Exam|5412,5418|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organism Function|General Exam|5412,5418|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Physiologic Function|General Exam|5412,5418|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Phenomenon|Phenomenon or Process|General Exam|5412,5418|true|false|false|C2911660|Growth action|GROWTH
Event|Event|General Exam|5433,5437|false|false|false|||Para
Finding|Finding|General Exam|5433,5437|false|false|false|C0030563|Parity|Para
Disorder|Disease or Syndrome|General Exam|5451,5458|false|false|false|C0003962|Ascites|ASCITES
Event|Event|General Exam|5451,5458|false|false|false|||ASCITES
Finding|Pathologic Function|General Exam|5451,5458|false|false|false|C5441966|Peritoneal Effusion|ASCITES
Disorder|Disease or Syndrome|General Exam|5480,5487|false|false|false|C0003962|Ascites|ASCITES
Event|Event|General Exam|5480,5487|false|false|false|||ASCITES
Finding|Pathologic Function|General Exam|5480,5487|false|false|false|C5441966|Peritoneal Effusion|ASCITES
Event|Event|General Exam|5493,5500|false|false|false|||IMAGING
Finding|Finding|General Exam|5493,5500|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|General Exam|5493,5500|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Event|Event|General Exam|5506,5509|true|false|false|||CXR
Procedure|Diagnostic Procedure|General Exam|5506,5509|true|false|false|C0039985|Plain chest X-ray|CXR
Finding|Intellectual Product|General Exam|5514,5519|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Location or Region|General Exam|5520,5535|true|false|false|C0553534|Cardiopulmonary|cardiopulmonary
Disorder|Disease or Syndrome|General Exam|5520,5535|true|false|false|C4072686|Cardiovascular disease+Pulmonary disease|cardiopulmonary
Disorder|Congenital Abnormality|General Exam|5536,5547|true|false|false|C0000768|Congenital Abnormality|abnormality
Event|Event|General Exam|5536,5547|true|false|false|||abnormality
Finding|Finding|General Exam|5536,5547|true|false|false|C1704258|Abnormality|abnormality
Anatomy|Body Location or Region|General Exam|5555,5558|false|false|false|C0230177|Structure of right upper quadrant of abdomen|RUQ
Event|Event|General Exam|5578,5584|false|false|false|||coarse
Anatomy|Body Part, Organ, or Organ Component|General Exam|5597,5602|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|General Exam|5597,5602|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|General Exam|5597,5602|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|General Exam|5597,5602|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|General Exam|5597,5602|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|General Exam|5597,5602|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Finding|Finding|General Exam|5597,5602|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|General Exam|5597,5602|false|false|false|C0872387|Procedures on liver|liver
Event|Event|General Exam|5615,5625|false|false|false|||consistent
Finding|Idea or Concept|General Exam|5615,5625|false|false|false|C0332290|Consistent with|consistent
Event|Event|General Exam|5634,5641|false|false|false|||history
Finding|Conceptual Entity|General Exam|5634,5641|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|General Exam|5634,5641|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|General Exam|5634,5641|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|General Exam|5634,5644|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|General Exam|5645,5654|false|false|false|C0023890;C1623038|Cirrhosis;Liver Cirrhosis|cirrhosis
Event|Event|General Exam|5645,5654|false|false|false|||cirrhosis
Finding|Finding|General Exam|5661,5669|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|General Exam|5661,5669|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Disorder|Disease or Syndrome|General Exam|5670,5677|false|false|false|C0003962|Ascites|ascites
Event|Event|General Exam|5670,5677|false|false|false|||ascites
Finding|Pathologic Function|General Exam|5670,5677|false|false|false|C5441966|Peritoneal Effusion|ascites
Finding|Intellectual Product|General Exam|5684,5690|false|false|false|C0030650|Legal patent|Patent
Anatomy|Body Location or Region|General Exam|5691,5697|false|false|false|C0205054|Hepatic|portal
Anatomy|Body Part, Organ, or Organ Component|General Exam|5691,5702|false|false|false|C0032718;C1305775;C4266644|Abdomen>Portal vein;Portal vein structure|portal vein
Anatomy|Body Part, Organ, or Organ Component|General Exam|5698,5702|false|false|false|C0042449|Veins|vein
Disorder|Disease or Syndrome|Hospital Course|5738,5741|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Disorder|Virus|Hospital Course|5738,5741|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Drug|Immunologic Factor|Hospital Course|5738,5741|false|false|false|C0086413|HIV Vaccine|HIV
Drug|Pharmacologic Substance|Hospital Course|5738,5741|false|false|false|C0086413|HIV Vaccine|HIV
Event|Event|Hospital Course|5738,5741|false|false|false|||HIV
Event|Event|Hospital Course|5745,5750|false|false|false|||HAART
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5745,5750|false|false|false|C0887947|Antiretroviral Therapy, Highly Active|HAART
Disorder|Disease or Syndrome|Hospital Course|5752,5755|false|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|HCV
Disorder|Virus|Hospital Course|5752,5755|false|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|HCV
Event|Event|Hospital Course|5752,5755|false|false|false|||HCV
Disorder|Disease or Syndrome|Hospital Course|5756,5765|false|false|false|C0023890;C1623038|Cirrhosis;Liver Cirrhosis|cirrhosis
Event|Event|Hospital Course|5756,5765|false|false|false|||cirrhosis
Disorder|Disease or Syndrome|Hospital Course|5771,5778|false|false|false|C0003962|Ascites|ascites
Event|Event|Hospital Course|5771,5778|false|false|false|||ascites
Finding|Pathologic Function|Hospital Course|5771,5778|false|false|false|C5441966|Peritoneal Effusion|ascites
Event|Event|Hospital Course|5783,5785|false|false|false|||HE
Event|Event|Hospital Course|5792,5796|false|false|false|||IVDU
Finding|Individual Behavior|Hospital Course|5792,5796|false|false|false|C0699778|intravenous drug use|IVDU
Disorder|Disease or Syndrome|Hospital Course|5798,5802|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|5798,5802|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|5798,5802|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|5798,5802|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Mental or Behavioral Dysfunction|Hospital Course|5804,5820|false|false|false|C0005586|Bipolar Disorder|bipolar disorder
Disorder|Disease or Syndrome|Hospital Course|5812,5820|false|false|false|C0012634|Disease|disorder
Event|Event|Hospital Course|5812,5820|false|false|false|||disorder
Event|Event|Hospital Course|5821,5829|false|false|false|||presents
Anatomy|Body Location or Region|Hospital Course|5835,5844|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|Hospital Course|5835,5855|false|false|false|C0232487|Abdominal discomfort|abdominal discomfort
Event|Event|Hospital Course|5845,5855|false|false|false|||discomfort
Finding|Sign or Symptom|Hospital Course|5845,5855|false|false|false|C2364135|Discomfort|discomfort
Disorder|Disease or Syndrome|Hospital Course|5868,5875|false|false|false|C0003962|Ascites|ascites
Event|Event|Hospital Course|5868,5875|false|false|false|||ascites
Finding|Pathologic Function|Hospital Course|5868,5875|false|false|false|C5441966|Peritoneal Effusion|ascites
Disorder|Disease or Syndrome|Hospital Course|5883,5890|false|false|false|C0003962|Ascites|ASCITES
Event|Event|Hospital Course|5883,5890|false|false|false|||ASCITES
Finding|Pathologic Function|Hospital Course|5883,5890|false|false|false|C5441966|Peritoneal Effusion|ASCITES
Drug|Pharmacologic Substance|Hospital Course|5896,5904|false|false|false|C0012798;C5399719|Diuretic [APC];Diuretics|diuretic
Event|Event|Hospital Course|5905,5915|false|false|false|||refractory
Finding|Functional Concept|Hospital Course|5905,5915|false|false|false|C0205269|Unresponsive to Treatment|refractory
Event|Event|Hospital Course|5927,5930|false|false|false|||tap
Finding|Gene or Genome|Hospital Course|5927,5930|false|false|false|C1414636;C1417898;C1419923;C1864009;C1865183|FLNB gene;NXF1 gene;SEC14L2 gene;TRACHEAL ANTIMICROBIAL PEPTIDE;USO1 gene|tap
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5927,5930|false|false|false|C0034115|Paracentesis|tap
Finding|Gene or Genome|Hospital Course|5947,5950|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|Hospital Course|5959,5966|false|false|false|||removed
Event|Event|Hospital Course|5987,5992|false|false|false|||built
Finding|Finding|Hospital Course|5996,6004|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|Hospital Course|5996,6004|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Disorder|Disease or Syndrome|Hospital Course|6006,6013|false|false|false|C0003962|Ascites|ascites
Event|Event|Hospital Course|6006,6013|false|false|false|||ascites
Finding|Pathologic Function|Hospital Course|6006,6013|false|false|false|C5441966|Peritoneal Effusion|ascites
Disorder|Disease or Syndrome|Hospital Course|6015,6025|false|false|false|C0009450|Communicable Diseases|Infectious
Event|Event|Hospital Course|6033,6041|false|false|false|||negative
Finding|Classification|Hospital Course|6033,6041|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|6033,6041|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|6033,6041|false|false|false|C5237010|Expression Negative|negative
Event|Event|Hospital Course|6048,6051|false|false|false|||CXR
Procedure|Diagnostic Procedure|Hospital Course|6048,6051|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|Hospital Course|6052,6057|false|false|false|||clear
Finding|Idea or Concept|Hospital Course|6052,6057|false|false|false|C1550016|Remote control command - Clear|clear
Event|Event|Hospital Course|6059,6061|false|false|false|||UA
Event|Event|Hospital Course|6063,6075|false|false|false|||contaminated
Finding|Finding|Hospital Course|6063,6075|false|false|false|C0205279;C1548222;C1548791;C2349974|Bed Status - Contaminated;Contaminated;Contamination;Specimen Condition - Contaminated|contaminated
Finding|Functional Concept|Hospital Course|6063,6075|false|false|false|C0205279;C1548222;C1548791;C2349974|Bed Status - Contaminated;Contaminated;Contamination;Specimen Condition - Contaminated|contaminated
Finding|Idea or Concept|Hospital Course|6063,6075|false|false|false|C0205279;C1548222;C1548791;C2349974|Bed Status - Contaminated;Contaminated;Contamination;Specimen Condition - Contaminated|contaminated
Disorder|Cell or Molecular Dysfunction|Hospital Course|6092,6100|true|true|false|C4727483|BRAF Gene Rearrangement|positive
Event|Event|Hospital Course|6092,6100|true|false|false|||positive
Finding|Classification|Hospital Course|6092,6100|true|true|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|Hospital Course|6092,6100|true|true|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Event|Event|Hospital Course|6109,6110|true|false|false|||f
Drug|Biomedical or Dental Material|Hospital Course|6113,6120|false|false|false|C1706355|Culture Dose Form|culture
Event|Event|Hospital Course|6113,6120|false|false|false|||culture
Finding|Functional Concept|Hospital Course|6113,6120|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Finding|Idea or Concept|Hospital Course|6113,6120|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Procedure|Laboratory Procedure|Hospital Course|6113,6120|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|culture
Drug|Indicator, Reagent, or Diagnostic Aid|Hospital Course|6123,6133|false|false|false|C0358514|Diagnostic agents|diagnostic
Event|Event|Hospital Course|6123,6133|false|false|false|||diagnostic
Finding|Functional Concept|Hospital Course|6123,6133|false|false|false|C0348026;C1547424|Diagnostic;Location Service Code - Diagnostic|diagnostic
Finding|Intellectual Product|Hospital Course|6123,6133|false|false|false|C0348026;C1547424|Diagnostic;Location Service Code - Diagnostic|diagnostic
Procedure|Diagnostic Procedure|Hospital Course|6123,6133|false|false|false|C0011900;C0430533|Diagnosis;Diagnostic dental procedure|diagnostic
Event|Event|Hospital Course|6134,6138|false|false|false|||para
Finding|Finding|Hospital Course|6134,6138|false|false|false|C0030563|Parity|para
Anatomy|Cell|Hospital Course|6153,6156|true|false|false|C0023516|Leukocytes|WBC
Anatomy|Body Location or Region|Hospital Course|6158,6161|true|false|false|C0230177|Structure of right upper quadrant of abdomen|RUQ
Event|Event|Hospital Course|6176,6184|true|false|false|||thrombus
Finding|Pathologic Function|Hospital Course|6176,6184|true|false|false|C0087086;C0302148|Blood Clot;Thrombus|thrombus
Event|Event|Hospital Course|6187,6196|false|false|false|||Compliant
Finding|Individual Behavior|Hospital Course|6187,6196|false|false|false|C1321605|Compliance behavior|Compliant
Drug|Pharmacologic Substance|Hospital Course|6202,6211|false|false|false|C0012798|Diuretics|diuretics
Event|Event|Hospital Course|6202,6211|false|false|false|||diuretics
Finding|Finding|Hospital Course|6230,6233|true|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Hospital Course|6230,6233|true|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Finding|Hospital Course|6230,6240|true|true|false|C0860871|Sodium decreased|low sodium
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6230,6240|true|true|false|C0012169|Low sodium diet|low sodium
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6230,6245|true|false|false|C0012169|Low sodium diet|low sodium diet
Drug|Biologically Active Substance|Hospital Course|6234,6240|true|true|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|Hospital Course|6234,6240|true|true|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|Hospital Course|6234,6240|true|true|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Event|Event|Hospital Course|6234,6240|true|false|false|||sodium
Finding|Physiologic Function|Hospital Course|6234,6240|true|true|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|Hospital Course|6234,6240|true|true|false|C0337443|Sodium measurement|sodium
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6234,6245|true|false|false|C0301592|Sodium diet|sodium diet
Drug|Food|Hospital Course|6241,6245|true|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|Hospital Course|6241,6245|true|false|false|||diet
Finding|Functional Concept|Hospital Course|6241,6245|true|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|Hospital Course|6241,6245|true|false|false|C0012159|Diet therapy|diet
Drug|Substance|Hospital Course|6250,6255|true|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|6250,6255|true|false|false|C1546638|Fluid Specimen Code|fluid
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6250,6267|true|false|false|C0204700|Fluid restriction|fluid restriction
Event|Event|Hospital Course|6256,6267|false|false|false|||restriction
Finding|Functional Concept|Hospital Course|6256,6267|false|false|false|C0443288|Restricted|restriction
Event|Event|Hospital Course|6277,6286|false|false|false|||discussed
Finding|Finding|Hospital Course|6287,6295|false|false|false|C0332149|Possible|possible
Event|Event|Hospital Course|6296,6300|false|false|false|||TIPS
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6296,6300|false|true|false|C0339897|Transjugular intrahepatic portosystemic shunt (procedure)|TIPS
Event|Event|Hospital Course|6309,6315|false|false|false|||office
Finding|Idea or Concept|Hospital Course|6309,6315|false|false|false|C1549636|Address type - Office|office
Anatomy|Body Location or Region|Hospital Course|6327,6331|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6327,6331|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Hospital Course|6327,6331|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Hospital Course|6327,6331|false|false|false|C0740941|Lung Problem|lung
Disorder|Disease or Syndrome|Hospital Course|6327,6339|false|false|false|C0024115|Lung diseases|lung disease
Disorder|Disease or Syndrome|Hospital Course|6332,6339|false|false|false|C0012634|Disease|disease
Event|Event|Hospital Course|6332,6339|false|false|false|||disease
Finding|Functional Concept|Hospital Course|6350,6357|false|false|false|C4520523|On hold|on hold
Event|Activity|Hospital Course|6353,6357|false|false|false|C1948035|Hold (action)|hold
Finding|Functional Concept|Hospital Course|6353,6357|false|false|false|C1553387;C3853841|Hold - dosing instruction fragment;hold - Data Operation|hold
Finding|Intellectual Product|Hospital Course|6353,6357|false|false|false|C1553387;C3853841|Hold - dosing instruction fragment;hold - Data Operation|hold
Event|Event|Hospital Course|6358,6365|false|false|false|||pending
Finding|Idea or Concept|Hospital Course|6358,6365|false|false|false|C1691786;C1704475|Pending - Allergy Clinical Status;Pending - referral status|pending
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6375,6382|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|Hospital Course|6375,6382|false|false|false|C1314974|Cardiac attachment|cardiac
Procedure|Diagnostic Procedure|Hospital Course|6375,6393|false|false|false|C2024217|cardiac evaluation|cardiac evaluation
Event|Event|Hospital Course|6383,6393|false|false|false|||evaluation
Finding|Idea or Concept|Hospital Course|6383,6393|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|Hospital Course|6383,6393|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Drug|Pharmacologic Substance|Hospital Course|6395,6404|false|false|false|C0012798|Diuretics|Diuretics
Event|Event|Hospital Course|6395,6404|false|false|false|||Diuretics
Event|Event|Hospital Course|6419,6428|false|false|false|||decreased
Disorder|Disease or Syndrome|Hospital Course|6437,6449|false|false|false|C0020625|Hyponatremia|hyponatremia
Event|Event|Hospital Course|6437,6449|false|false|false|||hyponatremia
Event|Event|Hospital Course|6454,6466|false|false|false|||hyperkalemia
Finding|Finding|Hospital Course|6454,6466|false|false|false|C0020461;C5700154|Hyperkalemia;Serum potassium level above reference range|hyperkalemia
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6468,6472|false|false|false|C0675390|ARID1A protein, human|Held
Drug|Biologically Active Substance|Hospital Course|6468,6472|false|false|false|C0675390|ARID1A protein, human|Held
Event|Event|Hospital Course|6468,6472|false|false|false|||Held
Finding|Gene or Genome|Hospital Course|6468,6472|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|Held
Finding|Idea or Concept|Hospital Course|6468,6472|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|Held
Drug|Organic Chemical|Hospital Course|6473,6487|false|false|false|C0037982|spironolactone|spironolactone
Drug|Pharmacologic Substance|Hospital Course|6473,6487|false|false|false|C0037982|spironolactone|spironolactone
Event|Event|Hospital Course|6473,6487|false|false|false|||spironolactone
Event|Event|Hospital Course|6497,6500|false|false|false|||due
Drug|Organic Chemical|Hospital Course|6524,6529|false|false|false|C0699992|Lasix|lasix
Drug|Pharmacologic Substance|Hospital Course|6524,6529|false|false|false|C0699992|Lasix|lasix
Event|Event|Hospital Course|6524,6529|false|false|false|||lasix
Event|Event|Hospital Course|6543,6551|true|false|false|||evidence
Finding|Idea or Concept|Hospital Course|6543,6551|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Hospital Course|6543,6554|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Finding|Finding|Hospital Course|6556,6562|true|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Hospital Course|6556,6562|true|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|Hospital Course|6563,6575|true|false|false|C0020625|Hyponatremia|hyponatremia
Event|Event|Hospital Course|6563,6575|true|false|false|||hyponatremia
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6588,6593|false|false|false|C0022646|Kidney|renal
Disorder|Disease or Syndrome|Hospital Course|6588,6593|false|false|false|C0042075|Urologic Diseases|renal
Disorder|Disease or Syndrome|Hospital Course|6588,6601|false|false|false|C0035078|Kidney Failure|renal failure
Event|Event|Hospital Course|6594,6601|false|false|false|||failure
Finding|Functional Concept|Hospital Course|6594,6601|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|Hospital Course|6594,6601|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|Hospital Course|6594,6601|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Drug|Inorganic Chemical|Hospital Course|6612,6616|false|false|false|C0723457|Stop brand of fluoride|stop
Drug|Pharmacologic Substance|Hospital Course|6612,6616|false|false|false|C0723457|Stop brand of fluoride|stop
Event|Activity|Hospital Course|6612,6616|false|false|false|C1947925|Stop (Instruction Imperative)|stop
Event|Event|Hospital Course|6612,6616|false|false|false|||stop
Finding|Gene or Genome|Hospital Course|6612,6616|false|false|false|C1417022|MAP6 gene|stop
Drug|Pharmacologic Substance|Hospital Course|6618,6627|false|false|false|C0012798|Diuretics|diuretics
Event|Event|Hospital Course|6618,6627|false|false|false|||diuretics
Event|Event|Hospital Course|6631,6638|false|false|false|||present
Finding|Finding|Hospital Course|6631,6638|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|Hospital Course|6631,6638|false|false|false|C0150312;C0449450|Present;Presentation|present
Drug|Indicator, Reagent, or Diagnostic Aid|Hospital Course|6640,6650|true|false|false|C0358514|Diagnostic agents|Diagnostic
Event|Event|Hospital Course|6640,6650|true|false|false|||Diagnostic
Finding|Functional Concept|Hospital Course|6640,6650|true|false|false|C0348026;C1547424|Diagnostic;Location Service Code - Diagnostic|Diagnostic
Finding|Intellectual Product|Hospital Course|6640,6650|true|false|false|C0348026;C1547424|Diagnostic;Location Service Code - Diagnostic|Diagnostic
Procedure|Diagnostic Procedure|Hospital Course|6640,6650|true|false|false|C0011900;C0430533|Diagnosis;Diagnostic dental procedure|Diagnostic
Event|Event|Hospital Course|6651,6663|true|false|false|||paracentesis
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6651,6663|true|false|false|C0034115|Paracentesis|paracentesis
Event|Event|Hospital Course|6664,6672|false|false|false|||negative
Finding|Classification|Hospital Course|6664,6672|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|6664,6672|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|6664,6672|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|Hospital Course|6664,6676|false|false|false|C0205160|Negative|negative for
Disorder|Disease or Syndrome|Hospital Course|6678,6687|true|false|false|C0009450|Communicable Diseases|infection
Event|Event|Hospital Course|6678,6687|true|false|false|||infection
Finding|Pathologic Function|Hospital Course|6678,6687|true|false|false|C3714514|Infection|infection
Finding|Physiologic Function|Hospital Course|6697,6710|false|false|false|C4553020|Total protein metabolic function|total protein
Lab|Laboratory or Test Result|Hospital Course|6697,6710|false|false|false|C1261360|Total protein result|total protein
Procedure|Laboratory Procedure|Hospital Course|6697,6710|false|false|false|C0555903|Total protein measurement|total protein
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6703,6710|false|false|false|C0033684|Proteins|protein
Drug|Biologically Active Substance|Hospital Course|6703,6710|false|false|false|C0033684|Proteins|protein
Event|Event|Hospital Course|6703,6710|false|false|false|||protein
Finding|Conceptual Entity|Hospital Course|6703,6710|false|false|false|C1521746|Protein Info|protein
Procedure|Laboratory Procedure|Hospital Course|6703,6710|false|false|false|C0202202|Protein measurement|protein
Attribute|Clinical Attribute|Hospital Course|6727,6730|false|false|false|C0871470|Systolic Pressure|SBP
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6727,6730|false|false|false|C0085805|Androgen Binding Protein|SBP
Drug|Biologically Active Substance|Hospital Course|6727,6730|false|false|false|C0085805|Androgen Binding Protein|SBP
Event|Event|Hospital Course|6727,6730|false|false|false|||SBP
Finding|Gene or Genome|Hospital Course|6727,6730|false|false|false|C1705296;C3274833|CCHCR1 wt Allele;SHBG wt Allele|SBP
Procedure|Diagnostic Procedure|Hospital Course|6727,6730|false|false|false|C1306620|Systolic blood pressure measurement|SBP
Event|Event|Hospital Course|6731,6742|false|false|false|||prophylaxis
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6731,6742|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Drug|Organic Chemical|Hospital Course|6778,6785|false|false|false|C0591139|Bactrim|Bactrim
Drug|Pharmacologic Substance|Hospital Course|6778,6785|false|false|false|C0591139|Bactrim|Bactrim
Event|Event|Hospital Course|6778,6785|false|false|false|||Bactrim
Disorder|Disease or Syndrome|Hospital Course|6790,6793|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6790,6793|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|Hospital Course|6790,6793|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6790,6793|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|Hospital Course|6790,6793|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|Hospital Course|6790,6793|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|Hospital Course|6790,6793|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|Hospital Course|6790,6793|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|Hospital Course|6790,6793|false|false|false|||PCP
Finding|Gene or Genome|Hospital Course|6790,6793|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|Hospital Course|6790,6793|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6790,6805|false|false|false|C0747314|pcp prophylaxis|PCP prophylaxis
Event|Event|Hospital Course|6794,6805|false|false|false|||prophylaxis
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6794,6805|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Event|Event|Hospital Course|6822,6833|false|false|false|||appropriate
Attribute|Clinical Attribute|Hospital Course|6838,6841|false|true|false|C0871470|Systolic Pressure|SBP
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6838,6841|false|true|false|C0085805|Androgen Binding Protein|SBP
Drug|Biologically Active Substance|Hospital Course|6838,6841|false|true|false|C0085805|Androgen Binding Protein|SBP
Event|Event|Hospital Course|6838,6841|false|false|false|||SBP
Finding|Gene or Genome|Hospital Course|6838,6841|false|true|false|C1705296;C3274833|CCHCR1 wt Allele;SHBG wt Allele|SBP
Procedure|Diagnostic Procedure|Hospital Course|6838,6841|false|true|false|C1306620|Systolic blood pressure measurement|SBP
Event|Event|Hospital Course|6842,6845|false|false|false|||ppx
Finding|Gene or Genome|Hospital Course|6842,6845|false|false|false|C1418850|PPP4C gene|ppx
Finding|Body Substance|Hospital Course|6852,6859|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|6852,6859|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|6852,6859|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|6864,6869|false|false|false|||admit
Procedure|Health Care Activity|Hospital Course|6864,6869|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admit
Event|Event|Hospital Course|6874,6880|false|false|false|||eating
Drug|Food|Hospital Course|6881,6886|false|false|false|C0453577|Pizza|pizza
Event|Event|Hospital Course|6881,6886|false|false|false|||pizza
Drug|Food|Hospital Course|6900,6904|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Drug|Immunologic Factor|Hospital Course|6900,6904|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Drug|Pharmacologic Substance|Hospital Course|6900,6904|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Event|Event|Hospital Course|6900,6904|false|false|false|||food
Event|Event|Hospital Course|6915,6924|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|6915,6924|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Drug|Organic Chemical|Hospital Course|6934,6945|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Drug|Pharmacologic Substance|Hospital Course|6934,6945|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Event|Event|Hospital Course|6934,6945|false|false|false|||therapeutic
Finding|Functional Concept|Hospital Course|6934,6945|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Finding|Intellectual Product|Hospital Course|6934,6945|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6934,6945|false|false|false|C0087111|Therapeutic procedure|therapeutic
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6934,6958|false|false|false|C2057774|Therapeutic abdominal paracentesis|therapeutic paracentesis
Event|Event|Hospital Course|6946,6958|false|false|false|||paracentesis
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6946,6958|false|false|false|C0034115|Paracentesis|paracentesis
Event|Event|Hospital Course|6969,6976|false|false|false|||removed
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6997,7004|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Drug|Biologically Active Substance|Hospital Course|6997,7004|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Drug|Pharmacologic Substance|Hospital Course|6997,7004|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Event|Event|Hospital Course|6997,7004|false|false|false|||albumin
Finding|Gene or Genome|Hospital Course|6997,7004|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|albumin
Finding|Physiologic Function|Hospital Course|6997,7004|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|albumin
Procedure|Laboratory Procedure|Hospital Course|6997,7004|false|false|false|C0201838|Albumin measurement|albumin
Attribute|Clinical Attribute|Hospital Course|7013,7022|false|false|false|C0945766||procedure
Event|Event|Hospital Course|7013,7022|false|false|false|||procedure
Event|Occupational Activity|Hospital Course|7013,7022|false|false|false|C1546467|Act Class - procedure|procedure
Finding|Functional Concept|Hospital Course|7013,7022|false|false|false|C2700391|Procedure (set of actions)|procedure
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7013,7022|false|false|false|C0184661|Interventional procedure|procedure
Event|Event|Hospital Course|7028,7032|false|false|false|||felt
Event|Event|Hospital Course|7033,7037|false|false|false|||much
Finding|Finding|Hospital Course|7033,7037|false|false|false|C4281574|Much|much
Event|Event|Hospital Course|7039,7045|false|false|false|||better
Finding|Idea or Concept|Hospital Course|7039,7045|false|false|false|C1550462|Observation Interpretation - better|better
Event|Event|Hospital Course|7051,7061|false|false|false|||resolution
Finding|Conceptual Entity|Hospital Course|7051,7061|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolution
Finding|Pathologic Function|Hospital Course|7051,7061|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolution
Anatomy|Body Location or Region|Hospital Course|7065,7074|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|Hospital Course|7065,7085|false|false|false|C0232487|Abdominal discomfort|abdominal discomfort
Event|Event|Hospital Course|7075,7085|false|false|false|||discomfort
Finding|Sign or Symptom|Hospital Course|7075,7085|false|false|false|C2364135|Discomfort|discomfort
Finding|Body Substance|Hospital Course|7087,7094|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|7087,7094|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|7087,7094|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|7099,7108|false|false|false|||scheduled
Finding|Functional Concept|Hospital Course|7113,7119|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Event|Event|Hospital Course|7120,7132|false|false|false|||paracentesis
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7120,7132|false|false|false|C0034115|Paracentesis|paracentesis
Event|Event|Hospital Course|7136,7146|false|false|false|||outpatient
Finding|Classification|Hospital Course|7136,7146|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|7136,7146|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Anatomy|Body Location or Region|Hospital Course|7160,7167|false|false|false|C0205054|Hepatic|HEPATIC
Disorder|Disease or Syndrome|Hospital Course|7160,7182|false|false|false|C0019151|Hepatic Encephalopathy|HEPATIC ENCEPHALOPATHY
Disorder|Disease or Syndrome|Hospital Course|7168,7182|false|false|false|C0085584|Encephalopathies|ENCEPHALOPATHY
Event|Event|Hospital Course|7168,7182|false|false|false|||ENCEPHALOPATHY
Event|Event|Hospital Course|7184,7191|false|false|false|||History
Finding|Conceptual Entity|Hospital Course|7184,7191|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|Hospital Course|7184,7191|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|Hospital Course|7184,7191|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|Hospital Course|7184,7194|false|false|false|C0262926|Medical History|History of
Anatomy|Body Location or Region|Hospital Course|7203,7206|false|false|false|C0449198|HEP (body structure)|Hep
Disorder|Disease or Syndrome|Hospital Course|7203,7206|false|false|false|C0162569|Hepatoerythropoietic Porphyria|Hep
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7203,7206|false|false|false|C0540659|EPHB6 protein, human|Hep
Drug|Enzyme|Hospital Course|7203,7206|false|false|false|C0540659|EPHB6 protein, human|Hep
Finding|Gene or Genome|Hospital Course|7203,7206|false|false|false|C0540659;C1414432;C1705569;C2239359;C4723683|DNLZ gene;EPHB6 gene;EPHB6 protein, human;EPHB6 wt Allele, Human;HPSE wt Allele|Hep
Finding|Receptor|Hospital Course|7203,7206|false|false|false|C0540659;C1414432;C1705569;C2239359;C4723683|DNLZ gene;EPHB6 gene;EPHB6 protein, human;EPHB6 wt Allele, Human;HPSE wt Allele|Hep
Drug|Immunologic Factor|Hospital Course|7203,7208|false|false|false|C2148557|hepatitis C vaccine|Hep C
Drug|Pharmacologic Substance|Hospital Course|7203,7208|false|false|false|C2148557|hepatitis C vaccine|Hep C
Disorder|Disease or Syndrome|Hospital Course|7209,7218|false|false|false|C0023890;C1623038|Cirrhosis;Liver Cirrhosis|cirrhosis
Event|Event|Hospital Course|7209,7218|false|false|false|||cirrhosis
Finding|Intellectual Product|Hospital Course|7230,7234|false|false|false|C1547225|Mild Severity of Illness Code|mild
Disorder|Disease or Syndrome|Hospital Course|7235,7249|false|false|false|C0085584|Encephalopathies|encephalopathy
Event|Event|Hospital Course|7235,7249|false|false|false|||encephalopathy
Disorder|Mental or Behavioral Dysfunction|Hospital Course|7251,7265|false|false|false|C0018524|Hallucinations|hallucinations
Event|Event|Hospital Course|7251,7265|false|false|false|||hallucinations
Event|Event|Hospital Course|7270,7283|false|false|false|||forgetfulness
Finding|Sign or Symptom|Hospital Course|7270,7283|false|false|false|C0542476|Forgetful|forgetfulness
Event|Event|Hospital Course|7286,7289|false|false|false|||due
Drug|Pharmacologic Substance|Hospital Course|7293,7303|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Hospital Course|7293,7303|false|false|false|||medication
Finding|Intellectual Product|Hospital Course|7293,7303|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Finding|Finding|Hospital Course|7293,7317|false|false|false|C0746935|Medication Nonadherence|medication noncompliance
Event|Event|Hospital Course|7304,7317|false|false|false|||noncompliance
Event|Event|Hospital Course|7335,7350|true|false|false|||encephalopathic
Event|Event|Hospital Course|7364,7373|true|false|false|||asterixis
Finding|Sign or Symptom|Hospital Course|7364,7373|true|false|false|C0232766|Asterixis|asterixis
Event|Event|Hospital Course|7377,7381|true|false|false|||exam
Finding|Functional Concept|Hospital Course|7377,7381|true|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|Hospital Course|7377,7381|true|false|false|C0582103|Medical Examination|exam
Disorder|Disease or Syndrome|Hospital Course|7383,7393|true|false|false|C0009450|Communicable Diseases|Infectious
Event|Event|Hospital Course|7394,7400|false|false|false|||workup
Event|Event|Hospital Course|7401,7409|false|false|false|||negative
Finding|Classification|Hospital Course|7401,7409|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|7401,7409|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|7401,7409|false|false|false|C5237010|Expression Negative|negative
Procedure|Laboratory Procedure|Hospital Course|7416,7419|false|false|false|C5400981|Fibrinogen to Albumin Ratio Measurement|far
Event|Event|Hospital Course|7421,7429|false|false|false|||Continue
Drug|Organic Chemical|Hospital Course|7430,7439|false|false|false|C0022957|lactulose|lactulose
Drug|Pharmacologic Substance|Hospital Course|7430,7439|false|false|false|C0022957|lactulose|lactulose
Event|Event|Hospital Course|7445,7448|false|false|false|||TID
Event|Event|Hospital Course|7453,7460|false|false|false|||titrate
Procedure|Health Care Activity|Hospital Course|7453,7460|false|false|false|C1883350|Titrate|titrate
Disorder|Disease or Syndrome|Hospital Course|7466,7469|false|false|false|C0006430|Burning Mouth Syndrome|BMs
Event|Event|Hospital Course|7466,7469|false|false|false|||BMs
Event|Event|Hospital Course|7481,7489|false|false|false|||continue
Drug|Organic Chemical|Hospital Course|7490,7499|false|false|false|C0073374|rifaximin|rifaximin
Drug|Pharmacologic Substance|Hospital Course|7490,7499|false|false|false|C0073374|rifaximin|rifaximin
Event|Event|Hospital Course|7500,7505|false|false|false|||550mg
Disorder|Mental or Behavioral Dysfunction|Hospital Course|7506,7509|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7506,7509|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|7506,7509|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|7506,7509|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|7506,7509|false|false|false|C1332410|BID gene|BID
Disorder|Disease or Syndrome|Hospital Course|7516,7528|false|false|false|C0020625|Hyponatremia|HYPONATREMIA
Event|Event|Hospital Course|7516,7528|false|false|false|||HYPONATREMIA
Event|Event|Hospital Course|7540,7549|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|7540,7549|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Gene or Genome|Hospital Course|7565,7568|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Finding|Idea or Concept|Hospital Course|7583,7588|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|Hospital Course|7583,7588|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Gene or Genome|Hospital Course|7589,7592|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|Hospital Course|7594,7600|false|false|false|||Likely
Finding|Finding|Hospital Course|7594,7600|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Idea or Concept|Hospital Course|7594,7600|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Event|Event|Hospital Course|7614,7621|false|false|false|||spacing
Event|Event|Hospital Course|7627,7636|false|false|false|||worsening
Finding|Idea or Concept|Hospital Course|7627,7636|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Disorder|Disease or Syndrome|Hospital Course|7638,7645|false|false|false|C0003962|Ascites|ascites
Event|Event|Hospital Course|7638,7645|false|false|false|||ascites
Finding|Pathologic Function|Hospital Course|7638,7645|false|false|false|C5441966|Peritoneal Effusion|ascites
Drug|Substance|Hospital Course|7650,7655|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|Hospital Course|7650,7655|false|false|false|||fluid
Finding|Intellectual Product|Hospital Course|7650,7655|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Finding|Hospital Course|7650,7664|false|false|false|C0546817;C5848920|Fluid Overload;Hypervolemia (finding)|fluid overload
Finding|Pathologic Function|Hospital Course|7650,7664|false|false|false|C0546817;C5848920|Fluid Overload;Hypervolemia (finding)|fluid overload
Event|Event|Hospital Course|7656,7664|false|false|false|||overload
Drug|Substance|Hospital Course|7671,7676|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|7671,7676|false|false|false|C1546638|Fluid Specimen Code|fluid
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7671,7688|false|false|false|C0204700|Fluid restriction|fluid restriction
Event|Event|Hospital Course|7677,7688|false|false|false|||restriction
Finding|Functional Concept|Hospital Course|7677,7688|false|false|false|C0443288|Restricted|restriction
Finding|Finding|Hospital Course|7690,7693|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Hospital Course|7690,7693|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Drug|Chemical Viewed Structurally|Hospital Course|7694,7698|false|false|false|C0036140;C0037494;C0206136|Salts;Sodium Chloride, Dietary;sodium chloride|salt
Drug|Food|Hospital Course|7694,7698|false|false|false|C0036140;C0037494;C0206136|Salts;Sodium Chloride, Dietary;sodium chloride|salt
Drug|Inorganic Chemical|Hospital Course|7694,7698|false|false|false|C0036140;C0037494;C0206136|Salts;Sodium Chloride, Dietary;sodium chloride|salt
Event|Event|Hospital Course|7694,7698|false|false|false|||salt
Drug|Food|Hospital Course|7700,7704|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|Hospital Course|7700,7704|false|false|false|||diet
Finding|Functional Concept|Hospital Course|7700,7704|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|Hospital Course|7700,7704|false|false|false|C0012159|Diet therapy|diet
Drug|Organic Chemical|Hospital Course|7710,7721|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Drug|Pharmacologic Substance|Hospital Course|7710,7721|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Event|Event|Hospital Course|7710,7721|false|false|false|||therapeutic
Finding|Functional Concept|Hospital Course|7710,7721|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Finding|Intellectual Product|Hospital Course|7710,7721|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7710,7721|false|false|false|C0087111|Therapeutic procedure|therapeutic
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7710,7734|false|false|false|C2057774|Therapeutic abdominal paracentesis|therapeutic paracentesis
Event|Event|Hospital Course|7722,7734|false|false|false|||paracentesis
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7722,7734|false|false|false|C0034115|Paracentesis|paracentesis
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7740,7747|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Drug|Biologically Active Substance|Hospital Course|7740,7747|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Drug|Pharmacologic Substance|Hospital Course|7740,7747|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Event|Event|Hospital Course|7740,7747|false|false|false|||albumin
Finding|Gene or Genome|Hospital Course|7740,7747|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|albumin
Finding|Physiologic Function|Hospital Course|7740,7747|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|albumin
Procedure|Laboratory Procedure|Hospital Course|7740,7747|false|false|false|C0201838|Albumin measurement|albumin
Event|Event|Hospital Course|7748,7759|false|false|false|||replacement
Finding|Functional Concept|Hospital Course|7748,7759|false|false|false|C0559956|Replacement|replacement
Procedure|Health Care Activity|Hospital Course|7748,7759|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7748,7759|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Disorder|Disease or Syndrome|Hospital Course|7764,7773|false|false|false|C0023890;C1623038|Cirrhosis;Liver Cirrhosis|CIRRHOSIS
Event|Event|Hospital Course|7764,7773|false|false|false|||CIRRHOSIS
Disorder|Disease or Syndrome|Hospital Course|7775,7784|false|false|false|C0019158;C0019159|Hepatitis;Hepatitis A|HEPATITIS
Finding|Intellectual Product|Hospital Course|7788,7792|false|false|false|C3826979;C4049616|Model for End Stage Liver Disease Clinical Classification;Model for End-Stage Liver Disease|MELD
Attribute|Clinical Attribute|Hospital Course|7788,7798|false|false|false|C1715987||MELD score
Finding|Intellectual Product|Hospital Course|7788,7798|false|false|false|C3826979|Model for End-Stage Liver Disease|MELD score
Procedure|Laboratory Procedure|Hospital Course|7788,7798|false|false|false|C4048785|Model for end stage liver disease score|MELD score
Event|Event|Hospital Course|7793,7798|false|false|false|||score
Finding|Finding|Hospital Course|7793,7798|false|false|false|C0449820|Score|score
Event|Event|Hospital Course|7809,7814|false|false|false|||Child
Finding|Idea or Concept|Hospital Course|7809,7814|false|false|false|C1546495|Relationship - Child|Child
Finding|Classification|Hospital Course|7822,7827|false|false|false|C0008902;C0008903;C0456387;C0489477;C1705943|Class;Classification;LOINC class types;Taxonomic;Taxonomic Class|class
Finding|Functional Concept|Hospital Course|7822,7827|false|false|false|C0008902;C0008903;C0456387;C0489477;C1705943|Class;Classification;LOINC class types;Taxonomic;Taxonomic Class|class
Finding|Intellectual Product|Hospital Course|7822,7827|false|false|false|C0008902;C0008903;C0456387;C0489477;C1705943|Class;Classification;LOINC class types;Taxonomic;Taxonomic Class|class
Event|Event|Hospital Course|7838,7847|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|7838,7847|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|Hospital Course|7853,7866|false|false|false|||decompensated
Disorder|Disease or Syndrome|Hospital Course|7874,7881|false|false|false|C0003962|Ascites|ascites
Event|Event|Hospital Course|7874,7881|false|false|false|||ascites
Finding|Pathologic Function|Hospital Course|7874,7881|false|false|false|C5441966|Peritoneal Effusion|ascites
Disorder|Disease or Syndrome|Hospital Course|7884,7893|false|false|false|C0019158;C0019159|Hepatitis;Hepatitis A|Hepatitis
Event|Event|Hospital Course|7884,7893|false|false|false|||Hepatitis
Disorder|Disease or Syndrome|Hospital Course|7884,7895|false|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|Hepatitis C
Disorder|Virus|Hospital Course|7884,7895|false|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|Hepatitis C
Event|Event|Hospital Course|7896,7904|false|false|false|||genotype
Procedure|Laboratory Procedure|Hospital Course|7896,7904|false|false|false|C1285573|Genotype determination|genotype
Event|Event|Hospital Course|7905,7909|false|false|false|||IIIB
Event|Event|Hospital Course|7919,7927|false|false|false|||starting
Finding|Body Substance|Hospital Course|7946,7953|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|7946,7953|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|7946,7953|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|7973,7982|false|false|false|||insurance
Finding|Idea or Concept|Hospital Course|7973,7982|false|false|false|C0021672|Insurance|insurance
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7983,7990|false|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|Hospital Course|7983,7990|false|false|false|C1951340|Process Pharmacologic Substance|process
Event|Event|Hospital Course|7983,7990|false|false|false|||process
Finding|Functional Concept|Hospital Course|7983,7990|false|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|Hospital Course|7983,7990|false|false|false|C1522240|Process|process
Event|Event|Hospital Course|7995,8002|false|false|false|||started
Event|Event|Hospital Course|8010,8016|false|false|false|||office
Finding|Idea or Concept|Hospital Course|8010,8016|false|false|false|C1549636|Address type - Office|office
Event|Event|Hospital Course|8021,8028|true|false|false|||history
Finding|Conceptual Entity|Hospital Course|8021,8028|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|8021,8028|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|8021,8028|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|8021,8031|true|false|false|C0262926|Medical History|history of
Event|Event|Hospital Course|8032,8035|true|false|false|||EGD
Procedure|Diagnostic Procedure|Hospital Course|8032,8035|true|false|false|C0079304|Esophagogastroduodenoscopy|EGD
Event|Event|Hospital Course|8038,8043|true|false|false|||needs
Event|Event|Hospital Course|8052,8062|false|false|false|||outpatient
Finding|Classification|Hospital Course|8052,8062|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|8052,8062|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Disorder|Disease or Syndrome|Hospital Course|8067,8074|false|false|false|C0042345|Varicosity|varices
Event|Event|Hospital Course|8075,8084|false|false|false|||screening
Finding|Finding|Hospital Course|8075,8084|false|false|false|C0220909;C1305399;C1409616|Aspects of disease screening;Screening - procedure intent;Special screening finding|screening
Finding|Functional Concept|Hospital Course|8075,8084|false|false|false|C0220909;C1305399;C1409616|Aspects of disease screening;Screening - procedure intent;Special screening finding|screening
Procedure|Diagnostic Procedure|Hospital Course|8075,8084|false|false|false|C0199230;C0220908;C1698960;C1710031;C1710032|Disease Screening;Screening;Screening for cancer;Screening procedure;research subject screening|screening
Procedure|Health Care Activity|Hospital Course|8075,8084|false|false|false|C0199230;C0220908;C1698960;C1710031;C1710032|Disease Screening;Screening;Screening for cancer;Screening procedure;research subject screening|screening
Procedure|Research Activity|Hospital Course|8075,8084|false|false|false|C0199230;C0220908;C1698960;C1710031;C1710032|Disease Screening;Screening;Screening for cancer;Screening procedure;research subject screening|screening
Event|Event|Hospital Course|8092,8101|false|false|false|||NUTRITION
Finding|Finding|Hospital Course|8092,8101|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|NUTRITION
Finding|Intellectual Product|Hospital Course|8092,8101|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|NUTRITION
Finding|Organism Function|Hospital Course|8092,8101|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|NUTRITION
Procedure|Research Activity|Hospital Course|8092,8101|false|false|false|C0600072;C1521729|Feeding and dietary regimes;Nutritional Study|NUTRITION
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8092,8101|false|false|false|C0600072;C1521729|Feeding and dietary regimes;Nutritional Study|NUTRITION
Event|Event|Hospital Course|8120,8129|false|false|false|||compliant
Finding|Individual Behavior|Hospital Course|8120,8129|false|false|false|C1321605|Compliance behavior|compliant
Finding|Finding|Hospital Course|8135,8138|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Hospital Course|8135,8138|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8135,8148|false|false|false|C0012169|Low sodium diet|low salt diet
Drug|Chemical Viewed Structurally|Hospital Course|8139,8143|false|false|false|C0036140;C0037494;C0206136|Salts;Sodium Chloride, Dietary;sodium chloride|salt
Drug|Food|Hospital Course|8139,8143|false|false|false|C0036140;C0037494;C0206136|Salts;Sodium Chloride, Dietary;sodium chloride|salt
Drug|Inorganic Chemical|Hospital Course|8139,8143|false|false|false|C0036140;C0037494;C0206136|Salts;Sodium Chloride, Dietary;sodium chloride|salt
Drug|Food|Hospital Course|8144,8148|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|Hospital Course|8144,8148|false|false|false|||diet
Finding|Functional Concept|Hospital Course|8144,8148|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|Hospital Course|8144,8148|false|false|false|C0012159|Diet therapy|diet
Finding|Intellectual Product|Hospital Course|8150,8154|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|Poor
Anatomy|Body Space or Junction|Hospital Course|8156,8160|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|8156,8160|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|8156,8160|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|8156,8160|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Finding|Hospital Course|8156,8167|false|false|false|C2137071|Oral intake|oral intake
Event|Event|Hospital Course|8161,8167|false|false|false|||intake
Finding|Functional Concept|Hospital Course|8161,8167|false|false|false|C1512806|Intake|intake
Procedure|Health Care Activity|Hospital Course|8161,8167|false|false|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|intake
Finding|Finding|Hospital Course|8169,8172|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|Low
Finding|Intellectual Product|Hospital Course|8169,8172|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|Low
Finding|Finding|Hospital Course|8169,8180|false|false|false|C0860864|Albumin below reference range|Low albumin
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8173,8180|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Drug|Biologically Active Substance|Hospital Course|8173,8180|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Drug|Pharmacologic Substance|Hospital Course|8173,8180|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Event|Event|Hospital Course|8173,8180|false|false|false|||albumin
Finding|Gene or Genome|Hospital Course|8173,8180|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|albumin
Finding|Physiologic Function|Hospital Course|8173,8180|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|albumin
Procedure|Laboratory Procedure|Hospital Course|8173,8180|false|false|false|C0201838|Albumin measurement|albumin
Event|Event|Hospital Course|8188,8197|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|8188,8197|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|Hospital Course|8199,8202|false|false|false|||Met
Event|Event|Hospital Course|8208,8217|false|false|false|||nutrition
Finding|Finding|Hospital Course|8208,8217|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|nutrition
Finding|Intellectual Product|Hospital Course|8208,8217|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|nutrition
Finding|Organism Function|Hospital Course|8208,8217|false|false|false|C0392209;C0518896;C1442959|Nutrition (function);Nutrition outcomes;Nutritional status|nutrition
Procedure|Research Activity|Hospital Course|8208,8217|false|false|false|C0600072;C1521729|Feeding and dietary regimes;Nutritional Study|nutrition
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8208,8217|false|false|false|C0600072;C1521729|Feeding and dietary regimes;Nutritional Study|nutrition
Disorder|Disease or Syndrome|Hospital Course|8224,8236|false|false|false|C0005779|Blood Coagulation Disorders|COAGULOPATHY
Event|Event|Hospital Course|8224,8236|false|false|false|||COAGULOPATHY
Attribute|Clinical Attribute|Hospital Course|8238,8241|false|false|false|C0368980|Coagulation tissue factor induced.INR|INR
Event|Event|Hospital Course|8238,8241|false|false|false|||INR
Procedure|Laboratory Procedure|Hospital Course|8238,8241|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8238,8241|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Finding|Gene or Genome|Hospital Course|8256,8259|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|Hospital Course|8264,8272|true|false|false|||evidence
Finding|Idea or Concept|Hospital Course|8264,8272|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Hospital Course|8264,8275|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Event|Event|Hospital Course|8284,8292|true|false|false|||bleeding
Finding|Pathologic Function|Hospital Course|8284,8292|true|false|false|C0019080|Hemorrhage|bleeding
Finding|Finding|Hospital Course|8294,8303|false|false|false|C4036115|Very mild|Very mild
Finding|Intellectual Product|Hospital Course|8299,8303|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Finding|Hospital Course|8299,8320|false|false|false|C1856453|Mild thrombocytopenia|mild thrombocytopenia
Disorder|Disease or Syndrome|Hospital Course|8304,8320|false|false|false|C0040034|Thrombocytopenia|thrombocytopenia
Event|Event|Hospital Course|8304,8320|false|false|false|||thrombocytopenia
Finding|Finding|Hospital Course|8304,8320|false|false|false|C0392386|Decreased platelet count|thrombocytopenia
Disorder|Disease or Syndrome|Hospital Course|8342,8345|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Disorder|Virus|Hospital Course|8342,8345|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Drug|Immunologic Factor|Hospital Course|8342,8345|false|false|false|C0086413|HIV Vaccine|HIV
Drug|Pharmacologic Substance|Hospital Course|8342,8345|false|false|false|C0086413|HIV Vaccine|HIV
Event|Event|Hospital Course|8342,8345|false|false|false|||HIV
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8359,8362|false|false|false|C0003323;C4048280|CD4 Antigens;T-Cell Surface Glycoprotein CD4, human|CD4
Drug|Biologically Active Substance|Hospital Course|8359,8362|false|false|false|C0003323;C4048280|CD4 Antigens;T-Cell Surface Glycoprotein CD4, human|CD4
Drug|Immunologic Factor|Hospital Course|8359,8362|false|false|false|C0003323;C4048280|CD4 Antigens;T-Cell Surface Glycoprotein CD4, human|CD4
Event|Event|Hospital Course|8359,8362|false|false|false|||CD4
Finding|Gene or Genome|Hospital Course|8359,8362|false|false|false|C0003323;C1332714|CD4 Antigens;CD4 gene|CD4
Finding|Receptor|Hospital Course|8359,8362|false|false|false|C0003323;C1332714|CD4 Antigens;CD4 gene|CD4
Event|Event|Hospital Course|8371,8376|false|false|false|||HAART
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8371,8376|false|false|false|C0887947|Antiretroviral Therapy, Highly Active|HAART
Event|Event|Hospital Course|8397,8405|true|false|false|||provider
Finding|Functional Concept|Hospital Course|8397,8405|true|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|provider
Finding|Intellectual Product|Hospital Course|8397,8405|true|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|provider
Event|Event|Hospital Course|8407,8415|false|false|false|||Continue
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Hospital Course|8416,8423|false|false|false|C1528494|Truvada|Truvada
Drug|Pharmacologic Substance|Hospital Course|8416,8423|false|false|false|C1528494|Truvada|Truvada
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Hospital Course|8428,8437|false|false|false|C1967563|Isentress|Isentress
Drug|Pharmacologic Substance|Hospital Course|8428,8437|false|false|false|C1967563|Isentress|Isentress
Event|Event|Hospital Course|8428,8437|false|false|false|||Isentress
Drug|Organic Chemical|Hospital Course|8439,8446|false|false|false|C0591139|Bactrim|Bactrim
Drug|Pharmacologic Substance|Hospital Course|8439,8446|false|false|false|C0591139|Bactrim|Bactrim
Drug|Organic Chemical|Hospital Course|8439,8449|false|false|false|C1154231|Bactrim DS|Bactrim DS
Drug|Pharmacologic Substance|Hospital Course|8439,8449|false|false|false|C1154231|Bactrim DS|Bactrim DS
Disorder|Disease or Syndrome|Hospital Course|8461,8464|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8461,8464|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|Hospital Course|8461,8464|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8461,8464|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|Hospital Course|8461,8464|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|Hospital Course|8461,8464|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|Hospital Course|8461,8464|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|Hospital Course|8461,8464|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|Hospital Course|8461,8464|false|false|false|||PCP
Finding|Gene or Genome|Hospital Course|8461,8464|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|Hospital Course|8461,8464|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|Hospital Course|8476,8486|false|false|false|||outpatient
Finding|Classification|Hospital Course|8476,8486|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|8476,8486|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Activity|Hospital Course|8490,8501|false|false|false|C0003629|Appointments|appointment
Event|Event|Hospital Course|8490,8501|false|false|false|||appointment
Disorder|Disease or Syndrome|Hospital Course|8507,8511|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|8507,8511|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|8507,8511|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|8507,8511|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|Hospital Course|8513,8519|false|false|false|||Stable
Finding|Intellectual Product|Hospital Course|8513,8519|false|false|false|C1547311|Patient Condition Code - Stable|Stable
Event|Event|Hospital Course|8521,8527|false|false|false|||States
Event|Event|Hospital Course|8551,8555|false|false|false|||home
Finding|Idea or Concept|Hospital Course|8551,8555|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|8551,8555|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|8551,8555|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|8564,8571|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Drug|Pharmacologic Substance|Hospital Course|8564,8571|false|false|false|C1310585|Comfort brand of hydroxyethyl cellulose|comfort
Event|Event|Hospital Course|8564,8571|false|false|false|||comfort
Finding|Mental Process|Hospital Course|8564,8571|false|false|false|C1331418|Comfort|comfort
Anatomy|Body Location or Region|Hospital Course|8590,8599|false|false|false|C0000726|Abdomen|abdominal
Event|Event|Hospital Course|8600,8610|false|false|false|||distentiom
Event|Event|Hospital Course|8622,8626|false|false|false|||home
Finding|Idea or Concept|Hospital Course|8622,8626|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|8622,8626|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|8622,8626|false|false|false|C1553498|home health encounter|home
Disorder|Disease or Syndrome|Hospital Course|8628,8632|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|8628,8632|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|8628,8632|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|8628,8632|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|Hospital Course|8633,8637|false|false|false|C3280240|MICROCEPHALY, EPILEPSY, AND DIABETES SYNDROME 1|meds
Event|Event|Hospital Course|8633,8637|false|false|false|||meds
Finding|Intellectual Product|Hospital Course|8633,8637|false|false|false|C4284232|Medications|meds
Event|Event|Hospital Course|8642,8646|false|false|false|||home
Finding|Idea or Concept|Hospital Course|8642,8646|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|8642,8646|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|8642,8646|false|false|false|C1553498|home health encounter|home
Event|Event|Hospital Course|8653,8659|false|false|false|||needed
Finding|Idea or Concept|Hospital Course|8664,8676|false|false|false|C1548597|Marketing basis - Transitional|Transitional
Event|Event|Hospital Course|8677,8683|false|false|false|||Issues
Drug|Organic Chemical|Hospital Course|8701,8715|false|false|false|C0037982|spironolactone|spironolactone
Drug|Pharmacologic Substance|Hospital Course|8701,8715|false|false|false|C0037982|spironolactone|spironolactone
Event|Event|Hospital Course|8701,8715|false|false|false|||spironolactone
Drug|Biologically Active Substance|Hospital Course|8729,8738|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Element, Ion, or Isotope|Hospital Course|8729,8738|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Food|Hospital Course|8729,8738|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Inorganic Chemical|Hospital Course|8729,8738|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Pharmacologic Substance|Hospital Course|8729,8738|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Event|Event|Hospital Course|8729,8738|false|false|false|||potassium
Finding|Physiologic Function|Hospital Course|8729,8738|false|false|false|C4553027|Potassium metabolic function|potassium
Procedure|Laboratory Procedure|Hospital Course|8729,8738|false|false|false|C0202194|Potassium measurement|potassium
Event|Event|Hospital Course|8741,8750|false|false|false|||Increased
Drug|Organic Chemical|Hospital Course|8751,8761|false|false|false|C0016860|furosemide|furosemide
Drug|Pharmacologic Substance|Hospital Course|8751,8761|false|false|false|C0016860|furosemide|furosemide
Event|Event|Hospital Course|8751,8761|false|false|false|||furosemide
Event|Event|Hospital Course|8785,8792|false|false|false|||recheck
Drug|Inorganic Chemical|Hospital Course|8793,8805|false|false|false|C0013832;C3536863|Electrolyte [EPC];Electrolytes|electrolytes
Drug|Pharmacologic Substance|Hospital Course|8793,8805|false|false|false|C0013832;C3536863|Electrolyte [EPC];Electrolytes|electrolytes
Event|Event|Hospital Course|8793,8805|false|false|false|||electrolytes
Finding|Idea or Concept|Hospital Course|8809,8813|false|false|false|C1552851|next - HtmlLinkType|next
Event|Event|Hospital Course|8814,8819|false|false|false|||visit
Finding|Social Behavior|Hospital Course|8814,8819|false|false|false|C0545082|Visit|visit
Event|Event|Hospital Course|8826,8838|false|false|false|||paracentesis
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8826,8838|false|false|false|C0034115|Paracentesis|paracentesis
Event|Event|Hospital Course|8854,8861|false|false|false|||removed
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8879,8886|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Drug|Biologically Active Substance|Hospital Course|8879,8886|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Drug|Pharmacologic Substance|Hospital Course|8879,8886|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Event|Event|Hospital Course|8879,8886|false|false|false|||albumin
Finding|Gene or Genome|Hospital Course|8879,8886|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|albumin
Finding|Physiologic Function|Hospital Course|8879,8886|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|albumin
Procedure|Laboratory Procedure|Hospital Course|8879,8886|false|false|false|C0201838|Albumin measurement|albumin
Event|Event|Hospital Course|8895,8905|false|false|false|||outpatient
Finding|Classification|Hospital Course|8895,8905|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|8895,8905|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|Hospital Course|8909,8917|false|false|false|||provider
Finding|Functional Concept|Hospital Course|8909,8917|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|provider
Finding|Intellectual Product|Hospital Course|8909,8917|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|provider
Event|Event|Hospital Course|8944,8956|false|false|false|||paracentesis
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8944,8956|false|false|false|C0034115|Paracentesis|paracentesis
Attribute|Clinical Attribute|Hospital Course|8959,8970|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|8959,8970|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|8959,8970|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|8959,8970|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|8959,8983|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|8974,8983|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|8974,8983|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|Hospital Course|9002,9012|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Hospital Course|9002,9012|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|Hospital Course|9002,9017|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|Hospital Course|9013,9017|false|false|false|||list
Finding|Intellectual Product|Hospital Course|9013,9017|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|Hospital Course|9021,9029|false|false|false|||accurate
Drug|Organic Chemical|Hospital Course|9034,9042|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Hospital Course|9034,9042|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Hospital Course|9034,9042|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|Hospital Course|9034,9042|false|false|false|||complete
Finding|Functional Concept|Hospital Course|9034,9042|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|9034,9042|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|Hospital Course|9047,9056|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|Hospital Course|9047,9056|false|false|false|C0001927|albuterol|Albuterol
Finding|Functional Concept|Hospital Course|9057,9064|false|false|false|C4319647|Inhaler (unit of presentation)|Inhaler
Finding|Gene or Genome|Hospital Course|9079,9082|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|9083,9091|false|false|false|||wheezing
Finding|Sign or Symptom|Hospital Course|9083,9091|false|false|false|C0043144|Wheezing|wheezing
Event|Event|Hospital Course|9093,9096|false|false|false|||SOB
Finding|Sign or Symptom|Hospital Course|9093,9096|false|false|false|C0013404|Dyspnea|SOB
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Hospital Course|9106,9113|false|false|false|C1528494|Truvada|Truvada
Drug|Pharmacologic Substance|Hospital Course|9106,9113|false|false|false|C1528494|Truvada|Truvada
Drug|Biomedical or Dental Material|Hospital Course|9117,9120|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|Hospital Course|9117,9120|false|false|false|||TAB
Drug|Organic Chemical|Hospital Course|9134,9144|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|Hospital Course|9134,9144|false|false|false|C0016860|furosemide|Furosemide
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Hospital Course|9164,9175|false|false|false|C1871526|raltegravir|Raltegravir
Drug|Pharmacologic Substance|Hospital Course|9164,9175|false|false|false|C1871526|raltegravir|Raltegravir
Event|Event|Hospital Course|9164,9175|false|false|false|||Raltegravir
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9186,9189|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9186,9189|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9186,9189|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|9186,9189|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|9186,9189|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|9194,9208|false|false|false|C0037982|spironolactone|Spironolactone
Drug|Pharmacologic Substance|Hospital Course|9194,9208|false|false|false|C0037982|spironolactone|Spironolactone
Drug|Organic Chemical|Hospital Course|9228,9241|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|9228,9241|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Hospital Course|9228,9241|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|9228,9241|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|Hospital Course|9256,9259|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|9260,9264|false|false|false|C2598155||pain
Event|Event|Hospital Course|9260,9264|false|false|false|||pain
Finding|Functional Concept|Hospital Course|9260,9264|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|9260,9264|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|9265,9270|false|false|false|||fever
Finding|Finding|Hospital Course|9265,9270|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|Hospital Course|9265,9270|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Drug|Organic Chemical|Hospital Course|9275,9285|false|false|false|C0213771|tiotropium|Tiotropium
Drug|Pharmacologic Substance|Hospital Course|9275,9285|false|false|false|C0213771|tiotropium|Tiotropium
Event|Event|Hospital Course|9275,9285|false|false|false|||Tiotropium
Drug|Organic Chemical|Hospital Course|9275,9293|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Pharmacologic Substance|Hospital Course|9275,9293|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Inorganic Chemical|Hospital Course|9286,9293|false|false|false|C0006222|Bromides|Bromide
Event|Event|Hospital Course|9286,9293|false|false|false|||Bromide
Procedure|Laboratory Procedure|Hospital Course|9286,9293|false|false|false|C0202341|Bromides measurement|Bromide
Disorder|Congenital Abnormality|Hospital Course|9296,9299|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|CAP
Drug|Biomedical or Dental Material|Hospital Course|9296,9299|false|false|false|C0006935|capsule (pharmacologic)|CAP
Event|Event|Hospital Course|9296,9299|false|false|false|||CAP
Finding|Gene or Genome|Hospital Course|9296,9299|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|CAP
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9296,9299|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|CAP
Drug|Organic Chemical|Hospital Course|9313,9322|false|false|false|C0073374|rifaximin|Rifaximin
Drug|Pharmacologic Substance|Hospital Course|9313,9322|false|false|false|C0073374|rifaximin|Rifaximin
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9333,9336|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9333,9336|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9333,9336|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|9333,9336|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|9333,9336|false|false|false|C1332410|BID gene|BID
Drug|Biologically Active Substance|Hospital Course|9341,9348|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|Hospital Course|9341,9348|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|Hospital Course|9341,9348|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|Hospital Course|9341,9348|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|Hospital Course|9341,9348|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|Hospital Course|9341,9348|false|false|false|||Calcium
Finding|Physiologic Function|Hospital Course|9341,9348|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|Hospital Course|9341,9348|false|false|false|C0201925|Calcium measurement|Calcium
Drug|Inorganic Chemical|Hospital Course|9341,9358|false|false|false|C0006681|calcium carbonate|Calcium Carbonate
Drug|Pharmacologic Substance|Hospital Course|9341,9358|false|false|false|C0006681|calcium carbonate|Calcium Carbonate
Drug|Element, Ion, or Isotope|Hospital Course|9349,9358|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|Carbonate
Drug|Organic Chemical|Hospital Course|9349,9358|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|Carbonate
Drug|Pharmacologic Substance|Hospital Course|9349,9358|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|Carbonate
Event|Event|Hospital Course|9349,9358|false|false|false|||Carbonate
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9370,9373|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9370,9373|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9370,9373|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|9370,9373|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|9370,9373|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|9379,9388|false|false|false|C0022957|lactulose|Lactulose
Drug|Pharmacologic Substance|Hospital Course|9379,9388|false|false|false|C0022957|lactulose|Lactulose
Event|Event|Hospital Course|9398,9401|false|false|false|||TID
Drug|Antibiotic|Hospital Course|9417,9429|false|false|false|C0041041|trimethoprim|Trimethoprim
Drug|Organic Chemical|Hospital Course|9417,9429|false|false|false|C0041041|trimethoprim|Trimethoprim
Drug|Biomedical or Dental Material|Hospital Course|9435,9438|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|Hospital Course|9435,9438|false|false|false|||TAB
Event|Event|Hospital Course|9452,9461|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|9452,9461|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|9452,9461|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|9452,9461|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|9452,9461|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|9452,9473|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|9462,9473|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|9462,9473|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|9462,9473|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|9462,9473|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|9478,9491|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|9478,9491|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Hospital Course|9478,9491|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|9478,9491|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|Hospital Course|9506,9509|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|9510,9514|false|false|false|C2598155||pain
Event|Event|Hospital Course|9510,9514|false|false|false|||pain
Finding|Functional Concept|Hospital Course|9510,9514|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|9510,9514|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|9515,9520|false|false|false|||fever
Finding|Finding|Hospital Course|9515,9520|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|Hospital Course|9515,9520|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Drug|Organic Chemical|Hospital Course|9525,9534|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|Hospital Course|9525,9534|false|false|false|C0001927|albuterol|Albuterol
Finding|Functional Concept|Hospital Course|9535,9542|false|false|false|C4319647|Inhaler (unit of presentation)|Inhaler
Finding|Gene or Genome|Hospital Course|9557,9560|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|9561,9569|false|false|false|||wheezing
Finding|Sign or Symptom|Hospital Course|9561,9569|false|false|false|C0043144|Wheezing|wheezing
Event|Event|Hospital Course|9571,9574|false|false|false|||SOB
Finding|Sign or Symptom|Hospital Course|9571,9574|false|false|false|C0013404|Dyspnea|SOB
Drug|Biologically Active Substance|Hospital Course|9579,9586|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|Hospital Course|9579,9586|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|Hospital Course|9579,9586|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|Hospital Course|9579,9586|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|Hospital Course|9579,9586|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|Hospital Course|9579,9586|false|false|false|||Calcium
Finding|Physiologic Function|Hospital Course|9579,9586|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|Hospital Course|9579,9586|false|false|false|C0201925|Calcium measurement|Calcium
Drug|Inorganic Chemical|Hospital Course|9579,9596|false|false|false|C0006681|calcium carbonate|Calcium Carbonate
Drug|Pharmacologic Substance|Hospital Course|9579,9596|false|false|false|C0006681|calcium carbonate|Calcium Carbonate
Drug|Element, Ion, or Isotope|Hospital Course|9587,9596|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|Carbonate
Drug|Organic Chemical|Hospital Course|9587,9596|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|Carbonate
Drug|Pharmacologic Substance|Hospital Course|9587,9596|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|Carbonate
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9608,9611|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9608,9611|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9608,9611|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|9608,9611|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|9608,9611|false|false|false|C1332410|BID gene|BID
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Hospital Course|9621,9628|false|false|false|C1528494|Truvada|Truvada
Drug|Pharmacologic Substance|Hospital Course|9621,9628|false|false|false|C1528494|Truvada|Truvada
Drug|Biomedical or Dental Material|Hospital Course|9632,9635|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|Hospital Course|9632,9635|false|false|false|||TAB
Drug|Organic Chemical|Hospital Course|9649,9659|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|Hospital Course|9649,9659|false|false|false|C0016860|furosemide|Furosemide
Drug|Organic Chemical|Hospital Course|9679,9688|false|false|false|C0022957|lactulose|Lactulose
Drug|Pharmacologic Substance|Hospital Course|9679,9688|false|false|false|C0022957|lactulose|Lactulose
Event|Event|Hospital Course|9698,9701|false|false|false|||TID
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Hospital Course|9706,9717|false|false|false|C1871526|raltegravir|Raltegravir
Drug|Pharmacologic Substance|Hospital Course|9706,9717|false|false|false|C1871526|raltegravir|Raltegravir
Event|Event|Hospital Course|9706,9717|false|false|false|||Raltegravir
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9728,9731|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9728,9731|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9728,9731|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|9728,9731|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|9728,9731|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|9736,9745|false|false|false|C0073374|rifaximin|Rifaximin
Drug|Pharmacologic Substance|Hospital Course|9736,9745|false|false|false|C0073374|rifaximin|Rifaximin
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9756,9759|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9756,9759|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9756,9759|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|9756,9759|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|9756,9759|false|false|false|C1332410|BID gene|BID
Drug|Antibiotic|Hospital Course|9774,9786|false|false|false|C0041041|trimethoprim|Trimethoprim
Drug|Organic Chemical|Hospital Course|9774,9786|false|false|false|C0041041|trimethoprim|Trimethoprim
Drug|Biomedical or Dental Material|Hospital Course|9792,9795|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|Hospital Course|9792,9795|false|false|false|||TAB
Drug|Organic Chemical|Hospital Course|9810,9820|false|false|false|C0213771|tiotropium|Tiotropium
Drug|Pharmacologic Substance|Hospital Course|9810,9820|false|false|false|C0213771|tiotropium|Tiotropium
Event|Event|Hospital Course|9810,9820|false|false|false|||Tiotropium
Drug|Organic Chemical|Hospital Course|9810,9828|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Pharmacologic Substance|Hospital Course|9810,9828|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Inorganic Chemical|Hospital Course|9821,9828|false|false|false|C0006222|Bromides|Bromide
Event|Event|Hospital Course|9821,9828|false|false|false|||Bromide
Procedure|Laboratory Procedure|Hospital Course|9821,9828|false|false|false|C0202341|Bromides measurement|Bromide
Disorder|Congenital Abnormality|Hospital Course|9831,9834|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|CAP
Drug|Biomedical or Dental Material|Hospital Course|9831,9834|false|false|false|C0006935|capsule (pharmacologic)|CAP
Event|Event|Hospital Course|9831,9834|false|false|false|||CAP
Finding|Gene or Genome|Hospital Course|9831,9834|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|CAP
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9831,9834|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|CAP
Event|Event|Hospital Course|9848,9857|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|9848,9857|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|9848,9857|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|9848,9857|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|9848,9857|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|9848,9869|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|9848,9869|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|9858,9869|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|9858,9869|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|9858,9869|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|Hospital Course|9871,9875|false|false|false|||Home
Finding|Idea or Concept|Hospital Course|9871,9875|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|9871,9875|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|9871,9875|false|false|false|C1553498|home health encounter|Home
Event|Event|Hospital Course|9878,9887|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|9878,9887|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|9878,9887|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|9878,9887|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|9878,9887|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|9878,9897|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|9888,9897|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|9888,9897|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|9888,9897|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|9888,9897|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|9888,9897|false|false|false|C0011900|Diagnosis|Diagnosis
Drug|Pharmacologic Substance|Hospital Course|9909,9917|false|false|false|C0012798;C5399719|Diuretic [APC];Diuretics|diuretic
Event|Event|Hospital Course|9909,9917|false|false|false|||diuretic
Finding|Functional Concept|Hospital Course|9918,9928|false|false|false|C0205269|Unresponsive to Treatment|refractory
Finding|Finding|Hospital Course|9918,9936|false|false|false|C3532188|Refractory ascites|refractory ascites
Disorder|Disease or Syndrome|Hospital Course|9929,9936|false|false|false|C0003962|Ascites|ascites
Event|Event|Hospital Course|9929,9936|false|false|false|||ascites
Finding|Pathologic Function|Hospital Course|9929,9936|false|false|false|C5441966|Peritoneal Effusion|ascites
Disorder|Neoplastic Process|Hospital Course|9937,9946|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Event|Event|Hospital Course|9937,9946|false|false|false|||Secondary
Finding|Functional Concept|Hospital Course|9937,9946|false|false|false|C1522484|metastatic qualifier|Secondary
Disorder|Disease or Syndrome|Hospital Course|9948,9951|false|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|HCV
Disorder|Virus|Hospital Course|9948,9951|false|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|HCV
Event|Event|Hospital Course|9948,9951|false|false|false|||HCV
Disorder|Disease or Syndrome|Hospital Course|9952,9961|false|false|false|C0023890;C1623038|Cirrhosis;Liver Cirrhosis|cirrhosis
Event|Event|Hospital Course|9952,9961|false|false|false|||cirrhosis
Disorder|Disease or Syndrome|Hospital Course|9963,9966|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Disorder|Virus|Hospital Course|9963,9966|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Drug|Immunologic Factor|Hospital Course|9963,9966|false|false|false|C0086413|HIV Vaccine|HIV
Drug|Pharmacologic Substance|Hospital Course|9963,9966|false|false|false|C0086413|HIV Vaccine|HIV
Event|Event|Hospital Course|9963,9966|false|false|false|||HIV
Disorder|Disease or Syndrome|Hospital Course|9968,9980|false|false|false|C0020625|Hyponatremia|hyponatremia
Event|Event|Hospital Course|9968,9980|false|false|false|||hyponatremia
Disorder|Disease or Syndrome|Hospital Course|9982,9986|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|9982,9986|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|9982,9986|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|9982,9986|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Mental Process|Discharge Condition|10011,10017|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|10011,10024|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|10011,10024|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|10018,10024|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|10018,10024|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|10026,10031|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|10026,10031|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|10036,10044|false|false|false|||coherent
Finding|Finding|Discharge Condition|10036,10044|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|10046,10051|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|10046,10068|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|10046,10068|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|10055,10068|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|10055,10068|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|10055,10068|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|10070,10075|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|10070,10075|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|10070,10075|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|10070,10075|false|false|false|||Alert
Finding|Finding|Discharge Condition|10070,10075|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|10070,10075|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|10070,10075|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|10080,10091|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|10080,10091|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|10093,10101|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|10093,10101|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|10093,10101|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|10102,10108|false|false|false|C5889824||Status
Event|Event|Discharge Condition|10102,10108|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|10102,10108|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|10110,10120|false|false|false|||Ambulatory
Finding|Functional Concept|Discharge Condition|10110,10120|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|10110,10120|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|10110,10120|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|10110,10120|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|10123,10134|false|false|false|||Independent
Finding|Finding|Discharge Condition|10123,10134|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Condition|10123,10134|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Gene or Genome|Discharge Instructions|10163,10167|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|Discharge Instructions|10184,10192|false|false|false|||pleasure
Finding|Intellectual Product|Discharge Instructions|10184,10192|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|Discharge Instructions|10184,10192|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|Discharge Instructions|10201,10205|false|false|false|C1947933|care activity|care
Event|Event|Discharge Instructions|10201,10205|false|false|false|||care
Finding|Finding|Discharge Instructions|10201,10205|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|10201,10205|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|10201,10208|false|false|false|C1555558|care of - AddressPartType|care of
Event|Event|Discharge Instructions|10235,10243|false|false|false|||admitted
Anatomy|Body Location or Region|Discharge Instructions|10249,10258|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|Discharge Instructions|10249,10267|false|false|false|C0235318|Fullness abdominal|abdominal fullness
Event|Event|Discharge Instructions|10259,10267|false|false|false|||fullness
Attribute|Clinical Attribute|Discharge Instructions|10273,10277|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|10273,10277|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|10273,10277|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|10273,10277|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Disorder|Disease or Syndrome|Discharge Instructions|10288,10295|false|false|false|C0003962|Ascites|ascites
Event|Event|Discharge Instructions|10288,10295|false|false|false|||ascites
Finding|Pathologic Function|Discharge Instructions|10288,10295|false|false|false|C5441966|Peritoneal Effusion|ascites
Drug|Indicator, Reagent, or Diagnostic Aid|Discharge Instructions|10307,10317|false|false|false|C0358514|Diagnostic agents|diagnostic
Event|Event|Discharge Instructions|10307,10317|false|false|false|||diagnostic
Finding|Functional Concept|Discharge Instructions|10307,10317|false|false|false|C0348026;C1547424|Diagnostic;Location Service Code - Diagnostic|diagnostic
Finding|Intellectual Product|Discharge Instructions|10307,10317|false|false|false|C0348026;C1547424|Diagnostic;Location Service Code - Diagnostic|diagnostic
Procedure|Diagnostic Procedure|Discharge Instructions|10307,10317|false|false|false|C0011900;C0430533|Diagnosis;Diagnostic dental procedure|diagnostic
Finding|Functional Concept|Discharge Instructions|10307,10333|false|false|false|C5817574|Combined diagnostic and therapeutic intent|diagnostic and therapeutic
Drug|Organic Chemical|Discharge Instructions|10322,10333|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Drug|Pharmacologic Substance|Discharge Instructions|10322,10333|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Event|Event|Discharge Instructions|10322,10333|false|false|false|||therapeutic
Finding|Functional Concept|Discharge Instructions|10322,10333|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Finding|Intellectual Product|Discharge Instructions|10322,10333|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10322,10333|false|false|false|C0087111|Therapeutic procedure|therapeutic
Event|Event|Discharge Instructions|10335,10347|false|false|false|||paracentesis
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10335,10347|false|false|false|C0034115|Paracentesis|paracentesis
Event|Event|Discharge Instructions|10359,10366|false|false|false|||removed
Drug|Organic Chemical|Discharge Instructions|10373,10387|false|false|false|C0037982|spironolactone|spironolactone
Drug|Pharmacologic Substance|Discharge Instructions|10373,10387|false|false|false|C0037982|spironolactone|spironolactone
Event|Event|Discharge Instructions|10373,10387|false|false|false|||spironolactone
Event|Event|Discharge Instructions|10393,10405|false|false|false|||discontinued
Drug|Biologically Active Substance|Discharge Instructions|10419,10428|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Element, Ion, or Isotope|Discharge Instructions|10419,10428|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Food|Discharge Instructions|10419,10428|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Inorganic Chemical|Discharge Instructions|10419,10428|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Pharmacologic Substance|Discharge Instructions|10419,10428|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Event|Event|Discharge Instructions|10419,10428|false|false|false|||potassium
Finding|Physiologic Function|Discharge Instructions|10419,10428|false|false|false|C4553027|Potassium metabolic function|potassium
Procedure|Laboratory Procedure|Discharge Instructions|10419,10428|false|false|false|C0202194|Potassium measurement|potassium
Event|Event|Discharge Instructions|10433,10437|false|false|false|||high
Finding|Finding|Discharge Instructions|10433,10437|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|Discharge Instructions|10433,10437|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|Discharge Instructions|10433,10437|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Drug|Organic Chemical|Discharge Instructions|10444,10449|false|false|false|C0699992|Lasix|lasix
Drug|Pharmacologic Substance|Discharge Instructions|10444,10449|false|false|false|C0699992|Lasix|lasix
Event|Event|Discharge Instructions|10444,10449|false|false|false|||lasix
Event|Event|Discharge Instructions|10455,10464|false|false|false|||increased
Event|Event|Discharge Instructions|10488,10497|false|false|false|||scheduled
Event|Event|Discharge Instructions|10511,10523|false|false|false|||paracentesis
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10511,10523|false|false|false|C0034115|Paracentesis|paracentesis
Event|Activity|Discharge Instructions|10551,10563|false|false|false|C0003629|Appointments|appointments
Event|Event|Discharge Instructions|10551,10563|false|false|false|||appointments
Finding|Idea or Concept|Discharge Instructions|10569,10572|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Discharge Instructions|10569,10572|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Discharge Instructions|10582,10586|false|false|false|||call
Event|Event|Discharge Instructions|10599,10603|false|false|false|||find
Finding|Finding|Discharge Instructions|10612,10616|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Discharge Instructions|10612,10616|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Discharge Instructions|10612,10616|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|Discharge Instructions|10624,10636|false|false|false|||paracentesis
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10624,10636|false|false|false|C0034115|Paracentesis|paracentesis
Event|Event|Discharge Instructions|10646,10654|false|false|false|||continue
Event|Event|Discharge Instructions|10658,10664|false|false|false|||follow
Finding|Finding|Discharge Instructions|10667,10670|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Discharge Instructions|10667,10670|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Finding|Discharge Instructions|10667,10677|false|false|false|C0860871|Sodium decreased|low sodium
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10667,10677|false|false|false|C0012169|Low sodium diet|low sodium
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10667,10682|false|false|false|C0012169|Low sodium diet|low sodium diet
Drug|Biologically Active Substance|Discharge Instructions|10671,10677|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|Discharge Instructions|10671,10677|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|Discharge Instructions|10671,10677|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Event|Event|Discharge Instructions|10671,10677|false|false|false|||sodium
Finding|Physiologic Function|Discharge Instructions|10671,10677|false|false|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|Discharge Instructions|10671,10677|false|false|false|C0337443|Sodium measurement|sodium
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10671,10682|false|false|false|C0301592|Sodium diet|sodium diet
Drug|Food|Discharge Instructions|10678,10682|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|Discharge Instructions|10678,10682|false|false|false|||diet
Finding|Functional Concept|Discharge Instructions|10678,10682|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|Discharge Instructions|10678,10682|false|false|false|C0012159|Diet therapy|diet
Drug|Substance|Discharge Instructions|10687,10692|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|Discharge Instructions|10687,10692|false|false|false|||fluid
Finding|Intellectual Product|Discharge Instructions|10687,10692|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|Discharge Instructions|10694,10705|false|false|false|||restriction
Finding|Functional Concept|Discharge Instructions|10694,10705|false|false|false|C0443288|Restricted|restriction
Event|Event|Discharge Instructions|10718,10722|false|false|false|||call
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|10728,10733|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Discharge Instructions|10728,10733|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Discharge Instructions|10728,10733|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Discharge Instructions|10728,10733|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Discharge Instructions|10728,10733|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Discharge Instructions|10728,10733|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Finding|Finding|Discharge Instructions|10728,10733|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Discharge Instructions|10728,10733|false|false|false|C0872387|Procedures on liver|liver
Event|Event|Discharge Instructions|10734,10740|false|false|false|||doctor
Finding|Intellectual Product|Discharge Instructions|10734,10740|false|false|false|C2348314|Doctor - Title|doctor
Event|Event|Discharge Instructions|10744,10750|false|false|false|||return
Finding|Finding|Discharge Instructions|10759,10768|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Idea or Concept|Discharge Instructions|10759,10768|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Intellectual Product|Discharge Instructions|10759,10768|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Pathologic Function|Discharge Instructions|10759,10768|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Phenomenon|Phenomenon or Process|Discharge Instructions|10759,10768|false|false|false|C0013956|Emergency Situation|emergency
Procedure|Health Care Activity|Discharge Instructions|10759,10768|false|false|false|C1553500|emergency encounter|emergency
Finding|Idea or Concept|Discharge Instructions|10759,10773|false|false|false|C1546435|Encounter Referral Source - emergency room|emergency room
Anatomy|Body Location or Region|Discharge Instructions|10786,10795|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|Discharge Instructions|10786,10800|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|Discharge Instructions|10796,10800|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|10796,10800|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|10796,10800|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|10796,10800|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Discharge Instructions|10802,10807|false|false|false|||fever
Finding|Finding|Discharge Instructions|10802,10807|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|Discharge Instructions|10802,10807|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|Discharge Instructions|10809,10815|false|false|false|||chills
Finding|Sign or Symptom|Discharge Instructions|10809,10815|false|false|false|C0085593|Chills|chills
Disorder|Mental or Behavioral Dysfunction|Discharge Instructions|10818,10827|false|false|false|C0009676|Confusion|confusion
Event|Event|Discharge Instructions|10818,10827|false|false|false|||confusion
Finding|Finding|Discharge Instructions|10818,10827|false|false|false|C0683369|Clouded consciousness|confusion
Event|Event|Discharge Instructions|10849,10857|false|false|false|||symptoms
Finding|Functional Concept|Discharge Instructions|10849,10857|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Discharge Instructions|10849,10857|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Functional Concept|Discharge Instructions|10880,10887|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|Discharge Instructions|10880,10887|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|Discharge Instructions|10880,10887|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|Discharge Instructions|10880,10887|false|false|false|C0199168|Medical service|medical
Procedure|Health Care Activity|Discharge Instructions|10895,10903|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|10904,10916|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|10904,10916|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|10904,10916|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

