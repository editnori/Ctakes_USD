CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|true|false||Unit
null|Unit device|Device|true|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|true|false||Unit
null|Unit of Measure|LabModifier|true|false||Unit
null|Unit|LabModifier|true|false||Unit
null|Enzyme Unit|LabModifier|true|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Urology|Title|false|false||UROLOGYnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Known|Modifier|true|false||Knownnull|Hypersensitivity|Finding|true|false||Allergiesnull|null|Attribute|true|false||Allergiesnull|Adverse reaction to drug|Finding|true|false||Adverse Drug Reactionsnull|Adverse reaction to drug|Finding|true|false||Drug Reactionsnull|Pharmaceutical Preparations|Drug|true|false||Drug
null|Pharmacologic Substance|Drug|true|false||Drugnull|Drug problem|Finding|true|false||Drugnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Chief complaint (finding)|Finding|false|false||Chief Complaintnull|Complaint (finding)|Finding|false|false||Complaintnull|null|Attribute|false|false||Complaintnull|Abdominal Pain|Finding|false|false||Abdominal painnull|Abdomen|Anatomy|false|false||Abdominalnull|Abdominal (qualifier value)|Modifier|false|false||Abdominalnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Distention|Finding|false|false||distention
null|Pathological Dilatation|Finding|false|false||distentionnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Interventional Radiology Procedure|Procedure|false|false||Interventional radiologynull|Interventional radiology|Title|false|false||Interventional radiologynull|interventional (invasive) radiology|Procedure|false|false||Interventional
null|Interventional procedure|Procedure|false|false||Interventionalnull|radiology referral type|Finding|false|false||radiology
null|Radiology Section ID|Finding|false|false||radiology
null|Encounter due to radiological examination|Finding|false|false||radiologynull|Radiology studies|Procedure|false|false||radiology
null|Diagnostic radiologic examination|Procedure|false|false||radiology
null|Radiographic imaging procedure|Procedure|false|false||radiologynull|Radiology Specialty|Title|false|false||radiologynull|Clinical act of insertion|Procedure|false|false||placement
null|Implantation procedure|Procedure|false|false||placement
null|null|Procedure|false|false||placementnull|Placement|Modifier|false|false||placementnull|Abdominal Abscess|Disorder|false|false||abdominal abscessnull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Abscess|Disorder|false|false||abscessnull|null|Finding|false|false||abscessnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|History of present illness (finding)|Finding|false|false||History of Present Illnessnull|null|Attribute|false|false||History of Present Illnessnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Present illness|Finding|false|false||Present Illnessnull|Present|Finding|false|false||Present
null|Presentation|Finding|false|false||Presentnull|Illness (finding)|Finding|false|false||Illnessnull|Muscle (organ)|Anatomy|false|false||muscle
null|Muscle Tissue|Anatomy|false|false||musclenull|Carcinoma of urinary bladder, invasive|Disorder|false|false||invasive bladder cancernull|Invasive|Modifier|false|false||invasivenull|Malignant neoplasm of urinary bladder|Disorder|false|false||bladder cancer
null|Carcinoma of bladder|Disorder|false|false||bladder cancer
null|Bladder Neoplasm|Disorder|false|false||bladder cancernull|Neoplasm of uncertain or unknown behavior of bladder|Disorder|false|false||bladder
null|Benign neoplasm of bladder|Disorder|false|false||bladder
null|Carcinoma in situ of bladder|Disorder|false|false||bladdernull|Procedures on bladder|Procedure|false|false||bladdernull|Urinary Bladder|Anatomy|false|false||bladdernull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Abdominal Pain|Finding|false|false||abdominal painnull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Pathological Dilatation|Finding|false|false||distension
null|Distention|Finding|false|false||distensionnull|Nearly|Modifier|false|false||nearlynull|day|Time|false|false||daysnull|X-Ray Computed Tomography|Procedure|false|false||CT scannull|Radionuclide Imaging|Procedure|false|false||scan
null|Scanning|Procedure|false|false||scannull|Dilated loops|Finding|false|false||dilated loopsnull|Dilated|Finding|false|false||dilatednull|null|Device|false|false||loopsnull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false||air
null|AIRN gene|Finding|false|false||air
null|AI/RHEUM|Finding|false|false||airnull|Liquid substance|Drug|true|false||fluidsnull|Mouse Body Fluid or Substance|Finding|true|false||fluidsnull|Fluid Therapy|Procedure|true|false||fluidsnull|Abdomen>Small bowel|Anatomy|true|false||small bowel
null|Intestines, Small|Anatomy|true|false||small bowelnull|Small|LabModifier|true|false||smallnull|Intestines|Anatomy|true|false||bowelnull|Obvious|Modifier|true|false||obviousnull|Transition Point|Finding|true|false||transition pointnull|Transition Mutation|Disorder|true|false||transitionnull|Transition (action)|Event|true|false||transitionnull|Point|Modifier|true|false||pointnull|point - UnitsOfMeasure|LabModifier|true|false||pointnull|Leukocytosis|Disorder|false|false||leukocytosisnull|Blood leukocyte number above reference range|Finding|false|false||leukocytosisnull|Small bowel obstruction|Disorder|false|false||small bowel obstructionnull|Abdomen>Small bowel|Anatomy|false|false||small bowel
null|Intestines, Small|Anatomy|false|false||small bowelnull|Small|LabModifier|false|false||smallnull|Intestinal Obstruction|Disorder|false|false||bowel obstructionnull|Intestines|Anatomy|false|false||bowelnull|Obstruction|Finding|false|false||obstructionnull|Intestinal obstruction co-occurrent and due to decreased peristalsis|Disorder|false|false||ileus
null|Ileus|Disorder|false|false||ileusnull|Providing presence (regime/therapy)|Procedure|false|false||presencenull|Presence (property)|Modifier|false|false||presencenull|Leukocytosis|Disorder|false|false||leukocytosisnull|Blood leukocyte number above reference range|Finding|false|false||leukocytosisnull|Ventricular Fibrillation, Paroxysmal Familial, 1|Disorder|false|false||IVFnull|SCN5A wt Allele|Finding|false|false||IVF
null|SCN5A gene|Finding|false|false||IVFnull|Fertilization in Vitro|Procedure|false|false||IVF
null|Assisted Reproductive Technologies|Procedure|false|false||IVFnull|Structure of interventricular foramen|Anatomy|false|false||IVFnull|Intestines|Anatomy|false|false||bowelnull|REST protein, human|Drug|false|false||rest
null|REST protein, human|Drug|false|false||restnull|REST gene|Finding|false|false||rest
null|site-specific telomere resolvase activity|Finding|false|false||rest
null|Rest|Finding|false|false||restnull|Decompression - action (qualifier value)|Finding|false|false||decompressionnull|Decompression|Procedure|false|false||decompression
null|Decompressive incision|Procedure|false|false||decompressionnull|external decompression|Phenomenon|false|false||decompressionnull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Hypertensive disease|Disorder|false|false||Hypertensionnull|Cholecystectomy, Laparoscopic|Procedure|false|false||laparoscopic cholecystectomynull|Laparoscopy|Procedure|false|false||laparoscopicnull|Laparoscopic approach|Modifier|false|false||laparoscopicnull|Cholecystectomy procedure|Procedure|false|false||cholecystectomynull|Structure of left knee region|Anatomy|false|false||left knee
null|Structure of left knee|Anatomy|false|false||left kneenull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Examination of knee joint|Procedure|false|false||kneenull|Knee region structure|Anatomy|false|false||knee
null|Knee|Anatomy|false|false||knee
null|Lower extremity>Knee|Anatomy|false|false||knee
null|Knee joint|Anatomy|false|false||kneenull|Replacement|Finding|false|false||replacementnull|Replacement - supply|Procedure|false|false||replacement
null|Surgical Replantation|Procedure|false|false||replacementnull|year|Time|false|false||yearsnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|Laminectomy|Procedure|false|false||laminectomynull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|Vaginal Dosage Form|Drug|false|false||vaginalnull|Vaginal Route of Administration|Finding|false|false||vaginal
null|Vaginal (intended site)|Finding|false|false||vaginalnull|Vagina|Anatomy|false|false||vaginalnull|Vaginal|Modifier|false|false||vaginalnull|Robot Device|Device|false|false||Robot
null|null|Device|false|false||Robotnull|Laparoscopy|Procedure|false|false||laparoscopicnull|Laparoscopic approach|Modifier|false|false||laparoscopicnull|Bilateral|Modifier|false|false||bilateralnull|Pelvic lymph node group|Anatomy|false|false||pelvic lymph nodenull|Pelvis|Anatomy|false|false||pelvicnull|lymph nodes|Anatomy|false|false||lymph nodenull|Lymph|Finding|false|false||lymphnull|Dissecting hemorrhage|Finding|false|false||dissectionnull|Tissue Dissection|Procedure|false|false||dissectionnull|Robot Device|Device|false|false||Robot
null|null|Device|false|false||Robotnull|Consent Type - Hysterectomy|Finding|false|false||hysterectomynull|Hysterectomy|Procedure|false|false||hysterectomynull|Bilateral oophorectomy|Procedure|false|false||bilateral oophorectomynull|Bilateral|Modifier|false|false||bilateralnull|Ovariectomy|Procedure|false|false||oophorectomynull|Enlarged uterus|Finding|false|false||large uterusnull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|Neoplasm of uncertain or unknown behavior of uterus|Disorder|false|false||uterus
null|Uterine Diseases|Disorder|false|false||uterusnull|examination of uterus|Procedure|false|false||uterusnull|Pelvis>Uterus|Anatomy|false|false||uterus
null|Mouse Uterus|Anatomy|false|false||uterus
null|Uterus|Anatomy|false|false||uterusnull|Greater Than|LabModifier|false|false||greater thannull|Greater|LabModifier|false|false||greaternull|gram|LabModifier|false|false||gramsnull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|Fibroid Tumor|Disorder|false|false||fibroidnull|Laparoscopic radical cystectomy|Procedure|false|false||Laparoscopic radical cystectomynull|Laparoscopy|Procedure|false|false||Laparoscopicnull|Laparoscopic approach|Modifier|false|false||Laparoscopicnull|Complete cystectomy|Procedure|false|false||radical cystectomynull|Radicals (chemistry)|Drug|false|false||radicalnull|Radical (qualifier value)|Modifier|false|false||radicalnull|Cystectomy|Procedure|false|false||cystectomynull|Adenohypophyseal Diseases|Disorder|false|false||anteriornull|Anterior|Modifier|false|false||anteriornull|Vaginectomy|Procedure|false|false||vaginectomynull|Reconstruction of vagina|Procedure|false|false||vaginal reconstructionnull|Vaginal Dosage Form|Drug|false|false||vaginalnull|Vaginal Route of Administration|Finding|false|false||vaginal
null|Vaginal (intended site)|Finding|false|false||vaginalnull|Vagina|Anatomy|false|false||vaginalnull|Vaginal|Modifier|false|false||vaginalnull|Optical Image Reconstruction|Procedure|false|false||reconstruction
null|Reconstructive Surgical Procedures|Procedure|false|false||reconstructionnull|Social and personal history|Finding|false|false||Social History
null|Social History|Finding|false|false||Social Historynull|Social|Finding|false|false||Socialnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Family Medical History|Finding|false|false||Family Historynull|Entity Name Part Type - family|Finding|false|false||Family
null|Last Name|Finding|false|false||Family
null|Living Arrangement - Family|Finding|false|false||Family
null|Family (taxonomic)|Finding|false|false||Family
null|Family Collection|Finding|false|false||Familynull|Family|Subject|false|false||Familynull|History of present illness (finding)|Finding|false|true||History
null|History of previous events|Finding|false|true||History
null|Historical aspects qualifier|Finding|false|true||History
null|Medical History|Finding|false|true||History
null|Concept History|Finding|false|true||Historynull|History|Subject|false|false||Historynull|Negative|Finding|false|false||Negative fornull|Rh Negative Blood Group|Finding|false|false||Negative
null|Negative|Finding|false|false||Negative
null|Negative Finding|Finding|false|false||Negativenull|Expression Negative|Lab|false|false||Negativenull|Negative - qualifier|Modifier|false|false||Negative
null|Negative Charge|Modifier|false|false||Negativenull|Negative Number|LabModifier|false|false||Negativenull|Malignant neoplasm of urinary bladder|Disorder|true|false||bladder CAnull|Neoplasm of uncertain or unknown behavior of bladder|Disorder|true|false||bladder
null|Benign neoplasm of bladder|Disorder|true|false||bladder
null|Carcinoma in situ of bladder|Disorder|true|false||bladdernull|Procedures on bladder|Procedure|true|false||bladdernull|Urinary Bladder|Anatomy|true|false||bladdernull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|Abdomen soft|Finding|false|false||Abdomen softnull|Malignant neoplasm of abdomen|Disorder|false|false||Abdomennull|Abdomen problem|Finding|false|false||Abdomennull|Abdomen|Anatomy|false|false||Abdomen
null|Abdominal Cavity|Anatomy|false|false||Abdomennull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|Tender|Modifier|false|false||tendernull|Surgical wound|Disorder|false|false||incisionnull|Surgical incisions|Procedure|false|false||incisionnull|Cranial incision point|Anatomy|false|false||incisionnull|Surgical wound|Disorder|false|false||Incisionnull|Surgical incisions|Procedure|false|false||Incisionnull|Cranial incision point|Anatomy|false|false||Incisionnull|Surgical Stoma|Anatomy|false|false||Stomanull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Color of urine|Finding|false|false||Urine colornull|Portion of urine|Finding|false|false||Urine
null|null|Finding|false|false||Urine
null|Urine|Finding|false|false||Urine
null|In Urine|Finding|false|false||Urine
null|Urine specimen|Finding|false|false||Urinenull|color additive|Drug|false|false||color
null|Coloring Excipient|Drug|false|false||colornull|color - solid dosage form|Modifier|false|false||color
null|Color|Modifier|false|false||colornull|Color quantity|LabModifier|false|false||colornull|Yellow color|Modifier|false|false||yellownull|Bilateral|Modifier|false|false||Bilateralnull|Lower Extremity|Anatomy|false|false||lower extremitiesnull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|Feels warm|Finding|false|false||warmnull|warming process|Phenomenon|false|false||warmnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Pain in calf|Finding|true|false||calf painnull|Structure of calf of leg|Anatomy|true|false||calf
null|null|Anatomy|true|false||calfnull|Cattle calf (organism)|Entity|true|false||calfnull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Deep palpation|Procedure|true|false||deep palpationnull|Deep Resection Margin|Attribute|true|false||deepnull|Deep (qualifier value)|Modifier|true|false||deepnull|Palpation|Procedure|true|false||palpationnull|Bilateral|Modifier|false|false||Bilateralnull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|2+ pitting edema|Finding|false|false||2+ pitting edemanull|Pitting edema|Finding|false|false||pitting edemanull|Pitting|Finding|false|false||pittingnull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Erythema|Disorder|true|false||erythemanull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Pigtail Drain|Device|false|false||Pigtail drainnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Dressing Dosage Form|Drug|false|false||dressingnull|null|Finding|false|false||dressing
null|Ability to dress|Finding|false|false||dressingnull|Dressing patient (procedure)|Procedure|false|false||dressing
null|Dressing of skin or wound|Procedure|false|false||dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Bands|Device|false|false||Bandsnull|Lymph|Finding|false|false||Lymphsnull|Monos|Drug|false|false||Monos
null|Mono-S|Drug|false|false||Monos
null|Monos|Drug|false|false||Monosnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||Eos
null|Familial eosinophilia|Disorder|false|false||Eosnull|PRSS33 gene|Finding|false|false||Eos
null|IKZF4 gene|Finding|false|false||Eosnull|Eos <Loriini>|Entity|false|false||Eosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||ASTnull|Atypical Spitz Nevus|Disorder|false|false||ASTnull|SLC17A5 wt Allele|Finding|false|false||AST
null|SLC17A5 gene|Finding|false|false||AST
null|GOT1 gene|Finding|false|false||ASTnull|Asterion|Anatomy|false|false||ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Alkaline Phosphatase|Drug|false|false||AlkPhos
null|Alkaline Phosphatase|Drug|false|false||AlkPhosnull|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood albumin|Procedure|false|false||BLOOD Albuminnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Albumin|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumin|Drug|false|false||Albuminnull|Albumin metabolic function|Finding|false|false||Albumin
null|ALB gene|Finding|false|false||Albuminnull|Albumin measurement|Procedure|false|false||Albuminnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Iron Drug Class|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||Ironnull|Iron measurement|Procedure|false|false||Ironnull|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Thyrotropin-Releasing Hormone, human|Drug|false|false||TRF
null|IL5 protein, human|Drug|false|false||TRF
null|IL5 protein, human|Drug|false|false||TRF
null|thyrotropin-releasing hormone|Drug|false|false||TRF
null|thyrotropin-releasing hormone|Drug|false|false||TRF
null|thyrotropin-releasing hormone|Drug|false|false||TRF
null|Tocotrienol-rich Fraction|Drug|false|false||TRF
null|Thyrotropin-Releasing Hormone, human|Drug|false|false||TRFnull|TERF1 wt Allele|Finding|false|false||TRF
null|TERF1 gene|Finding|false|false||TRF
null|IL5 gene|Finding|false|false||TRFnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|lactate in blood (lab test)|Procedure|false|false||BLOOD Lactatenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|lactate|Drug|false|false||Lactate
null|lactate|Drug|false|false||Lactate
null|Lactates|Drug|false|false||Lactatenull|Lactic acid measurement|Procedure|false|false||Lactatenull|Ascites|Disorder|false|false||ASCITESnull|Peritoneal Effusion|Finding|false|false||ASCITESnull|amylase|Drug|false|false||Amylase
null|amylase|Drug|false|false||Amylase
null|amylase|Drug|false|false||Amylasenull|Amylase measurement|Procedure|false|false||Amylasenull|lipase|Drug|false|false||Lipase
null|lipase|Drug|false|false||Lipase
null|lipase|Drug|false|false||Lipasenull|Lipase measurement|Procedure|false|false||Lipasenull|Body Fluids|Finding|false|false||BODY FLUIDnull|Document Body|Finding|false|false||BODYnull|Structure of body of caudate nucleus|Anatomy|false|false||BODY
null|Human body structure|Anatomy|false|false||BODY
null|Body structure|Anatomy|false|false||BODY
null|Adult human body|Anatomy|false|false||BODY
null|Whole body|Anatomy|false|false||BODYnull|Human body|Subject|false|false||BODYnull|fluid - substance|Drug|false|false||FLUID
null|Liquid substance|Drug|false|false||FLUIDnull|Fluid Specimen Code|Finding|false|false||FLUIDnull|Fluid behavior|Modifier|false|false||FLUIDnull|Blood culture|Procedure|false|false||BLOOD CULTUREnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Final report|Finding|false|false||FINAL REPORTnull|Diagnosis Type - Final|Finding|false|false||FINALnull|Final|Time|false|false||FINALnull|End-stage|Modifier|false|false||FINALnull|Report (document)|Finding|false|false||REPORTnull|Reporting|Procedure|false|false||REPORTnull|null|Attribute|false|false||REPORTnull|Blood culture|Procedure|false|false||Blood Culturenull|Blood and lymphatic system disorders|Disorder|false|false||Bloodnull|peripheral blood|Finding|false|false||Blood
null|Blood|Finding|false|false||Blood
null|In Blood|Finding|false|false||Bloodnull|Culture Dose Form|Drug|false|false||Culturenull|Culture (Anthropological)|Finding|false|false||Culture
null|Cultural aspects|Finding|false|false||Culturenull|Microbial culture (procedure)|Procedure|false|false||Culture
null|Laboratory culture|Procedure|false|false||Culturenull|Extended Priority Codes - Routine|Finding|false|false||Routine
null|Report priority - Routine|Finding|false|false||Routine
null|Admission Type - Routine|Finding|false|false||Routine
null|Level of Care - Routine|Finding|false|false||Routine
null|Processing priority - Routine|Finding|false|false||Routine
null|Referral priority - Routine|Finding|false|false||Routinenull|Routine coag|Procedure|false|false||Routinenull|Priority - Routine|Time|false|false||Routinenull|Routine|Modifier|false|false||Routinenull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Citrobacter koseri|Entity|false|false||CITROBACTER KOSERInull|Citrobacter|Entity|false|false||CITROBACTERnull|Diagnosis Type - Final|Finding|false|false||FINALnull|Final|Time|false|false||FINALnull|End-stage|Modifier|false|false||FINALnull|Antimicrobial susceptibility|Finding|false|false||SENSITIVITIESnull|Antimicrobial susceptibility|Finding|false|false||SENSITIVITIESnull|methyl isocyanate|Drug|false|false||MIC
null|methyl isocyanate|Drug|false|false||MICnull|Ductal Carcinoma In Situ with Microinvasion|Disorder|false|false||MICnull|cisplatin/ifosfamide/mitomycin protocol|Procedure|false|false||MIC
null|Minimum Inhibitory Concentration Test|Procedure|false|false||MICnull|Micmac language|Entity|false|false||MICnull|Microgram per Milliliter|LabModifier|false|false||MCG/MLnull|microgram|LabModifier|false|false||MCGnull|per milliliter|LabModifier|false|false||/MLnull|Citrobacter koseri|Entity|false|false||CITROBACTER KOSERInull|Citrobacter|Entity|false|false||CITROBACTERnull|cefepime|Drug|false|false||CEFEPIME
null|cefepime|Drug|false|false||CEFEPIMEnull|ceftazidime|Drug|false|false||CEFTAZIDIME
null|ceftazidime|Drug|false|false||CEFTAZIDIMEnull|ceftriaxone|Drug|false|false||CEFTRIAXONE
null|ceftriaxone|Drug|false|false||CEFTRIAXONEnull|ciprofloxacin|Drug|false|false||CIPROFLOXACIN
null|ciprofloxacin|Drug|false|false||CIPROFLOXACINnull|gentamicin|Drug|false|false||GENTAMICIN
null|gentamicin|Drug|false|false||GENTAMICINnull|Gentamicin measurement|Procedure|false|false||GENTAMICINnull|INJECTION, MEROPENEM, 100 MG ADMINISTERED|Drug|false|false||MEROPENEM
null|meropenem|Drug|false|false||MEROPENEM
null|meropenem|Drug|false|false||MEROPENEMnull|piperacillin|Drug|false|false||PIPERACILLIN
null|piperacillin|Drug|false|false||PIPERACILLINnull|tazobactam|Drug|false|false||TAZO
null|tazobactam|Drug|false|false||TAZOnull|tobramycin|Drug|false|false||TOBRAMYCIN
null|tobramycin|Drug|false|false||TOBRAMYCINnull|Tobramycin measurement|Procedure|false|false||TOBRAMYCINnull|trimethoprim|Drug|false|false||TRIMETHOPRIM
null|trimethoprim|Drug|false|false||TRIMETHOPRIMnull|sulfa|Drug|false|false||SULFAnull|Aerobic|Modifier|false|false||Aerobicnull|null|Device|false|false||Bottlenull|Bottle (unit of presentation)|LabModifier|false|false||Bottle
null|Bottle Dosing Unit|LabModifier|false|false||Bottlenull|Gram's stain|Drug|false|false||Gram Stain
null|Gram's stain|Drug|false|false||Gram Stainnull|Bacterial stain, routine|Procedure|false|false||Gram Stainnull|gram|LabModifier|false|false||Gramnull|Stains|Drug|false|false||Stainnull|Staining method|Procedure|false|false||Stainnull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Gram-negative bacillus|Entity|false|false||GRAM NEGATIVE RODnull|gram|LabModifier|false|false||GRAMnull|Rh Negative Blood Group|Finding|false|false||NEGATIVE
null|Negative|Finding|false|false||NEGATIVE
null|Negative Finding|Finding|false|false||NEGATIVEnull|Expression Negative|Lab|false|false||NEGATIVEnull|Negative - qualifier|Modifier|false|false||NEGATIVE
null|Negative Charge|Modifier|false|false||NEGATIVEnull|Negative Number|LabModifier|false|false||NEGATIVEnull|Renal Osteodystrophy|Disorder|true|false||RODnull|KNTC1 gene|Finding|true|false||RODnull|Rod Photoreceptors|Anatomy|false|false||RODnull|Rod Device|Device|true|false||RODnull|Form-bacillus|Entity|true|false||RODnull|Rod Shape|Modifier|false|false||RODnull|Abscess|Disorder|false|false||ABSCESSnull|null|Finding|false|false||ABSCESSnull|Pelvis|Anatomy|false|false||PELVICnull|Respiratory Aspiration|Disorder|false|false||ASPIRATIONnull|Aspiration into respiratory tract|Finding|false|false||ASPIRATION
null|Endotracheal aspiration|Finding|false|false||ASPIRATION
null|Pulmonary aspiration|Finding|false|false||ASPIRATIONnull|null|Procedure|false|false||ASPIRATIONnull|Final report|Finding|false|false||FINAL REPORTnull|Diagnosis Type - Final|Finding|false|false||FINALnull|Final|Time|false|false||FINALnull|End-stage|Modifier|false|false||FINALnull|Report (document)|Finding|false|false||REPORTnull|Reporting|Procedure|false|false||REPORTnull|null|Attribute|false|false||REPORTnull|Gram's stain|Drug|false|false||GRAM STAIN
null|Gram's stain|Drug|false|false||GRAM STAINnull|Bacterial stain, routine|Procedure|false|false||GRAM STAINnull|gram|LabModifier|false|false||GRAMnull|Stains|Drug|false|false||STAINnull|Staining method|Procedure|false|false||STAINnull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Knowledge Field|Finding|false|false||FIELD
null|Force Field|Finding|false|false||FIELD
null|Field|Finding|false|false||FIELDnull|field - patient encounter|Procedure|false|false||FIELDnull|Specimen Type - Leukocytes|Finding|false|false||LEUKOCYTES
null|null|Finding|false|false||LEUKOCYTESnull|Leukocytes|Anatomy|false|false||LEUKOCYTESnull|Knowledge Field|Finding|true|false||FIELD
null|Force Field|Finding|true|false||FIELD
null|Field|Finding|true|false||FIELDnull|field - patient encounter|Procedure|true|false||FIELDnull|Gram-negative bacillus|Entity|false|false||GRAM NEGATIVE RODnull|gram|LabModifier|false|false||GRAMnull|Rh Negative Blood Group|Finding|false|false||NEGATIVE
null|Negative|Finding|false|false||NEGATIVE
null|Negative Finding|Finding|false|false||NEGATIVEnull|Expression Negative|Lab|false|false||NEGATIVEnull|Negative - qualifier|Modifier|false|false||NEGATIVE
null|Negative Charge|Modifier|false|false||NEGATIVEnull|Negative Number|LabModifier|false|false||NEGATIVEnull|Renal Osteodystrophy|Disorder|true|false||RODnull|KNTC1 gene|Finding|true|false||RODnull|Rod Photoreceptors|Anatomy|false|false||RODnull|Rod Device|Device|true|false||RODnull|Form-bacillus|Entity|true|false||RODnull|Rod Shape|Modifier|false|false||RODnull|Wound Culture|Procedure|false|false||WOUND CULTUREnull|Traumatic Wound|Disorder|false|false||WOUND
null|Wounds and Injuries|Disorder|false|false||WOUND
null|Traumatic injury|Disorder|false|false||WOUNDnull|Route of Administration - Wound|Finding|false|false||WOUND
null|null|Finding|false|false||WOUND
null|Specimen Type - Wound|Finding|false|false||WOUNDnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Growth & development aspects|Finding|true|false||GROWTH
null|Tissue Growth|Finding|true|false||GROWTH
null|Growth|Finding|true|false||GROWTH
null|growth aspects|Finding|true|false||GROWTHnull|Growth action|Phenomenon|true|false||GROWTHnull|Anaerobic microbial culture|Procedure|false|false||ANAEROBIC CULTUREnull|Anaerobic|Modifier|false|false||ANAEROBICnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Bacteroides fragilis group|Entity|false|false||BACTEROIDES FRAGILIS GROUPnull|Bacteroides fragilis infection in conditions classified elsewhere and of unspecified site|Disorder|false|false||BACTEROIDES FRAGILISnull|Bacteroides fragilis|Entity|false|false||BACTEROIDES FRAGILISnull|Bacteroides|Entity|false|false||BACTEROIDESnull|Group Specimen|Finding|false|false||GROUP
null|Stage Grouping|Finding|false|false||GROUP
null|Group Object|Finding|false|false||GROUP
null|Groups|Finding|false|false||GROUPnull|Population Group|Subject|false|false||GROUP
null|Social group|Subject|false|false||GROUP
null|User Group|Subject|false|false||GROUPnull|Growth & development aspects|Finding|false|false||GROWTH
null|Tissue Growth|Finding|false|false||GROWTH
null|Growth|Finding|false|false||GROWTH
null|growth aspects|Finding|false|false||GROWTHnull|Growth action|Phenomenon|false|false||GROWTHnull|beta-Lactamase|Drug|false|false||BETA LACTAMASE
null|beta-Lactamase|Drug|false|false||BETA LACTAMASEnull|Greek letter beta|Finding|false|false||BETAnull|Beta <eudicots>|Entity|false|false||BETAnull|Beta Distribution|LabModifier|false|false||BETAnull|lactamase|Drug|false|false||LACTAMASE
null|lactamase|Drug|false|false||LACTAMASEnull|BRAF Gene Rearrangement|Disorder|false|false||POSITIVEnull|Rh Positive Blood Group|Finding|false|false||POSITIVE
null|Positive Finding|Finding|false|false||POSITIVE
null|Positive|Finding|false|false||POSITIVEnull|Positive Charge|Modifier|false|false||POSITIVEnull|Positive Number|LabModifier|false|false||POSITIVEnull|Consistency of stool|Finding|false|false||STOOL     CONSISTENCYnull|Feces|Finding|false|false||STOOLnull|Stool seat|Device|false|false||STOOLnull|Consistency|Modifier|false|false||CONSISTENCYnull|Kind of quantity - Consistency|LabModifier|false|false||CONSISTENCYnull|Applicable|Modifier|true|false||APPLICABLE
null|null|Modifier|true|false||APPLICABLEnull|Source (property) (qualifier value)|Finding|true|false||Source
null|Term Source|Finding|true|false||Source
null|Source|Finding|true|false||Sourcenull|Feces|Finding|false|false||Stoolnull|Stool seat|Device|false|false||Stoolnull|Final report|Finding|false|false||FINAL REPORTnull|Diagnosis Type - Final|Finding|false|false||FINALnull|Final|Time|false|false||FINALnull|End-stage|Modifier|false|false||FINALnull|Report (document)|Finding|false|false||REPORTnull|Reporting|Procedure|false|false||REPORTnull|null|Attribute|false|false||REPORTnull|dna amplification|Finding|false|false||DNA amplificationnull|DNA|Drug|false|false||DNA
null|DNA|Drug|false|false||DNAnull|Gene Amplification Abnormality|Disorder|false|false||amplificationnull|Gene Amplification Technique|Procedure|false|false||amplificationnull|Amplification|Phenomenon|false|false||amplificationnull|Biological Assay|Procedure|false|false||assay
null|Assay|Procedure|false|false||assaynull|assay qualifier|Modifier|false|false||assaynull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Negative|Finding|false|false||Negative fornull|Rh Negative Blood Group|Finding|false|false||Negative
null|Negative|Finding|false|false||Negative
null|Negative Finding|Finding|false|false||Negativenull|Expression Negative|Lab|false|false||Negativenull|Negative - qualifier|Modifier|false|false||Negative
null|Negative Charge|Modifier|false|false||Negativenull|Negative Number|LabModifier|false|false||Negativenull|Toxigenic|Finding|true|false||toxigenicnull|DNA|Drug|false|false||DNA
null|DNA|Drug|false|false||DNAnull|Gene Amplification Abnormality|Disorder|false|false||amplificationnull|Gene Amplification Technique|Procedure|false|false||amplificationnull|Amplification|Phenomenon|false|false||amplificationnull|Biological Assay|Procedure|false|false||assay
null|Assay|Procedure|false|false||assaynull|assay qualifier|Modifier|false|false||assaynull|Reference range (qualifier value)|Modifier|false|false||Reference Rangenull|null|LabModifier|false|false||Reference Rangenull|Reference - MdfHmdMetSourceType|Finding|false|false||Reference
null|Reference Object|Finding|false|false||Reference
null|Reference source|Finding|false|false||Reference
null|Bibliographic Reference|Finding|false|false||Reference
null|Reference - HL7UpdateMode|Finding|false|false||Referencenull|Concept model range (foundation metadata concept)|Finding|false|false||Rangenull|Sample Range|LabModifier|false|false||Range
null|Range|LabModifier|false|false||Rangenull|Rh Negative Blood Group|Finding|false|false||Negative
null|Negative|Finding|false|false||Negative
null|Negative Finding|Finding|false|false||Negativenull|Expression Negative|Lab|false|false||Negativenull|Negative - qualifier|Modifier|false|false||Negative
null|Negative Charge|Modifier|false|false||Negativenull|Negative Number|LabModifier|false|false||Negativenull|BRIEF Health Literacy Screening Tool|Finding|false|false||Brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||Briefnull|Brief|Time|false|false||Briefnull|Shortened|Modifier|false|false||Briefnull|Hospital course|Finding|false|false||Hospital Coursenull|null|Attribute|false|false||Hospital Coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||Coursenull|ActInformationPrivacyReason - service|Finding|false|false||servicenull|Software Service|Device|false|false||servicenull|Services|Event|false|false||servicenull|Disease Management|Procedure|false|false||managementnull|Management Occupations|Subject|false|false||managementnull|Management procedure|Event|false|false||management
null|Administration occupational activities|Event|false|false||managementnull|Ileus|Disorder|false|false||ileus
null|Intestinal obstruction co-occurrent and due to decreased peristalsis|Disorder|false|false||ileusnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Nasogastric tube procedures|Procedure|false|false||nasogastric tubenull|Nasogastric tube|Device|false|false||nasogastric tubenull|Nasogastric Route of Administration|Finding|false|false||nasogastricnull|Nasogastric|Anatomy|false|false||nasogastricnull|Unspecified tube|Finding|false|false||tube
null|TUBE1 gene|Finding|false|false||tubenull|biomedical tube device|Device|false|false||tube
null|Packaging Tube|Device|false|false||tubenull|tube|Modifier|false|false||tubenull|Tube (unit of presentation)|LabModifier|false|false||tube
null|Tube Dosing Unit|LabModifier|false|false||tubenull|Decompression - action (qualifier value)|Finding|false|false||decompressionnull|Decompression|Procedure|false|false||decompression
null|Decompressive incision|Procedure|false|false||decompressionnull|external decompression|Phenomenon|false|false||decompressionnull|Peripherally Inserted Central Catheter Line Insertion|Procedure|false|false||PICCnull|Peripherally inserted central catheter (physical object)|Device|false|false||PICCnull|TAPBP protein, human|Drug|false|false||TPN
null|NADP|Drug|false|false||TPN
null|NADP|Drug|false|false||TPN
null|TAPBP protein, human|Drug|false|false||TPNnull|TAPBP wt Allele|Finding|false|false||TPN
null|TAPBP gene|Finding|false|false||TPNnull|Parenteral Nutrition, Total|Procedure|false|false||TPNnull|Blood culture|Procedure|true|false||Blood culturesnull|Blood and lymphatic system disorders|Disorder|false|false||Bloodnull|peripheral blood|Finding|false|false||Blood
null|Blood|Finding|false|false||Blood
null|In Blood|Finding|false|false||Bloodnull|Culture (Anthropological)|Finding|false|false||culturesnull|Gram-negative bacillus|Entity|false|false||gram negative rodsnull|gram|LabModifier|false|false||gramnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Rod Photoreceptors|Anatomy|false|false||rodsnull|ceftriaxone|Drug|true|false||ceftriaxone
null|ceftriaxone|Drug|true|false||ceftriaxonenull|Small amount|LabModifier|false|false||small amountnull|Small|LabModifier|false|false||smallnull|Amount class - Amount|Finding|false|false||amountnull|Quantity|LabModifier|false|false||amountnull|Flatulence|Finding|false|false||flatusnull|X-Ray Computed Tomography|Procedure|false|false||CT scannull|Radionuclide Imaging|Procedure|false|false||scan
null|Scanning|Procedure|false|false||scannull|Ileus|Disorder|false|false||ileus
null|Intestinal obstruction co-occurrent and due to decreased peristalsis|Disorder|false|false||ileusnull|Concern|Finding|false|false||concernnull|Possible|Finding|false|false||possiblenull|Possible diagnosis|Modifier|false|false||possible
null|Possibly Related to Intervention|Modifier|false|false||possiblenull|Urinary Incontinence|Finding|false|false||urine leaknull|Portion of urine|Finding|false|false||urine
null|null|Finding|false|false||urine
null|Urine|Finding|false|false||urine
null|In Urine|Finding|false|false||urine
null|Urine specimen|Finding|false|false||urinenull|Leaking|Finding|false|false||leaknull|effusion|Finding|false|false||free fluidnull|Free of (attribute)|Finding|false|false||freenull|Empty (qualifier)|Modifier|false|false||freenull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Structure of left lower quadrant of abdomen|Anatomy|false|false||LLQnull|Left lower quadrant|Modifier|false|false||LLQnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Interventional Radiology Procedure|Procedure|false|false||interventional radiologynull|Interventional radiology|Title|false|false||interventional radiologynull|interventional (invasive) radiology|Procedure|false|false||interventional
null|Interventional procedure|Procedure|false|false||interventionalnull|radiology referral type|Finding|false|false||radiology
null|Radiology Section ID|Finding|false|false||radiology
null|Encounter due to radiological examination|Finding|false|false||radiologynull|Radiology studies|Procedure|false|false||radiology
null|Diagnostic radiologic examination|Procedure|false|false||radiology
null|Radiographic imaging procedure|Procedure|false|false||radiologynull|Radiology Specialty|Title|false|false||radiologynull|Clamping Activity|Finding|false|false||clamp
null|PDZK1 wt Allele|Finding|false|false||clamp
null|PDZK1 gene|Finding|false|false||clamp
null|SPEF1 gene|Finding|false|false||clampnull|null|Device|false|false||clampnull|Clinical Trials|Procedure|false|false||trialnull|Pass (indicator)|Finding|false|false||passnull|Flatulence|Finding|false|false||flatusnull|Defecation|Finding|false|false||bowel movementsnull|Intestines|Anatomy|false|false||bowelnull|Movement|Finding|false|false||movementsnull|Clear liquid diet|Procedure|false|false||clear liquid dietnull|Clear liquid|Finding|false|false||clear liquidnull|Remote control command - Clear|Finding|false|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Liquid diet|Procedure|false|false||liquid dietnull|Liquid Dosage Form|Drug|false|false||liquid
null|Liquid substance|Drug|false|false||liquidnull|Liquid (finding)|Finding|false|false||liquidnull|Liquid diet|Procedure|false|false||liquidnull|Liquid (state of matter)|Modifier|false|false||liquidnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Repeat Object|Finding|false|false||Repeat
null|Repeat|Finding|false|false||Repeatnull|Repeat Pattern|Time|false|false||Repeatnull|Blood culture|Procedure|false|false||blood culturesnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Culture (Anthropological)|Finding|false|false||culturesnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Organism isolated in blood by culture|Lab|false|false||positive blood culturenull|BRAF Gene Rearrangement|Disorder|false|false||positivenull|Rh Positive Blood Group|Finding|false|false||positive
null|Positive Finding|Finding|false|false||positive
null|Positive|Finding|false|false||positivenull|Positive Charge|Modifier|false|false||positivenull|Positive Number|LabModifier|false|false||positivenull|Blood culture|Procedure|false|false||blood culturenull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Culture Dose Form|Drug|false|false||culturenull|Culture (Anthropological)|Finding|false|false||culture
null|Cultural aspects|Finding|false|false||culturenull|Microbial culture (procedure)|Procedure|false|false||culture
null|Laboratory culture|Procedure|false|false||culturenull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Citrobacter|Entity|false|false||citrobacternull|Diet (animal life circumstance)|Drug|false|false||Diet
null|Diet|Drug|false|false||Dietnull|diet - supply|Finding|false|false||Dietnull|Diet therapy|Procedure|false|false||Dietnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Diagnostic Service Section ID - Physical Therapy|Finding|false|false||physical therapynull|Physical therapy|Procedure|false|false||physical therapynull|Physical therapy (field)|Title|false|false||physical therapynull|physical examination (physical finding)|Finding|false|false||physical
null|Physical|Finding|false|false||physicalnull|Physical Examination|Procedure|false|false||physicalnull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|Rehabilitative Services|Finding|false|false||rehabilitative servicesnull|Rehabilitation therapy|Procedure|false|false||rehabilitativenull|Clinical Service|Procedure|false|false||servicesnull|Services|Event|false|false||servicesnull|Walkers|Device|false|false||walkernull|Helping Behavior|Finding|false|false||assistancenull|Assisted (qualifier value)|Modifier|false|false||assistancenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|ADMIN.FACILITY|Finding|false|false||facilitynull|Facility (object)|Device|false|false||facilitynull|TAPBP protein, human|Drug|false|false||TPN
null|NADP|Drug|false|false||TPN
null|NADP|Drug|false|false||TPN
null|TAPBP protein, human|Drug|false|false||TPNnull|TAPBP wt Allele|Finding|false|false||TPN
null|TAPBP gene|Finding|false|false||TPNnull|Parenteral Nutrition, Total|Procedure|false|false||TPNnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|null|Finding|false|false||regular dietnull|Regular|Modifier|false|false||regularnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Flatulence|Finding|false|false||passing flatusnull|null|Attribute|false|false||passing flatusnull|Flatulence|Finding|false|false||flatusnull|Defecation|Finding|false|false||bowel movementsnull|Intestines|Anatomy|false|false||bowelnull|Movement|Finding|false|false||movementsnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Accurate (qualifier value)|Modifier|false|false||accuratenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|levothyroxine sodium|Drug|false|false||Levothyroxine Sodium
null|levothyroxine sodium|Drug|false|false||Levothyroxine Sodium
null|levothyroxine sodium|Drug|false|false||Levothyroxine Sodiumnull|Synthetic Levothyroxine|Drug|false|false||Levothyroxine
null|Synthetic Levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxinenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|microgram|LabModifier|false|false||mcgnull|Daily|Time|false|false||DAILYnull|losartan potassium|Drug|false|false||Losartan Potassium
null|losartan potassium|Drug|false|false||Losartan Potassiumnull|losartan|Drug|false|false||Losartan
null|losartan|Drug|false|false||Losartannull|Potassium Drug Class|Drug|false|false||Potassium
null|Dietary Potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassiumnull|Potassium metabolic function|Finding|false|false||Potassiumnull|Potassium measurement|Procedure|false|false||Potassiumnull|Daily|Time|false|false||DAILYnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every six hours|Time|false|false||Q6Hnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|enoxaparin sodium|Drug|false|false||Enoxaparin Sodium
null|enoxaparin sodium|Drug|false|false||Enoxaparin Sodiumnull|enoxaparin|Drug|false|false||Enoxaparin
null|enoxaparin|Drug|false|false||Enoxaparinnull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|Daily|Time|false|false||DAILYnull|nitrofurantoin|Drug|false|false||Nitrofurantoin
null|nitrofurantoin|Drug|false|false||Nitrofurantoinnull|Macrobid|Drug|false|false||MacroBID
null|Macrobid|Drug|false|false||MacroBIDnull|Daily|Time|false|false||DAILYnull|oxycodone|Drug|false|false||OxyCODONE
null|oxycodone|Drug|false|false||OxyCODONEnull|Oxycodone measurement|Procedure|false|false||OxyCODONEnull|Immediate Release Dosage Form|Drug|false|false||Immediate Releasenull|Query Priority - Immediate|Finding|false|false||Immediate
null|immediate - ResponseCode|Finding|false|false||Immediatenull|Immediate|Time|false|false||Immediate
null|Stat (do immediately)|Time|false|false||Immediatenull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Every four hours|Time|false|false||Q4Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Moderate - Severity of Illness Code|Finding|false|false||Moderate
null|Moderate|Finding|false|false||Moderatenull|Moderate (severity modifier)|Modifier|false|false||Moderate
null|Moderate - Allergy Severity|Modifier|false|false||Moderate
null|Moderation|Modifier|false|false||Moderatenull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|ciprofloxacin hydrochloride|Drug|false|false||Ciprofloxacin HCl
null|ciprofloxacin hydrochloride|Drug|false|false||Ciprofloxacin HClnull|ciprofloxacin|Drug|false|false||Ciprofloxacin
null|ciprofloxacin|Drug|false|false||Ciprofloxacinnull|Flinders medical centre-7 marker|Drug|false|false||HCl
null|hydrochloride|Drug|false|false||HCl
null|hydrochloride|Drug|false|false||HClnull|Hairy Cell Leukemia|Disorder|false|false||HClnull|Every twelve hours|Time|false|false||Q12Hnull|Duration brand of oxymetazoline|Drug|false|false||Durationnull|Duration (temporal concept)|Time|false|false||Durationnull|7 days|Time|false|false||7 Daysnull|day|Time|false|false||Daysnull|Last|Modifier|false|false||Lastnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|metronidazole|Drug|false|false||MetroNIDAZOLE
null|metronidazole|Drug|false|false||MetroNIDAZOLEnull|Every six hours|Time|false|false||Q6Hnull|Duration brand of oxymetazoline|Drug|false|false||Durationnull|Duration (temporal concept)|Time|false|false||Durationnull|7 days|Time|false|false||7 Daysnull|day|Time|false|false||Daysnull|Last|Modifier|false|false||Lastnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|sennosides, USP|Drug|false|false||Senna
null|sennosides, USP|Drug|false|false||Sennanull|Senna alexandrina|Entity|false|false||Senna
null|Senna Plant|Entity|false|false||Sennanull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every six hours|Time|false|false||Q6Hnull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|enoxaparin sodium|Drug|false|false||Enoxaparin Sodium
null|enoxaparin sodium|Drug|false|false||Enoxaparin Sodiumnull|enoxaparin|Drug|false|false||Enoxaparin
null|enoxaparin|Drug|false|false||Enoxaparinnull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|Daily|Time|false|false||DAILYnull|Firstly|Modifier|false|false||Firstnull|First (number)|LabModifier|false|false||Firstnull|Unit dose|LabModifier|false|false||Dose
null|Dosage|LabModifier|false|false||Dosenull|next - HtmlLinkType|Finding|false|false||Nextnull|Following|Time|false|false||Next
null|Then|Time|false|false||Nextnull|Adjacent|Modifier|false|false||Nextnull|Extended Priority Codes - Routine|Finding|false|false||Routine
null|Report priority - Routine|Finding|false|false||Routine
null|Admission Type - Routine|Finding|false|false||Routine
null|Level of Care - Routine|Finding|false|false||Routine
null|Processing priority - Routine|Finding|false|false||Routine
null|Referral priority - Routine|Finding|false|false||Routinenull|Routine coag|Procedure|false|false||Routinenull|Priority - Routine|Time|false|false||Routinenull|Routine|Modifier|false|false||Routinenull|Administration (procedure)|Procedure|false|false||Administrationnull|Administration occupational activities|Event|false|false||Administrationnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||Time
null|Time (foundation metadata concept)|Finding|false|false||Time
null|Value type - Time|Finding|false|false||Time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||Time
null|Data types - Time|Finding|false|false||Time
null|null|Finding|false|false||Timenull|Time|Time|false|false||Timenull|levothyroxine sodium|Drug|false|false||Levothyroxine Sodium
null|levothyroxine sodium|Drug|false|false||Levothyroxine Sodium
null|levothyroxine sodium|Drug|false|false||Levothyroxine Sodiumnull|Synthetic Levothyroxine|Drug|false|false||Levothyroxine
null|Synthetic Levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxinenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|microgram|LabModifier|false|false||mcgnull|Daily|Time|false|false||DAILYnull|lorazepam|Drug|false|false||LORazepam
null|lorazepam|Drug|false|false||LORazepamnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Anxiety Disorders|Disorder|false|false||anxiety
null|Anxiety|Disorder|false|false||anxietynull|Anxiety symptoms|Finding|false|false||anxietynull|losartan potassium|Drug|false|false||Losartan Potassium
null|losartan potassium|Drug|false|false||Losartan Potassiumnull|losartan|Drug|false|false||Losartan
null|losartan|Drug|false|false||Losartannull|Potassium Drug Class|Drug|false|false||Potassium
null|Dietary Potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassiumnull|Potassium metabolic function|Finding|false|false||Potassiumnull|Potassium measurement|Procedure|false|false||Potassiumnull|Daily|Time|false|false||DAILYnull|nitrofurantoin|Drug|false|false||Nitrofurantoin
null|nitrofurantoin|Drug|false|false||Nitrofurantoinnull|Macrobid|Drug|false|false||MacroBID
null|Macrobid|Drug|false|false||MacroBIDnull|Daily|Time|false|false||DAILYnull|oxycodone|Drug|false|false||OxyCODONE
null|oxycodone|Drug|false|false||OxyCODONEnull|Oxycodone measurement|Procedure|false|false||OxyCODONEnull|Immediate Release Dosage Form|Drug|false|false||Immediate Releasenull|Query Priority - Immediate|Finding|false|false||Immediate
null|immediate - ResponseCode|Finding|false|false||Immediatenull|Immediate|Time|false|false||Immediate
null|Stat (do immediately)|Time|false|false||Immediatenull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Every four hours|Time|false|false||Q4Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Moderate - Severity of Illness Code|Finding|false|false||Moderate
null|Moderate|Finding|false|false||Moderatenull|Moderate (severity modifier)|Modifier|false|false||Moderate
null|Moderate - Allergy Severity|Modifier|false|false||Moderate
null|Moderation|Modifier|false|false||Moderatenull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|long-term care|Procedure|false|false||Extended Carenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Malignant neoplasm of urinary bladder|Disorder|false|false||bladder cancer
null|Carcinoma of bladder|Disorder|false|false||bladder cancer
null|Bladder Neoplasm|Disorder|false|false||bladder cancernull|Neoplasm of uncertain or unknown behavior of bladder|Disorder|false|false||bladder
null|Benign neoplasm of bladder|Disorder|false|false||bladder
null|Carcinoma in situ of bladder|Disorder|false|false||bladdernull|Procedures on bladder|Procedure|false|false||bladdernull|Urinary Bladder|Anatomy|false|false||bladdernull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Postoperative Period|Time|false|false||post-operativenull|Ileus|Disorder|false|false||ileus
null|Intestinal obstruction co-occurrent and due to decreased peristalsis|Disorder|false|false||ileusnull|Bacteremia|Finding|false|false||bacteremianull|Citrobacter|Entity|false|false||CITROBACTERnull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Pelvic abscess|Disorder|false|false||pelvic abscessnull|Pelvis|Anatomy|false|false||pelvicnull|Abscess|Disorder|false|false||abscessnull|null|Finding|false|false||abscessnull|Bacteroides fragilis infection in conditions classified elsewhere and of unspecified site|Disorder|false|false||BACTEROIDES FRAGILISnull|Bacteroides fragilis|Entity|false|false||BACTEROIDES FRAGILISnull|Bacteroides|Entity|false|false||BACTEROIDESnull|Group Specimen|Finding|false|false||GROUP
null|Stage Grouping|Finding|false|false||GROUP
null|Group Object|Finding|false|false||GROUP
null|Groups|Finding|false|false||GROUPnull|Population Group|Subject|false|false||GROUP
null|Social group|Subject|false|false||GROUP
null|User Group|Subject|false|false||GROUPnull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Disease|Disorder|false|false||Conditionnull|Logical Condition|Finding|false|false||Conditionnull|null|Attribute|false|false||Conditionnull|Condition|Modifier|false|false||Conditionnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Helping Behavior|Finding|false|false||assistancenull|Assisted (qualifier value)|Modifier|false|false||assistancenull|AICDA protein, human|Drug|false|false||aid
null|AICDA protein, human|Drug|false|false||aidnull|AICDA wt Allele|Finding|false|false||aid
null|AICDA gene|Finding|false|false||aidnull|AID - Artificial insemination by donor|Procedure|false|false||aid
null|dacarbazine/doxorubicin/ifosfamide protocol|Procedure|false|false||aidnull|Aid (attribute)|Modifier|false|false||aid
null|Assisted (qualifier value)|Modifier|false|false||aidnull|Walkers|Device|false|false||walkernull|CANE, INCLUDES CANES OF ALL MATERIALS, ADJUSTABLE OR FIXED, WITH TIP|Device|false|false||canenull|Cane - plant part|Entity|false|false||canenull|Discharge instructions|Finding|false|false||Discharge Instructionsnull|hospital discharge instructions (treatment)|Procedure|false|false||Discharge Instructionsnull|null|Attribute|false|false||Discharge Instructionsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|Instructions provided|Finding|false|false||instructions providednull|null|Attribute|false|false||instructions providednull|Instructions|Finding|false|false||instructions
null|Instruction [Publication Type]|Finding|false|false||instructionsnull|null|Attribute|false|false||instructionsnull|Ostomy|Procedure|false|false||Ostomynull|Nurse Specialists|Subject|false|false||nurse specialistnull|Nurses|Subject|false|false||nursenull|United States Military enlisted E4 (qualifier value)|Finding|false|false||specialistnull|Specialist Physician|Subject|false|false||specialist
null|Hospital specialist|Subject|false|false||specialist
null|Specialist|Subject|false|false||specialistnull|Details|Modifier|false|false||detailsnull|required - HL7ConformanceInclusion|Finding|false|false||required
null|Required - Escort Required|Finding|false|false||required
null|required - HL7V3Conformance|Finding|false|false||required
null|Requirement|Finding|false|false||required
null|required - ParticipationSignature|Finding|false|false||required
null|required - CodingRationale|Finding|false|false||requirednull|Continuity Assessment Record and Evaluation|Finding|false|false||care
null|In care (finding)|Finding|false|false||carenull|care activity|Event|false|false||carenull|Disease Management|Procedure|false|false||managementnull|Management Occupations|Subject|false|false||managementnull|Management procedure|Event|false|false||management
null|Administration occupational activities|Event|false|false||managementnull|Urostomy procedure|Procedure|false|false||Urostomynull|Urological stoma|Anatomy|false|false||Urostomynull|Resume - Remote control command|Finding|false|false||Resume
null|Curriculum Vitae|Finding|false|false||Resume
null|resume - DataOperation|Finding|false|false||Resumenull|Pre-admission Encounter|Finding|false|false||pre-admissionnull|Pre-admission|Time|false|false||pre-admissionnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Always - AcknowledgementCondition|Finding|false|false||Always
null|All of the Time|Finding|false|false||Alwaysnull|Always (frequency)|Time|false|false||Alwaysnull|Call - dosing instruction fragment|Finding|true|false||call
null|Call (Instruction)|Finding|true|false||call
null|Decision|Finding|true|false||call
null|CHL1 gene|Finding|true|false||callnull|Reporting|Procedure|true|false||informnull|inform|Event|true|false||informnull|Review (Publication Type)|Finding|true|false||review
null|Act Class - review|Finding|true|false||reviewnull|Pharmaceutical Preparations|Drug|true|false||medicationnull|medication - HL7 publishing domain|Finding|true|false||medication
null|Medications|Finding|true|false||medicationnull|Changing|Finding|true|false||changesnull|Changed status|LabModifier|true|false||changesnull|Postoperative Period|Time|true|false||post-operativenull|Course|Time|true|false||coursenull|Primary care provider|Subject|false|false||primary care doctornull|Location Service Code - Primary Care|Finding|false|false||primary carenull|Primary Health Care|Procedure|false|false||primary carenull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|Continuity Assessment Record and Evaluation|Finding|false|false||care
null|In care (finding)|Finding|false|false||carenull|care activity|Event|false|false||carenull|Doctor - Title|Finding|false|false||doctornull|Physicians|Subject|false|false||doctornull|Acetaminophen [EPC]|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophennull|Acetaminophen measurement|Procedure|false|false||acetaminophennull|ibuprofen|Drug|false|false||Ibuprofen
null|ibuprofen|Drug|false|false||Ibuprofennull|Demonstrates adequate pain control|Finding|false|false||pain controlnull|Pain control|Procedure|false|false||pain control
null|Pain management (procedure)|Procedure|false|false||pain controlnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Control brand of phenylpropanolamine|Drug|false|false||control
null|CONTROL veterinary product|Drug|false|false||control
null|control substance|Drug|false|false||control
null|Control brand of phenylpropanolamine|Drug|false|false||controlnull|Control - Relationship modifier|Finding|false|false||control
null|Control function|Finding|false|false||control
null|Scientific Control|Finding|false|false||controlnull|Control Groups|Subject|false|false||controlnull|True Control Status|Modifier|false|false||control
null|control aspects|Modifier|false|false||controlnull|ciprofloxacin and metronidazole|Drug|false|false||Ciprofloxacin and Metronidazolenull|ciprofloxacin|Drug|false|false||Ciprofloxacin
null|ciprofloxacin|Drug|false|false||Ciprofloxacinnull|metronidazole|Drug|false|false||Metronidazole
null|metronidazole|Drug|false|false||Metronidazolenull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Antibiotics|Drug|false|false||ANTIBIOTICnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|7 days|Time|false|false||7 daysnull|day|Time|false|false||daysnull|Act Relationship Subset - maximum|LabModifier|false|false||MAXIMUM
null|Maximum|LabModifier|false|false||MAXIMUMnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Tylenol|Drug|false|false||Tylenol
null|Tylenol|Drug|false|false||Tylenolnull|Acetaminophen [EPC]|Drug|false|false||ACETAMINOPHEN
null|acetaminophen|Drug|false|false||ACETAMINOPHEN
null|acetaminophen|Drug|false|false||ACETAMINOPHENnull|Acetaminophen measurement|Procedure|false|false||ACETAMINOPHENnull|gram|LabModifier|false|false||gramsnull|Source|Finding|false|false||sourcesnull|per day|Time|false|false||PER DAYnull|Transaction counts and value totals - day|Finding|false|false||DAY
null|Precision - day|Finding|false|false||DAYnull|Land Dayak Languages|Entity|false|false||DAYnull|day|Time|false|false||DAY
null|Daily|Time|false|false||DAYnull|ibuprofen|Drug|false|false||Ibuprofen
null|ibuprofen|Drug|false|false||Ibuprofennull|Proprietary Name|Finding|false|false||Brand namesnull|Name|Finding|false|false||namesnull|Always - AcknowledgementCondition|Finding|false|false||always
null|All of the Time|Finding|false|false||alwaysnull|Always (frequency)|Time|false|false||alwaysnull|With Food|Modifier|false|false||with foodnull|Food allergenic extracts|Drug|false|false||food
null|Food|Drug|false|false||food
null|Food allergenic extracts|Drug|false|false||foodnull|Neoplasm of uncertain or unknown behavior of stomach|Disorder|false|false||stomach
null|Stomach Diseases|Disorder|false|false||stomach
null|Benign neoplasm of stomach|Disorder|false|false||stomach
null|Carcinoma in situ of stomach|Disorder|false|false||stomachnull|Stomach problem|Finding|false|false||stomachnull|Procedure on stomach|Procedure|false|false||stomachnull|Stomach structure|Anatomy|false|false||stomach
null|Abdomen>Stomach|Anatomy|false|false||stomach
null|Stomach|Anatomy|false|false||stomachnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|null|Finding|false|false||black stool
null|Melena|Finding|false|false||black stoolnull|Black - ethnic group (ethnic group)|Subject|false|false||black
null|Black race|Subject|false|false||black
null|African|Subject|false|false||blacknull|Black - Structured Product Labeling Color|Modifier|false|false||black
null|Black color|Modifier|false|false||blacknull|Feces|Finding|false|false||stoolnull|Stool seat|Device|false|false||stoolnull|ibuprofen|Drug|false|false||Ibuprofen
null|ibuprofen|Drug|false|false||Ibuprofennull|Contact with machinery|Disorder|true|false||machinerynull|Industrial machine|Device|true|false||machinerynull|Alcohols|Drug|false|false||alcohol
null|Alcohols|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcoholnull|Alcohol - Recreational Drug Use Code|Finding|false|false||alcoholnull|Narcotics|Drug|false|false||narcotic
null|Narcotics|Drug|false|false||narcoticnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|activities (history)|Finding|false|false||activitiesnull|Activities|Event|false|false||activitiesnull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Urologists|Subject|false|false||urologistnull|Passenger|Subject|false|false||passengernull|Colace|Drug|false|false||Colace
null|Colace|Drug|false|false||Colacenull|Operative Surgical Procedures|Procedure|false|false||surgical
null|Surgical service|Procedure|false|false||surgicalnull|Constipation|Finding|false|false||constipationnull|Constipation|Finding|false|false||constipationnull|Relate - vinyl resin|Drug|false|false||relatednull|Role Link Type - related|Finding|false|false||related
null|Related (finding)|Finding|false|false||relatednull|Definitely Related to Intervention|Modifier|false|false||related
null|Relationships|Modifier|false|false||relatednull|Narcotics|Drug|false|false||narcotic
null|Narcotics|Drug|false|false||narcoticnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Loose stool|Finding|false|false||loose stoolnull|Loose|Modifier|false|false||loosenull|Feces|Finding|false|false||stoolnull|Stool seat|Device|false|false||stoolnull|rectal discharge diarrhea (physical finding)|Finding|false|false||diarrhea
null|Diarrhea|Finding|false|false||diarrheanull|Colace|Drug|true|false||Colace
null|Colace|Drug|true|false||Colacenull|Feces|Finding|true|false||stoolnull|Stool seat|Device|true|false||stoolnull|Laxatives|Drug|true|false||laxativenull|Heavy (weight) (qualifier value)|Modifier|true|false||heavy
null|Heavy (amount)|Modifier|true|false||heavynull|Lifting|Event|true|false||liftingnull|4 Weeks|Time|true|false||4 weeksnull|week|Time|true|false||weeksnull|Greater Than|LabModifier|true|false||more thannull|More|LabModifier|true|false||morenull|10 pounds|Finding|true|false||10 poundsnull|Pounds|LabModifier|true|false||poundsnull|Sedentary lifestyle|Finding|true|false||sedentarynull|Sedentary|Modifier|true|false||sedentarynull|Walking (function)|Finding|false|false||Walknull|Frequently|Time|false|false||frequentlynull|TNFSF14 protein, human|Drug|false|false||Light
null|TNFSF14 protein, human|Drug|false|false||Lightnull|Light - subjective measurement|Finding|false|false||Light
null|TNFSF14 wt Allele|Finding|false|false||Light
null|TNFSF14 gene|Finding|false|false||Light
null|Light color|Finding|false|false||Lightnull|Phototherapy|Procedure|false|false||Lightnull|Light|Phenomenon|false|false||Lightnull|Light (qualifier)|Modifier|false|false||Lightnull|activity level doing household chores|Finding|false|false||household choresnull|Households|Subject|false|false||householdnull|Cooking (activity)|Finding|false|false||cookingnull|Laundry|Finding|false|false||laundrynull|null|Attribute|false|false||laundrynull|Washing Dishes question|Finding|false|false||washing dishesnull|Wash (cleansing action)|Event|false|false||washingnull|Straining (finding)|Finding|true|false||strainingnull|Pulling|Finding|true|false||pulling
null|Does pull|Finding|true|false||pullingnull|Musculoskeletal torsion (function)|Finding|true|false||twisting
null|Torsion (malposition)|Finding|true|false||twistingnull|Vacuum (physical force)|Phenomenon|true|false||vacuumnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions