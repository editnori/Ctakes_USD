CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|Known|Modifier|false|false||Knownnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Adverse reaction to drug|Finding|true|false||Adverse Drug Reactionsnull|Adverse reaction to drug|Finding|true|false||Drug Reactionsnull|Pharmaceutical Preparations|Drug|false|false||Drug
null|Pharmacologic Substance|Drug|false|false||Drugnull|Drug problem|Finding|false|false||Drugnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Dyspnea on exertion|Finding|false|false||dyspnea on exertionnull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|Exertion|Finding|false|false||exertionnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Hypertensive disease|Disorder|false|false||HTNnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|DES protein, human|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|DES protein, human|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DESnull|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|Disorder|false|false||DESnull|DES gene|Finding|false|false||DESnull|Ischemic|Finding|false|false||ischemicnull|Systolic dysfunction|Finding|false|false||systolic dysfunctionnull|Systole|Finding|false|false||systolicnull|DYSFUNCTION - SKIN DISORDERS|Disorder|false|false||dysfunctionnull|Dysfunction|Finding|false|false||dysfunction
null|physiopathological|Finding|false|false||dysfunction
null|Functional disorder|Finding|false|false||dysfunctionnull|torsemide|Drug|false|false||torsemide
null|torsemide|Drug|false|false||torsemidenull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|4 Days|Time|false|false||4 daysnull|day|Time|false|false||daysnull|Dyspnea on exertion|Finding|false|false||dyspnea on exertionnull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|Exertion|Finding|false|false||exertionnull|Swelling of lower limb|Finding|false|false||leg swellingnull|Leg|Anatomy|false|false||leg
null|Lower Extremity|Anatomy|false|false||legnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|Gain|LabModifier|false|false||gainnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Congestive heart failure|Disorder|false|false||Heart Failure
null|Heart failure|Disorder|false|false||Heart Failurenull|Malignant neoplasm of heart|Disorder|false|false||Heart
null|benign neoplasm of heart|Disorder|false|false||Heartnull|HEART PROBLEM|Finding|false|false||Heartnull|Chest>Heart|Anatomy|false|false||Heart
null|Heart|Anatomy|false|false||Heartnull|Failure (biologic function)|Finding|false|false||Failure
null|Failure|Finding|false|false||Failure
null|Personal failure|Finding|false|false||Failurenull|Clinic|Device|false|false||Clinic
null|Ambulatory Care Facilities|Device|false|false||Clinicnull|Clinic|Entity|false|false||Clinic
null|Ambulatory Care Facilities|Entity|false|false||Clinicnull|Patient location type - Clinic|Modifier|false|false||Clinic
null|Person location type - Clinic|Modifier|false|false||Clinicnull|Persistent|Time|false|false||persistentnull|Dyspnea on exertion|Finding|false|false||dyspnea on exertionnull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|Exertion|Finding|false|false||exertionnull|Paroxysmal nocturnal dyspnea|Disorder|false|false||PNDnull|NPPA wt Allele|Finding|false|false||PND
null|NPPA gene|Finding|false|false||PNDnull|null|Time|false|false||priornull|Hospitalization|Procedure|false|false||hospitalizationnull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|torsemide|Drug|false|false||torsemide
null|torsemide|Drug|false|false||torsemidenull|Initially|Time|false|false||initiallynull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Holidays|Event|false|false||holidaynull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Sodium Chloride, Dietary|Drug|false|false||salt
null|sodium chloride|Drug|false|false||salt
null|Salts|Drug|false|false||saltnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Slow|Modifier|false|false||slownull|Onset of (contextual qualifier)|Modifier|false|false||onsetnull|Age of Onset|LabModifier|false|false||onsetnull|Dyspnea on exertion|Finding|false|false||dyspnea on exertionnull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|Exertion|Finding|false|false||exertionnull|Pharmaceutical Preparations|Drug|true|false||medicationnull|medication - HL7 publishing domain|Finding|true|false||medication
null|Medications|Finding|true|false||medicationnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Palpitations|Finding|false|false||palpitationsnull|Palpitations|Finding|false|false||palpitationsnull|Paroxysmal nocturnal dyspnea|Disorder|false|false||PNDnull|NPPA wt Allele|Finding|false|false||PND
null|NPPA gene|Finding|false|false||PNDnull|null|Finding|false|false||exercise tolerancenull|null|Attribute|false|false||exercise tolerance
null|Exercise Tolerance|Attribute|false|false||exercise tolerancenull|Exercise|Finding|false|false||exercisenull|Exercise Pain Management|Procedure|false|false||exercisenull|Physiologic tolerance|Finding|false|false||tolerance
null|Mental tolerance|Finding|false|false||tolerance
null|Immune Tolerance|Finding|false|false||tolerance
null|Drug Tolerance|Finding|false|false||tolerancenull|Tolerance|Modifier|false|false||tolerancenull|Unable|Finding|false|false||unablenull|Foot|Anatomy|false|false||feetnull|Foot Unit of Length|LabModifier|false|false||feetnull|sleeping upright or using specific number of extra pillows (orthopnea)|Finding|false|false||orthopnea
null|Orthopnea|Finding|false|false||orthopneanull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Bilateral|Modifier|false|false||bilateralnull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Peripheral edema|Finding|false|false||extremity edemanull|Limb structure|Anatomy|false|false||extremitynull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Basilar Rales|Finding|false|false||crackles
null|Rales|Finding|false|false||cracklesnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Plain chest X-ray|Procedure|false|false||CXRnull|NPPB protein, human|Drug|false|false||BNP
null|NPPB protein, human|Drug|false|false||BNP
null|nesiritide|Drug|false|false||BNP
null|nesiritide|Drug|false|false||BNP
null|nesiritide|Drug|false|false||BNPnull|NPPB wt Allele|Finding|false|false||BNP
null|NPPB gene|Finding|false|false||BNPnull|Brain natriuretic peptide measurement|Procedure|false|false||BNPnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Lasix|Drug|false|false||Lasix
null|Lasix|Drug|false|false||Lasixnull|Initial (abbreviation)|Finding|false|false||initialnull|Initially|Time|false|false||initialnull|Firstly|Modifier|false|false||initialnull|null|Time|false|false||Prior tonull|null|Time|false|false||Priornull|Transfer - product ownership|Finding|false|false||transfer
null|Transfer Technique|Finding|false|false||transfer
null|ActClass - transfer|Finding|false|false||transfer
null|null|Finding|false|false||transfernull|Transfer (immobility management)|Procedure|false|false||transfernull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Laboratory test finding|Lab|false|false||labsnull|Sodium supplements|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|Sodium Drug Class|Drug|false|false||sodiumnull|Sodium metabolic function|Finding|false|false||sodiumnull|Sodium measurement|Procedure|false|false||sodiumnull|chloride ion|Drug|false|false||Chloride
null|Chlorides|Drug|false|false||Chloridenull|Chloride metabolic function|Finding|false|false||Chloridenull|Chloride measurement|Procedure|false|false||Chloridenull|sodium bicarbonate|Drug|false|false||Bicarb
null|sodium bicarbonate|Drug|false|false||Bicarbnull|Blood Urea Nitrogen|Drug|false|false||BUN
null|Blood Urea Nitrogen|Drug|false|false||BUNnull|Blood urea nitrogen measurement|Procedure|false|false||BUNnull|creatinine|Drug|false|false||Creatinine
null|creatinine|Drug|false|false||Creatininenull|Creatinine metabolic function|Finding|false|false||Creatininenull|Creatinine measurement|Procedure|false|false||Creatininenull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|NPPB protein, human|Drug|false|false||BNP
null|NPPB protein, human|Drug|false|false||BNP
null|nesiritide|Drug|false|false||BNP
null|nesiritide|Drug|false|false||BNP
null|nesiritide|Drug|false|false||BNPnull|NPPB wt Allele|Finding|false|false||BNP
null|NPPB gene|Finding|false|false||BNPnull|Brain natriuretic peptide measurement|Procedure|false|false||BNPnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Blood Platelets|Anatomy|false|false||Plateletnull|Leukocytes|Anatomy|false|false||WBCnull|Urinalysis; qualitative or semiquantitative, except immunoassays|Procedure|false|false||Urinalysis
null|Urinalysis|Procedure|false|false||Urinalysisnull|Still|Disorder|false|false||stillnull|Pending - Allergy Clinical Status|Finding|false|false||pending
null|Pending - referral status|Finding|false|false||pendingnull|Pending - status|Time|false|false||pendingnull|pending - ManagedParticipationStatus|Modifier|false|false||pending
null|pending - RoleStatus|Modifier|false|false||pending
null|Pending - Day type|Modifier|false|false||pendingnull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|Leukocyte adhesion deficiency type 1|Disorder|false|false||LAD
null|Leukocyte adhesion deficiency|Disorder|false|false||LADnull|ITGB2 wt Allele|Finding|false|false||LAD
null|DLD gene|Finding|false|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false||LADnull|Ladino Language|Entity|false|false||LADnull|Twi language|Entity|false|false||TWInull|inferiority|Finding|false|false||inferiornull|Inferior|Modifier|false|false||inferiornull|Lead Device|Device|false|false||leadsnull|null|Finding|false|false||unchangednull|About The Same|Modifier|false|false||unchangednull|null|Time|false|false||priornull|Floor (anatomic)|Anatomy|false|false||floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Hypertensive disease|Disorder|false|false||hypertensionnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||diabetes
null|Diabetes|Disorder|false|false||diabetes
null|Diabetes Mellitus|Disorder|false|false||diabetesnull|Cyclophosphamide/Doxorubicin/Vincristine|Drug|false|false||CVAnull|Acute ill-defined cerebrovascular disease|Disorder|false|false||CVA
null|Cerebrovascular accident|Disorder|false|false||CVAnull|Cerebellum|Anatomy|false|false||cerebellarnull|Medullary - body parts|Anatomy|false|false||medullary
null|Medulla Oblongata|Anatomy|false|false||medullary
null|Adrenal Medulla|Anatomy|false|false||medullarynull|Cerebrovascular accident|Disorder|false|false||strokenull|Stroke (heart beat)|Finding|false|false||strokenull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Burning Mouth Syndrome|Disorder|false|false||BMSnull|Circumflex|Modifier|false|false||circumflexnull|Peripheral Arterial Diseases|Disorder|false|false||peripheral arterial disease
null|Peripheral Vascular Diseases|Disorder|false|false||peripheral arterial diseasenull|Peripheral|Modifier|false|false||peripheralnull|Arteriopathic disease|Disorder|false|false||arterial diseasenull|Arteries|Anatomy|false|false||arterialnull|Arterial|Modifier|false|false||arterialnull|Disease|Disorder|false|false||diseasenull|Intermittent Claudication|Disorder|false|false||claudicationnull|Claudication (finding)|Finding|false|false||claudication
null|Lameness|Finding|false|false||claudicationnull|Blood Vessel|Anatomy|false|false||vascularnull|Vascular|Modifier|false|false||vascularnull|Stage level 4|Finding|false|false||stage IVnull|Tumor stage|Attribute|false|false||stagenull|Stage|Time|false|false||stage
null|Phase|Time|false|false||stagenull|Chronic Kidney Diseases|Disorder|false|false||CKDnull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Gastroesophageal reflux disease|Disorder|false|false||GERDnull|Terminal esophageal web|Disorder|false|false||esophageal ringsnull|Esophageal Diseases|Disorder|false|false||esophagealnull|Esophageal|Modifier|false|false||esophagealnull|Ring device|Device|false|false||ringsnull|ring form of protozoa|Entity|false|false||ringsnull|Indirect exposure mechanism - Father|Finding|false|false||Father
null|Relationship - Father|Finding|false|false||Father
null|Father - courtesy title|Finding|false|false||Fathernull|Father (person)|Subject|false|false||Fathernull|Lung diseases|Disorder|false|false||lung diseasenull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|Disease|Disorder|false|false||diseasenull|Relationship - Mother|Finding|false|false||Mothernull|Mother (person)|Subject|false|false||Mothernull|unknown vaccine or immune globulin|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|unknown vaccine or immune globulin|Drug|false|false||unknownnull|Unknown - Patient_s Relationship to Insured|Finding|false|false||unknown
null|Unknown - Special Program Code|Finding|false|false||unknown
null|Unknown - Production Class Code|Finding|false|false||unknown
null|Unknown - Patient Outcome|Finding|false|false||unknown
null|Unknown - Recreational Drug Use Code|Finding|false|false||unknown
null|Unknown - Escort Required|Finding|false|false||unknown
null|Unknown - Transport Arranged|Finding|false|false||unknown
null|Unknown - Living Arrangement|Finding|false|false||unknown
null|Unknown - Employment Status|Finding|false|false||unknown
null|Unknown - Relationship|Finding|false|false||unknown
null|Unknown - publishing section|Finding|false|false||unknown
null|Unknown Publicity Code|Finding|false|false||unknown
null|Unknown - Event reason|Finding|false|false||unknown
null|Unknown - Religion|Finding|false|false||unknown
null|Unknown - Organ Donor Code|Finding|false|false||unknown
null|unknown - NullFlavor|Finding|false|false||unknown
null|Unknown - Notify Clergy Code|Finding|false|false||unknown
null|Unknown - Administrative Gender|Finding|false|false||unknown
null|Unknown - Patient Condition Code|Finding|false|false||unknown
null|Unknown - Living Will Code|Finding|false|false||unknown
null|Marital Status - Unknown|Finding|false|false||unknown
null|Unknown - mode of arrival code|Finding|false|false||unknown
null|Unknown - Patient Class|Finding|false|false||unknown
null|Unknown - Event Expected|Finding|false|false||unknown
null|Unknown - Expanded yes/no indicator|Finding|false|false||unknown
null|Unknown - Immunization Registry Status|Finding|false|false||unknown
null|Unknown - Container status|Finding|false|false||unknown
null|Unknown - CWE statuses|Finding|false|false||unknown
null|Unknown - Job Status|Finding|false|false||unknown
null|Unknown - Precaution Code|Finding|false|false||unknown
null|Unknown - Contact Role|Finding|false|false||unknown
null|Unknown - Living Dependency|Finding|false|false||unknownnull|Ethnic group unknown|Subject|false|false||unknownnull|Unknown - Allergy Severity|Modifier|false|false||unknown
null|Unknown - HL7 update mode|Modifier|false|false||unknown
null|Unknown|Modifier|false|false||unknownnull|Science of Etiology|Finding|false|false||cause
null|Etiology aspects|Finding|false|false||causenull|Early|Time|false|false||earlynull|DFFB protein, human|Drug|true|false||CAD
null|DFFB protein, human|Drug|true|false||CADnull|Cold Hemagglutinin Disease|Disorder|true|false||CAD
null|Coronary heart disease|Disorder|true|false||CAD
null|Coronary Artery Disease|Disorder|true|false||CADnull|CAD gene|Finding|true|false||CAD
null|CALD1 wt Allele|Finding|true|false||CAD
null|B4GALNT2 gene|Finding|true|false||CAD
null|DFFB wt Allele|Finding|true|false||CAD
null|ACOD1 gene|Finding|true|false||CAD
null|DFFB gene|Finding|true|false||CADnull|cytarabine/daunorubicin protocol|Procedure|true|false||CAD
null|Computer Assisted Diagnosis|Procedure|true|false||CAD
null|Collision-Induced Dissociation|Procedure|true|false||CAD
null|CyADIC regimen|Procedure|true|false||CADnull|Caddo language|Entity|true|false||CADnull|Sudden (qualifier value)|Modifier|false|false||suddennull|Cardiac attachment|Finding|true|false||cardiacnull|Heart|Anatomy|false|false||cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||cardiacnull|Event Consequence - Death|Finding|false|false||death
null|Death (finding)|Finding|false|false||death
null|Cessation of life|Finding|false|false||deathnull|Known|Modifier|false|false||knownnull|History of malignant neoplasm|Finding|true|false||history of cancernull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Malignant Neoplasms|Disorder|true|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|true|false||cancernull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|physical examination (physical finding)|Finding|false|false||PHYSICAL EXAMINATIONnull|Physical Examination|Procedure|false|false||PHYSICAL EXAMINATIONnull|physical examination (physical finding)|Finding|false|false||PHYSICAL
null|Physical|Finding|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||EXAMINATION
null|Medical Examination|Procedure|false|false||EXAMINATIONnull|Examination|Event|false|false||EXAMINATIONnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GENERALnull|General medical service|Procedure|false|false||GENERALnull|Generalized|Modifier|false|false||GENERALnull|Obesity|Disorder|false|false||obesenull|Sitting upright|Finding|false|false||sitting uprightnull|Special Handling Code - Upright|Finding|false|false||uprightnull|Entity Handling - upright|Phenomenon|false|false||uprightnull|Upright|Modifier|false|false||uprightnull|BORNHOLM EYE DISEASE|Disorder|false|false||bednull|Bachelor of Education|Finding|false|false||bednull|Beds|Device|false|false||bednull|Patient Location - Bed|Modifier|false|false||bednull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|Mood (psychological function)|Finding|false|false||Mood
null|mood (physical finding)|Finding|false|false||Mood
null|Mood (attribute)|Finding|false|false||Moodnull|null|Attribute|false|false||Moodnull|Appropriate|Modifier|false|false||appropriatenull|HEENT|Anatomy|false|false||HEENTnull|Scleral Diseases|Disorder|false|false||Scleranull|examination of sclera|Procedure|false|false||Scleranull|Sclera|Anatomy|false|false||Scleranull|Anicteric|Finding|false|false||anictericnull|Pupil equal round and reacting to light|Finding|false|false||PERRLnull|Malignant neoplasm of conjunctiva|Disorder|false|false||Conjunctiva
null|Benign neoplasm of conjunctiva|Disorder|false|false||Conjunctiva
null|Conjunctival Diseases|Disorder|false|false||Conjunctivanull|Specimen Type - Conjunctiva|Finding|false|false||Conjunctiva
null|null|Finding|false|false||Conjunctivanull|examination of conjunctiva|Procedure|false|false||Conjunctiva
null|Procedure on conjunctiva|Procedure|false|false||Conjunctivanull|Structure of palpebral conjunctiva|Anatomy|false|false||Conjunctiva
null|conjunctiva|Anatomy|false|false||Conjunctivanull|Pink color|Modifier|false|false||pinknull|Pallor of skin|Finding|true|false||pallornull|Cyanosis|Finding|true|false||cyanosisnull|Oral mucous membrane structure|Anatomy|false|false||oral mucosanull|Oral Dosage Form|Drug|false|false||oralnull|Oral Route of Administration|Finding|false|false||oral
null|Oral (intended site)|Finding|false|false||oralnull|Oral cavity|Anatomy|false|false||oralnull|Oral|Modifier|false|false||oralnull|null|Finding|false|false||mucosanull|Mucous Membrane|Anatomy|false|false||mucosanull|Passive joint movement of neck (finding)|Finding|false|false||NECK
null|Neck problem|Finding|false|false||NECKnull|dendritic spine neck|Anatomy|false|false||NECK
null|Neck|Anatomy|false|false||NECKnull|Supple|Finding|false|false||Supplenull|Jugular venous pressure|Finding|false|false||JVPnull|Cardiac attachment|Finding|false|false||CARDIACnull|Heart|Anatomy|false|false||CARDIACnull|Cardiac - anatomy qualifier|Modifier|false|false||CARDIACnull|Point of Maximum Impulse|Finding|false|false||PMI
null|TMEM11 gene|Finding|false|false||PMI
null|PMM2 wt Allele|Finding|false|false||PMI
null|PMM2 gene|Finding|false|false||PMI
null|MPI gene|Finding|false|false||PMInull|Prostate Mechanical Imager|Device|false|false||PMInull|Space of intercostal compartment|Anatomy|false|false||intercostal space
null|Structure of intercostal space|Anatomy|false|false||intercostal spacenull|Intercostal|Modifier|false|false||intercostalnull|Space (Astronomy)|Phenomenon|false|false||spacenull|Space - property|Modifier|false|false||spacenull|Midclavicular|Modifier|false|false||midclavicularnull|Line Specimen|Drug|false|false||line
null|Long Interspersed Elements|Drug|false|false||line
null|Long Interspersed Elements|Drug|false|false||linenull|line source specimen code|Finding|false|false||linenull|Intravascular line|Device|false|false||linenull|Linear|Modifier|false|false||linenull|Line Unit of Length|LabModifier|false|false||linenull|Heart murmur|Finding|true|false||murmursnull|Pericardial friction rub|Finding|true|false||rubsnull|Cardiac thrill (finding)|Finding|false|false||thrillsnull|hoist [device]|Device|false|false||liftsnull|Lung|Anatomy|false|false||LUNGSnull|Respiratory, thoracic and mediastinal disorders|Disorder|false|false||Respnull|Respiratory rate|Attribute|false|false||Respnull|Unlabored|Finding|false|false||unlaborednull|Use of accessory muscles|Finding|true|false||accessory muscle usenull|Accessory skeletal muscle|Disorder|true|false||accessory musclenull|Accessory|Device|true|false||accessorynull|Muscle (organ)|Anatomy|false|false||muscle
null|Muscle Tissue|Anatomy|false|false||musclenull|Use - dosing instruction imperative|Finding|true|false||use
null|utilization qualifier|Finding|true|false||use
null|Usage|Finding|true|false||usenull|dyspneic|Finding|false|false||dyspneicnull|Endoglin, human|Drug|false|false||end
null|Endoglin, human|Drug|false|false||endnull|end - ActRelationshipCheckpoint|Finding|false|false||end
null|ENG gene|Finding|false|false||end
null|ENG wt Allele|Finding|false|false||endnull|Stop (qualifier value)|Time|false|false||endnull|End|Modifier|false|false||endnull|Long Variable|Modifier|false|false||long
null|Long|Modifier|false|false||longnull|Sentence|Finding|false|false||sentencenull|Basilar Rales|Finding|false|false||crackles
null|Rales|Finding|false|false||cracklesnull|Malignant neoplasm of thorax|Disorder|false|false||thoraxnull|Chest|Anatomy|false|false||thoraxnull|diffuse wheezing|Finding|false|false||diffuse wheezingnull|Diffuse|Modifier|false|false||diffusenull|Wheezing|Finding|false|false||wheezingnull|Malignant neoplasm of abdomen|Disorder|false|false||ABDOMENnull|Abdomen problem|Finding|false|false||ABDOMENnull|Abdomen|Anatomy|false|false||ABDOMEN
null|Abdominal Cavity|Anatomy|false|false||ABDOMENnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|LRRC4B gene|Finding|true|false||HSMnull|Emotional tenderness|Finding|true|false||tenderness
null|Sore to touch|Finding|true|false||tendernessnull|All extremities|Anatomy|false|false||EXTREMITIES
null|Limb structure|Anatomy|false|false||EXTREMITIESnull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Shin|Anatomy|false|false||shinsnull|Femur|Anatomy|false|false||femoralnull|Bruit|Finding|true|false||bruitsnull|null|Drug|false|false||PULSESnull|Physiologic pulse|Finding|false|false||PULSESnull|Pulse taking|Procedure|false|false||PULSESnull|Distal Resection Margin|Attribute|false|false||Distalnull|Distal (qualifier value)|Modifier|false|false||Distalnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Palpable|Modifier|false|false||palpablenull|Symmetric Relationship|Finding|false|false||symmetric
null|Symmetrical|Finding|false|false||symmetricnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|physical examination (physical finding)|Finding|false|false||PHYSICAL EXAMINATIONnull|Physical Examination|Procedure|false|false||PHYSICAL EXAMINATIONnull|physical examination (physical finding)|Finding|false|false||PHYSICAL
null|Physical|Finding|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||EXAMINATION
null|Medical Examination|Procedure|false|false||EXAMINATIONnull|Examination|Event|false|false||EXAMINATIONnull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GENERALnull|General medical service|Procedure|false|false||GENERALnull|Generalized|Modifier|false|false||GENERALnull|Obesity|Disorder|false|false||obesenull|Sitting upright|Finding|false|false||sitting uprightnull|Special Handling Code - Upright|Finding|false|false||uprightnull|Entity Handling - upright|Phenomenon|false|false||uprightnull|Upright|Modifier|false|false||uprightnull|BORNHOLM EYE DISEASE|Disorder|false|false||bednull|Bachelor of Education|Finding|false|false||bednull|Beds|Device|false|false||bednull|Patient Location - Bed|Modifier|false|false||bednull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|Mood (psychological function)|Finding|false|false||Mood
null|mood (physical finding)|Finding|false|false||Mood
null|Mood (attribute)|Finding|false|false||Moodnull|null|Attribute|false|false||Moodnull|Appropriate|Modifier|false|false||appropriatenull|HEENT|Anatomy|false|false||HEENTnull|Scleral Diseases|Disorder|false|false||Scleranull|examination of sclera|Procedure|false|false||Scleranull|Sclera|Anatomy|false|false||Scleranull|Anicteric|Finding|false|false||anictericnull|Pupil equal round and reacting to light|Finding|false|false||PERRLnull|Malignant neoplasm of conjunctiva|Disorder|false|false||Conjunctiva
null|Benign neoplasm of conjunctiva|Disorder|false|false||Conjunctiva
null|Conjunctival Diseases|Disorder|false|false||Conjunctivanull|Specimen Type - Conjunctiva|Finding|false|false||Conjunctiva
null|null|Finding|false|false||Conjunctivanull|examination of conjunctiva|Procedure|false|false||Conjunctiva
null|Procedure on conjunctiva|Procedure|false|false||Conjunctivanull|Structure of palpebral conjunctiva|Anatomy|false|false||Conjunctiva
null|conjunctiva|Anatomy|false|false||Conjunctivanull|Pink color|Modifier|false|false||pinknull|Pallor of skin|Finding|true|false||pallornull|Cyanosis|Finding|true|false||cyanosisnull|Oral mucous membrane structure|Anatomy|false|false||oral mucosanull|Oral Dosage Form|Drug|false|false||oralnull|Oral Route of Administration|Finding|false|false||oral
null|Oral (intended site)|Finding|false|false||oralnull|Oral cavity|Anatomy|false|false||oralnull|Oral|Modifier|false|false||oralnull|null|Finding|false|false||mucosanull|Mucous Membrane|Anatomy|false|false||mucosanull|Passive joint movement of neck (finding)|Finding|false|false||NECK
null|Neck problem|Finding|false|false||NECKnull|dendritic spine neck|Anatomy|false|false||NECK
null|Neck|Anatomy|false|false||NECKnull|Supple|Finding|false|false||Supplenull|Jugular venous pressure|Finding|false|false||JVPnull|Cardiac attachment|Finding|false|false||CARDIACnull|Heart|Anatomy|false|false||CARDIACnull|Cardiac - anatomy qualifier|Modifier|false|false||CARDIACnull|Point of Maximum Impulse|Finding|false|false||PMI
null|TMEM11 gene|Finding|false|false||PMI
null|PMM2 wt Allele|Finding|false|false||PMI
null|PMM2 gene|Finding|false|false||PMI
null|MPI gene|Finding|false|false||PMInull|Prostate Mechanical Imager|Device|false|false||PMInull|Space of intercostal compartment|Anatomy|false|false||intercostal space
null|Structure of intercostal space|Anatomy|false|false||intercostal spacenull|Intercostal|Modifier|false|false||intercostalnull|Space (Astronomy)|Phenomenon|false|false||spacenull|Space - property|Modifier|false|false||spacenull|Midclavicular|Modifier|false|false||midclavicularnull|Line Specimen|Drug|false|false||line
null|Long Interspersed Elements|Drug|false|false||line
null|Long Interspersed Elements|Drug|false|false||linenull|line source specimen code|Finding|false|false||linenull|Intravascular line|Device|false|false||linenull|Linear|Modifier|false|false||linenull|Line Unit of Length|LabModifier|false|false||linenull|Heart murmur|Finding|true|false||murmursnull|Pericardial friction rub|Finding|true|false||rubsnull|Cardiac thrill (finding)|Finding|false|false||thrillsnull|hoist [device]|Device|false|false||liftsnull|Lung|Anatomy|false|false||LUNGSnull|Respiratory, thoracic and mediastinal disorders|Disorder|false|false||Respnull|Respiratory rate|Attribute|false|false||Respnull|Unlabored|Finding|false|false||unlaborednull|Use of accessory muscles|Finding|true|false||accessory muscle usenull|Accessory skeletal muscle|Disorder|true|false||accessory musclenull|Accessory|Device|true|false||accessorynull|Muscle (organ)|Anatomy|false|false||muscle
null|Muscle Tissue|Anatomy|false|false||musclenull|Use - dosing instruction imperative|Finding|true|false||use
null|utilization qualifier|Finding|true|false||use
null|Usage|Finding|true|false||usenull|Basilar Rales|Finding|false|false||crackles
null|Rales|Finding|false|false||cracklesnull|Sequence Chromatogram|Finding|false|false||tracenull|Trace Dosing Unit|LabModifier|false|false||trace
null|trace amount|LabModifier|false|false||trace
null|unknown - trace|LabModifier|false|false||tracenull|diffuse wheezing|Finding|false|false||diffuse wheezingnull|Diffuse|Modifier|false|false||diffusenull|Wheezing|Finding|false|false||wheezingnull|Malignant neoplasm of abdomen|Disorder|false|false||ABDOMENnull|Abdomen problem|Finding|false|false||ABDOMENnull|Abdomen|Anatomy|false|false||ABDOMEN
null|Abdominal Cavity|Anatomy|false|false||ABDOMENnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|LRRC4B gene|Finding|true|false||HSMnull|Emotional tenderness|Finding|true|false||tenderness
null|Sore to touch|Finding|true|false||tendernessnull|All extremities|Anatomy|false|false||EXTREMITIES
null|Limb structure|Anatomy|false|false||EXTREMITIESnull|Femur|Anatomy|false|false||femoralnull|Bruit|Finding|true|false||bruitsnull|null|Drug|false|false||PULSESnull|Physiologic pulse|Finding|false|false||PULSESnull|Pulse taking|Procedure|false|false||PULSESnull|Distal Resection Margin|Attribute|false|false||Distalnull|Distal (qualifier value)|Modifier|false|false||Distalnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Palpable|Modifier|false|false||palpablenull|Symmetric Relationship|Finding|false|false||symmetric
null|Symmetrical|Finding|false|false||symmetricnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Lymph|Finding|false|false||Lymphsnull|Monos|Drug|false|false||Monos
null|Mono-S|Drug|false|false||Monos
null|Monos|Drug|false|false||Monosnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||Eos
null|Familial eosinophilia|Disorder|false|false||Eosnull|PRSS33 gene|Finding|false|false||Eos
null|IKZF4 gene|Finding|false|false||Eosnull|Eos <Loriini>|Entity|false|false||Eosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|RET protein, human|Drug|false|false||Retnull|RET protein, human|Finding|false|false||Ret
null|RET gene|Finding|false|false||Ret
null|Oncogene RET|Finding|false|false||Ret
null|RET wt Allele|Finding|false|false||Retnull|ret unit of radiation dose|LabModifier|false|false||Retnull|CONSTRICTING BANDS, CONGENITAL|Disorder|false|false||Abs
null|Amniotic Band Syndrome|Disorder|false|false||Absnull|DDX41 wt Allele|Finding|false|false||Abs
null|DDX41 gene|Finding|false|false||Absnull|RET protein, human|Drug|false|false||Retnull|RET protein, human|Finding|false|false||Ret
null|RET gene|Finding|false|false||Ret
null|Oncogene RET|Finding|false|false||Ret
null|RET wt Allele|Finding|false|false||Retnull|ret unit of radiation dose|LabModifier|false|false||Retnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MB
null|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MBnull|creatine kinase activity|Finding|false|false||CK-MBnull|Serum creatine phosphokinase MB isoenzyme measurement|Procedure|false|false||CK-MB
null|Creatine kinase MB measurement|Procedure|false|false||CK-MBnull|MB-6|Drug|false|false||MB-6null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MB
null|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MBnull|creatine kinase activity|Finding|false|false||CK-MBnull|Serum creatine phosphokinase MB isoenzyme measurement|Procedure|false|false||CK-MB
null|Creatine kinase MB measurement|Procedure|false|false||CK-MBnull|MB-6|Drug|false|false||MB-6null|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Imaging problem|Finding|false|false||IMAGINGnull|Diagnostic Imaging|Procedure|false|false||IMAGING
null|Imaging Techniques|Procedure|false|false||IMAGINGnull|Imaging Technology|Title|false|false||IMAGINGnull|Plain chest X-ray|Procedure|false|false||CXRnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Pulmonary Edema|Finding|false|false||pulmonary edemanull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Protein Domain|Drug|false|false||regionnull|Geographic Locations|Entity|false|false||regionnull|regional|Modifier|false|false||regionnull|More|LabModifier|false|false||morenull|Confluent|Modifier|false|false||confluentnull|Lung consolidation|Disorder|false|false||consolidationnull|Consolidation|Modifier|false|false||consolidationnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|Possible|Finding|false|false||possiblenull|Possible diagnosis|Modifier|false|false||possible
null|Possibly Related to Intervention|Modifier|false|false||possiblenull|Small|LabModifier|false|false||smallnull|Bilateral|Modifier|false|false||bilateralnull|Pleural effusion (disorder)|Finding|false|false||pleural effusionsnull|Pleural Diseases|Disorder|false|false||pleuralnull|Pleura|Anatomy|false|false||pleuralnull|Pleural|Modifier|false|false||pleuralnull|effusion|Finding|false|false||effusionsnull|Moderate - Severity of Illness Code|Finding|false|false||Moderate
null|Moderate|Finding|false|false||Moderatenull|Moderate (severity modifier)|Modifier|false|false||Moderate
null|Moderate - Allergy Severity|Modifier|false|false||Moderate
null|Moderation|Modifier|false|false||Moderatenull|Cardiomegaly|Finding|false|false||cardiomegalynull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Tortuosity|Modifier|false|false||tortuositynull|Descending thoracic aorta|Anatomy|false|false||descending thoracic aorta
null|Thoracic aorta|Anatomy|false|false||descending thoracic aortanull|Sequencing - Descending|Finding|false|false||descendingnull|Descending|Modifier|false|false||descendingnull|Chest>Aorta.thoracic|Anatomy|false|false||thoracic aorta
null|Thoracic aorta|Anatomy|false|false||thoracic aortanull|Dissecting Thoracic Aortic Aneurysm|Disorder|false|false||thoracicnull|Chest|Anatomy|false|false||thoracicnull|Procedure on aorta|Procedure|false|false||aortanull|Chest+Abdomen>Aorta|Anatomy|false|false||aorta
null|Aorta|Anatomy|false|false||aortanull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|false|false||acutenull|Bone Tissue, Human|Anatomy|false|false||osseous
null|Skeletal bone|Anatomy|false|false||osseousnull|Congenital Abnormality|Disorder|true|false||abnormalitiesnull|teratologic|Finding|true|false||abnormalitiesnull|Mild Severity of Illness Code|Finding|false|false||Mildnull|Mild (qualifier value)|Modifier|false|false||Mild
null|Mild Allergy Severity|Modifier|false|false||Mildnull|Pulmonary Edema|Finding|false|false||pulmonary edemanull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|Lung consolidation|Disorder|false|false||consolidationnull|Consolidation|Modifier|false|false||consolidationnull|More|LabModifier|false|false||morenull|Confluent|Modifier|false|false||confluentnull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Old|Time|false|false||oldnull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|null|Finding|false|false||history of hypertensionnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Hypertensive disease|Disorder|false|false||hypertensionnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|DES protein, human|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|DES protein, human|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DESnull|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|Disorder|false|false||DESnull|DES gene|Finding|false|false||DESnull|Ischemic|Finding|false|false||ischemicnull|Systolic dysfunction|Finding|false|false||systolic dysfunctionnull|Systole|Finding|false|false||systolicnull|DYSFUNCTION - SKIN DISORDERS|Disorder|false|false||dysfunctionnull|Dysfunction|Finding|false|false||dysfunction
null|physiopathological|Finding|false|false||dysfunction
null|Functional disorder|Finding|false|false||dysfunctionnull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|Congestive heart failure|Disorder|false|false||CHFnull|Choroidal fissure|Anatomy|false|false||CHFnull|Exacerbation|Finding|false|false||exacerbationnull|Acute-on-chronic|Time|false|false||Acute on chronicnull|Admission Level of Care Code - Acute|Finding|false|false||Acute
null|Acute - Triage Code|Finding|false|false||Acutenull|acute|Time|false|false||Acutenull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Decompensated cardiac failure|Disorder|false|false||decompensated heart failurenull|Decompensated|Modifier|false|false||decompensatednull|Congestive heart failure|Disorder|false|false||heart failure
null|Heart failure|Disorder|false|false||heart failurenull|Malignant neoplasm of heart|Disorder|false|false||heart
null|benign neoplasm of heart|Disorder|false|false||heartnull|HEART PROBLEM|Finding|false|false||heartnull|Chest>Heart|Anatomy|false|false||heart
null|Heart|Anatomy|false|false||heartnull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Sodium Chloride, Dietary|Drug|false|false||salt
null|sodium chloride|Drug|false|false||salt
null|Salts|Drug|false|false||saltnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Dyspnea on exertion|Finding|false|false||dyspnea on exertionnull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|Exertion|Finding|false|false||exertionnull|null|Finding|false|false||exercise tolerancenull|null|Attribute|false|false||exercise tolerance
null|Exercise Tolerance|Attribute|false|false||exercise tolerancenull|Exercise|Finding|false|false||exercisenull|Exercise Pain Management|Procedure|false|false||exercisenull|Physiologic tolerance|Finding|false|false||tolerance
null|Mental tolerance|Finding|false|false||tolerance
null|Immune Tolerance|Finding|false|false||tolerance
null|Drug Tolerance|Finding|false|false||tolerancenull|Tolerance|Modifier|false|false||tolerancenull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Basilar Rales|Finding|false|false||crackles
null|Rales|Finding|false|false||cracklesnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Elevated|Modifier|false|false||elevated
null|High|Modifier|false|false||elevatednull|NPPB protein, human|Drug|false|false||BNP
null|NPPB protein, human|Drug|false|false||BNP
null|nesiritide|Drug|false|false||BNP
null|nesiritide|Drug|false|false||BNP
null|nesiritide|Drug|false|false||BNPnull|NPPB wt Allele|Finding|false|false||BNP
null|NPPB gene|Finding|false|false||BNPnull|Brain natriuretic peptide measurement|Procedure|false|false||BNPnull|Dry body weight (observable entity)|Subject|false|false||dry weightnull|dry weight (physical finding)|LabModifier|false|false||dry weightnull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|Pulmonary congestion|Disorder|false|false||pulmonary congestionnull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Congestion|Finding|false|false||congestionnull|Plain chest X-ray|Procedure|false|false||CXRnull|Late|Time|false|false||Laternull|Diagnostic Service Section ID - Pharmacy|Finding|false|false||pharmacy
null|Pharmacy domain|Finding|false|false||pharmacynull|Pharmaceutical Services|Procedure|false|false||pharmacynull|Pharmacy facility|Device|false|false||pharmacynull|Pharmacy (field)|Title|false|false||pharmacynull|Pharmacy facility|Entity|false|false||pharmacynull|Review (Publication Type)|Finding|false|false||review
null|Act Class - review|Finding|false|false||reviewnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|torsemide|Drug|false|false||torsemide
null|torsemide|Drug|false|false||torsemidenull|Last|Modifier|false|false||lastnull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Cardiovascular system|Anatomy|false|false||Cardiologynull|cardiology (field)|Title|false|false||Cardiologynull|Cardiology service|Entity|false|false||Cardiologynull|Appointments|Event|false|false||appointmentnull|Troponin|Drug|false|false||Troponins
null|Troponin|Drug|false|false||Troponinsnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|On admission|Time|false|false||On admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Sodium Chloride, Dietary|Drug|false|false||salt
null|sodium chloride|Drug|false|false||salt
null|Salts|Drug|false|false||saltnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Dietary Restriction|Procedure|false|false||restricted dietnull|Document Confidentiality Status - Restricted|Finding|false|false||restricted
null|Confidentiality - restricted|Finding|false|false||restricted
null|Confidentiality code - Restricted|Finding|false|false||restricted
null|Restricted|Finding|false|false||restrictednull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Lasix|Drug|false|false||Lasix
null|Lasix|Drug|false|false||Lasixnull|2 Days|Time|false|false||2 daysnull|day|Time|false|false||daysnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|torsemide|Drug|false|false||torsemide
null|torsemide|Drug|false|false||torsemidenull|Steady|Modifier|false|false||steadynull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|Ephrin Type-B Receptor 1, human|Drug|false|false||net
null|SLC6A2 protein, human|Drug|false|false||net
null|SLC6A2 protein, human|Drug|false|false||net
null|Ephrin Type-B Receptor 1, human|Drug|false|false||netnull|NET questionnaire|Finding|false|false||net
null|SLC6A2 gene|Finding|false|false||net
null|SLC6A2 wt Allele|Finding|false|false||net
null|EPHB1 wt Allele|Finding|false|false||net
null|ELK3 wt Allele|Finding|false|false||net
null|ELK3 gene|Finding|false|false||net
null|EPHB1 gene|Finding|false|false||net
null|Ephrin Type-B Receptor 1, human|Finding|false|false||netnull|Neutrophil Extracellular Traps|Anatomy|false|false||netnull|Net (qualifier)|Modifier|false|false||netnull|Negative fluid balance|Finding|false|false||negative fluid balancenull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Fluid Balance|Finding|false|false||fluid balancenull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Balance (substance)|Drug|false|false||balance
null|Balance (substance)|Drug|false|false||balancenull|Ability to balance|Finding|false|false||balance
null|Equilibrium|Finding|false|false||balancenull|examination of balance|Procedure|false|false||balancenull|balance device|Device|false|false||balancenull|Balanced (qualifier value)|Modifier|false|false||balancenull|objective (goal)|Finding|false|false||goal
null|Act Mood - Goal|Finding|false|false||goalnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Renal function|Finding|false|false||renal functionnull|Kidney Function Tests|Procedure|false|false||renal functionnull|Urologic Diseases|Disorder|false|false||renalnull|Kidney|Anatomy|false|false||renalnull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|Electrolytes|Drug|false|false||Electrolytes
null|Electrolytes|Drug|false|false||Electrolytes
null|Electrolyte [EPC]|Drug|false|false||Electrolytesnull|objective (goal)|Finding|false|false||goal
null|Act Mood - Goal|Finding|false|false||goalnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|carvedilol|Drug|false|false||carvedilol
null|carvedilol|Drug|false|false||carvedilolnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|atorvastatin|Drug|false|false||atorvastatin
null|atorvastatin|Drug|false|false||atorvastatinnull|Daily|Time|false|false||dailynull|lisinopril|Drug|false|false||lisinopril
null|lisinopril|Drug|false|false||lisinoprilnull|Daily|Time|false|false||dailynull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Control brand of phenylpropanolamine|Drug|false|false||control
null|CONTROL veterinary product|Drug|false|false||control
null|control substance|Drug|false|false||control
null|Control brand of phenylpropanolamine|Drug|false|false||controlnull|Control - Relationship modifier|Finding|false|false||control
null|Control function|Finding|false|false||control
null|Scientific Control|Finding|false|false||controlnull|Control Groups|Subject|false|false||controlnull|True Control Status|Modifier|false|false||control
null|control aspects|Modifier|false|false||controlnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|nifedipine|Drug|false|false||nifedipine
null|nifedipine|Drug|false|false||nifedipinenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|objective (goal)|Finding|false|false||goal
null|Act Mood - Goal|Finding|false|false||goalnull|Androgen Binding Protein|Drug|false|false||SBP
null|Androgen Binding Protein|Drug|false|false||SBPnull|CCHCR1 wt Allele|Finding|false|false||SBP
null|SHBG wt Allele|Finding|false|false||SBPnull|Systolic blood pressure measurement|Procedure|false|false||SBPnull|Systolic Pressure|Attribute|false|false||SBPnull|Close|Finding|false|false||close
null|Closed|Finding|false|false||closenull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Weights - exercise activity|Finding|false|false||weightsnull|Weight|LabModifier|false|false||weightsnull|Blood pressure finding|Finding|false|false||blood pressure
null|Systemic arterial pressure|Finding|false|false||blood pressure
null|Blood Pressure|Finding|false|false||blood pressurenull|Blood pressure determination|Procedure|false|false||blood pressurenull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Control brand of phenylpropanolamine|Drug|false|false||control
null|CONTROL veterinary product|Drug|false|false||control
null|control substance|Drug|false|false||control
null|Control brand of phenylpropanolamine|Drug|false|false||controlnull|Control - Relationship modifier|Finding|false|false||control
null|Control function|Finding|false|false||control
null|Scientific Control|Finding|false|false||controlnull|Control Groups|Subject|false|false||controlnull|True Control Status|Modifier|false|false||control
null|control aspects|Modifier|false|false||controlnull|Hypertensive disease|Disorder|false|false||Hypertensionnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|carvedilol|Drug|false|false||carvedilol
null|carvedilol|Drug|false|false||carvedilolnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|atorvastatin|Drug|false|false||atorvastatin
null|atorvastatin|Drug|false|false||atorvastatinnull|Daily|Time|false|false||dailynull|lisinopril|Drug|false|false||lisinopril
null|lisinopril|Drug|false|false||lisinoprilnull|Daily|Time|false|false||dailynull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Control brand of phenylpropanolamine|Drug|false|false||control
null|CONTROL veterinary product|Drug|false|false||control
null|control substance|Drug|false|false||control
null|Control brand of phenylpropanolamine|Drug|false|false||controlnull|Control - Relationship modifier|Finding|false|false||control
null|Control function|Finding|false|false||control
null|Scientific Control|Finding|false|false||controlnull|Control Groups|Subject|false|false||controlnull|True Control Status|Modifier|false|false||control
null|control aspects|Modifier|false|false||controlnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|nifedipine|Drug|false|false||nifedipine
null|nifedipine|Drug|false|false||nifedipinenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|objective (goal)|Finding|false|false||goal
null|Act Mood - Goal|Finding|false|false||goalnull|Androgen Binding Protein|Drug|false|false||SBP
null|Androgen Binding Protein|Drug|false|false||SBPnull|CCHCR1 wt Allele|Finding|false|false||SBP
null|SHBG wt Allele|Finding|false|false||SBPnull|Systolic blood pressure measurement|Procedure|false|false||SBPnull|Systolic Pressure|Attribute|false|false||SBPnull|BRAF Gene Rearrangement|Disorder|false|false||Positivenull|Rh Positive Blood Group|Finding|false|false||Positive
null|Positive Finding|Finding|false|false||Positive
null|Positive|Finding|false|false||Positivenull|Positive Charge|Modifier|false|false||Positivenull|Positive Number|LabModifier|false|false||Positivenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Asymptomatic diagnosis of|Finding|false|false||asymptomatic
null|Asymptomatic (finding)|Finding|false|false||asymptomaticnull|bacteria aspects|Finding|false|false||bacterianull|Bacteria <walking sticks>|Entity|false|false||bacteria
null|Bacteria|Entity|false|false||bacterianull|Asymptomatic diagnosis of|Finding|false|false||Asymptomatic
null|Asymptomatic (finding)|Finding|false|false||Asymptomaticnull|Fever|Finding|false|false||feversnull|Dysuria|Finding|false|false||dysurianull|Malaise|Finding|false|false||malaisenull|Culture urine negative|Lab|false|false||Urine culture negativenull|Urine culture|Procedure|false|false||Urine culturenull|Portion of urine|Finding|false|false||Urine
null|null|Finding|false|false||Urine
null|Urine|Finding|false|false||Urine
null|In Urine|Finding|false|false||Urine
null|Urine specimen|Finding|false|false||Urinenull|Culture negative|Lab|false|false||culture negativenull|Culture Dose Form|Drug|false|false||culturenull|Culture (Anthropological)|Finding|false|false||culture
null|Cultural aspects|Finding|false|false||culturenull|Microbial culture (procedure)|Procedure|false|false||culture
null|Laboratory culture|Procedure|false|false||culturenull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Lung consolidation|Disorder|false|false||lung consolidationnull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|Lung consolidation|Disorder|false|false||consolidationnull|Consolidation|Modifier|false|false||consolidationnull|Administration Method - Infiltrate|Finding|false|false||infiltrate
null|null|Finding|false|false||infiltrate
null|Infiltration|Finding|false|false||infiltratenull|radiology referral type|Finding|false|false||Radiology
null|Radiology Section ID|Finding|false|false||Radiology
null|Encounter due to radiological examination|Finding|false|false||Radiologynull|Radiology studies|Procedure|false|false||Radiology
null|Diagnostic radiologic examination|Procedure|false|false||Radiology
null|Radiographic imaging procedure|Procedure|false|false||Radiologynull|Radiology Specialty|Title|false|false||Radiologynull|Reading (datum presentation)|Finding|false|false||read
null|Do Reading Question|Finding|false|false||read
null|Reading (activity)|Finding|false|false||readnull|Nucleotide Sequence Read|Procedure|false|false||readnull|On admission|Time|false|false||on admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Plain chest X-ray|Procedure|false|false||CXRnull|Cough (guaifenesin)|Drug|true|false||cough
null|Cough (guaifenesin)|Drug|true|false||coughnull|Coughing|Finding|true|false||coughnull|Fever|Finding|true|false||feversnull|Leukocytosis|Disorder|true|false||leukocytosisnull|Blood leukocyte number above reference range|Finding|true|false||leukocytosisnull|Call - dosing instruction fragment|Finding|false|false||call
null|Call (Instruction)|Finding|false|false||call
null|Decision|Finding|false|false||call
null|CHL1 gene|Finding|false|false||callnull|Procedure Practitioner Identifier Code Type - Radiologist|Finding|false|false||radiologistnull|radiologist|Subject|false|false||radiologistnull|Pulmonary Edema|Finding|false|false||pulmonary edemanull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Repeat Object|Finding|false|false||repeat
null|Repeat|Finding|false|false||repeatnull|Repeat Pattern|Time|false|false||repeatnull|Imaging problem|Finding|false|false||imagingnull|Diagnostic Imaging|Procedure|false|false||imaging
null|Imaging Techniques|Procedure|false|false||imagingnull|Imaging Technology|Title|false|false||imagingnull|Peptide Nucleic Acids|Drug|false|false||PNAnull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Signs and Symptoms|Finding|true|false||clinical findingsnull|Clinical NEC (not elsewhere classified in LNC)|Finding|false|false||clinicalnull|Clinical|Modifier|false|false||clinicalnull|findings aspects|Finding|true|false||findingsnull|null|Attribute|true|false||findingsnull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|Coumadin|Drug|false|false||Coumadin
null|Coumadin|Drug|false|false||Coumadinnull|objective (goal)|Finding|false|false||goal
null|Act Mood - Goal|Finding|false|false||goalnull|Aspects of signs|Finding|true|false||signs
null|Physical findings|Finding|true|false||signsnull|Manufactured sign|Device|true|false||signsnull|Thrombus|Finding|false|false||thrombus
null|Blood Clot|Finding|false|false||thrombusnull|Thrombus <Thrombidae>|Entity|false|false||thrombusnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Daily|Time|false|false||Dailynull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Coumadin|Drug|false|false||Coumadin
null|Coumadin|Drug|false|false||Coumadinnull|Daily|Time|false|false||dailynull|Anemia|Disorder|false|false||Anemianull|Anemia <Anemiaceae>|Entity|false|false||Anemianull|Aspects of signs|Finding|true|false||signs
null|Physical findings|Finding|true|false||signsnull|Manufactured sign|Device|true|false||signsnull|External route|Finding|false|false||externalnull|Body Site Modifier - External|Anatomy|false|false||externalnull|Code System Type - External|Modifier|false|false||external
null|External|Modifier|false|false||externalnull|Loss (adaptation)|Finding|true|false||lossnull|Loss (quantitative)|LabModifier|false|false||lossnull|Melena|Finding|false|false||melenanull|Anemic|Finding|false|false||anemicnull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Probable diagnosis|Finding|false|false||Likely
null|Probably|Finding|false|false||Likelynull|Kidney Diseases|Disorder|false|false||renal diseasenull|Urologic Diseases|Disorder|false|false||renalnull|Kidney|Anatomy|false|false||renalnull|Disease|Disorder|false|false||diseasenull|ACD protein, human|Drug|false|false||ACD
null|ACD protein, human|Drug|false|false||ACD
null|acid citrate dextrose|Drug|false|false||ACD
null|acid citrate dextrose|Drug|false|false||ACDnull|Anemia of chronic disease|Disorder|false|false||ACD
null|Avellino corneal dystrophy|Disorder|false|false||ACD
null|Amyloidosis cutis dyschromia|Disorder|false|false||ACD
null|Angiokeratoma Corporis Diffusum|Disorder|false|false||ACDnull|ACD gene|Finding|false|false||ACDnull|Advisory Committee to the Director, National Cancer Institute|Subject|false|false||ACDnull|Before Lunch|Time|false|false||ACDnull|Mean corpuscular volume above reference range|Finding|false|false||elevated MCVnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|Possible|Finding|false|false||possiblenull|Possible diagnosis|Modifier|false|false||possible
null|Possibly Related to Intervention|Modifier|false|false||possiblenull|Reticulocytosis|Finding|false|false||reticulocytosisnull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Suspicion|Finding|false|false||suspicionnull|Coumadin|Drug|false|false||Coumadin
null|Coumadin|Drug|false|false||Coumadinnull|Reticulocytes|Anatomy|false|false||Reticulocytesnull|Inappropriate component (foundation metadata concept)|Modifier|false|false||inappropriate
null|Inappropriate|Modifier|false|false||inappropriate
null|Inappropriate Specimen|Modifier|false|false||inappropriatenull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Loss (adaptation)|Finding|false|false||lossnull|Loss (quantitative)|LabModifier|false|false||lossnull|Daily|Time|false|false||dailynull|Complete Blood Count|Procedure|false|false||CBCnull|Nuclear cap binding complex location|Anatomy|false|false||CBCnull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|chronic kidney disease stage|Finding|false|false||Chronic kidney disease, stagenull|Chronic Kidney Diseases|Disorder|false|false||Chronic kidney diseasenull|Chronic - Admission Level of Care Code|Finding|false|false||Chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||Chronicnull|chronic|Time|false|false||Chronicnull|Kidney Diseases|Disorder|false|false||kidney diseasenull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false||kidney
null|Benign neoplasm of kidney|Disorder|false|false||kidneynull|Kidney problem|Finding|false|false||kidneynull|examination of kidney|Procedure|false|false||kidney
null|Procedures on Kidney|Procedure|false|false||kidneynull|Kidney|Anatomy|false|false||kidney
null|Both kidneys|Anatomy|false|false||kidneynull|Disease|Disorder|false|false||diseasenull|Stage level 4|Finding|false|false||stage IVnull|Tumor stage|Attribute|false|false||stagenull|Stage|Time|false|false||stage
null|Phase|Time|false|false||stagenull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Hypertensive disease|Disorder|false|false||HTNnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Changing|Finding|false|false||changenull|Change - procedure|Procedure|false|false||changenull|Delta (difference)|LabModifier|false|false||change
null|Changed status|LabModifier|false|false||changenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|atorvastatin|Drug|false|false||atorvastatin
null|atorvastatin|Drug|false|false||atorvastatinnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|insulin aspart, human|Drug|false|false||aspart
null|insulin aspart, human|Drug|false|false||aspart
null|insulin aspart, human|Drug|false|false||aspartnull|SHORT STATURE, IDIOPATHIC, X-LINKED|Disorder|false|false||ISSnull|insulin glargine|Drug|false|false||glargine
null|insulin glargine|Drug|false|false||glargine
null|insulin glargine|Drug|false|false||glarginenull|Once a day, at bedtime|Time|false|false||qHSnull|Language Ability Proficiency - Good|Finding|false|false||good
null|Language Proficiency - Good|Finding|false|false||goodnull|Specimen Quality - Good|Modifier|false|false||good
null|Good|Modifier|false|false||goodnull|Glycemic Control|Procedure|false|false||glycemic controlnull|Control brand of phenylpropanolamine|Drug|false|false||control
null|CONTROL veterinary product|Drug|false|false||control
null|control substance|Drug|false|false||control
null|Control brand of phenylpropanolamine|Drug|false|false||controlnull|Control - Relationship modifier|Finding|false|false||control
null|Control function|Finding|false|false||control
null|Scientific Control|Finding|false|false||controlnull|Control Groups|Subject|false|false||controlnull|True Control Status|Modifier|false|false||control
null|control aspects|Modifier|false|false||controlnull|Marketing basis - Transitional|Finding|false|false||TRANSITIONALnull|Transitional cell morphology|Modifier|false|false||TRANSITIONALnull|Congestive heart failure|Disorder|false|false||CHFnull|Choroidal fissure|Anatomy|false|false||CHFnull|Lasix|Drug|false|false||lasix
null|Lasix|Drug|false|false||lasixnull|Diuretics|Drug|false|false||diureticsnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|torsemide|Drug|false|false||torsemide
null|torsemide|Drug|false|false||torsemidenull|Take|Procedure|false|false||takenull|banana allergenic extract|Drug|false|false||banana
null|Banana|Drug|false|false||banana
null|banana allergenic extract|Drug|false|false||banana
null|banana extract|Drug|false|false||banana
null|banana extract|Drug|false|false||banananull|Musa x paradisiaca|Entity|false|false||banana
null|Musa acuminata|Entity|false|false||banananull|Unilateral|Modifier|false|false||unilateralnull|Document Completion - incomplete|Finding|false|false||incompletenull|Incomplete|Modifier|false|false||incompletenull|Partial|LabModifier|false|false||incompletenull|outcomes otolaryngology hearing|Finding|false|false||hearing
null|Hearing finding|Finding|false|false||hearing
null|Hearing|Finding|false|false||hearingnull|Loss (adaptation)|Finding|false|false||lossnull|Loss (quantitative)|LabModifier|false|false||lossnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Relate - vinyl resin|Drug|false|false||relatednull|Role Link Type - related|Finding|false|false||related
null|Related (finding)|Finding|false|false||relatednull|Definitely Related to Intervention|Modifier|false|false||related
null|Relationships|Modifier|false|false||relatednull|Diuretics|Drug|false|false||diureticsnull|Hypertensive disease|Disorder|false|false||HTNnull|nifedipine|Drug|false|false||nifedipine
null|nifedipine|Drug|false|false||nifedipinenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Elevated|Modifier|false|false||elevated
null|High|Modifier|false|false||elevatednull|Structure of subparietal sulcus|Anatomy|false|false||SBPsnull|next - HtmlLinkType|Finding|false|false||nextnull|Following|Time|false|false||next
null|Then|Time|false|false||nextnull|Adjacent|Modifier|false|false||nextnull|Appointments|Event|false|false||appointmentsnull|Anemia|Disorder|false|false||Anemianull|Anemia <Anemiaceae>|Entity|false|false||Anemianull|Numerous|LabModifier|false|false||multiplenull|null|Time|false|false||priornull|ACD protein, human|Drug|false|false||ACD
null|ACD protein, human|Drug|false|false||ACD
null|acid citrate dextrose|Drug|false|false||ACD
null|acid citrate dextrose|Drug|false|false||ACDnull|Angiokeratoma Corporis Diffusum|Disorder|false|false||ACD
null|Avellino corneal dystrophy|Disorder|false|false||ACD
null|Anemia of chronic disease|Disorder|false|false||ACD
null|Amyloidosis cutis dyschromia|Disorder|false|false||ACDnull|ACD gene|Finding|false|false||ACDnull|Advisory Committee to the Director, National Cancer Institute|Subject|false|false||ACDnull|Before Lunch|Time|false|false||ACDnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|null|Time|false|false||Priornull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|on warfarin|Procedure|false|false||on warfarinnull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|Continuous|Finding|false|false||continuednull|Preventive monitoring|Procedure|false|false||monitoringnull|null|Event|false|false||monitoringnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|In-House|Finding|false|false||in-housenull|House (environment)|Device|false|false||housenull|Home environment|Modifier|false|false||housenull|insulin aspart, human|Drug|false|false||aspart
null|insulin aspart, human|Drug|false|false||aspart
null|insulin aspart, human|Drug|false|false||aspartnull|insulin glargine|Drug|false|false||glargine
null|insulin glargine|Drug|false|false||glargine
null|insulin glargine|Drug|false|false||glarginenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|GDC Regimen Terminology|Finding|false|false||regimennull|Treatment Protocols|Procedure|false|false||regimennull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Accurate (qualifier value)|Modifier|false|false||accuratenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||DAILYnull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|carvedilol|Drug|false|false||Carvedilol
null|carvedilol|Drug|false|false||Carvedilolnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|gabapentin|Drug|false|false||Gabapentin
null|gabapentin|Drug|false|false||Gabapentinnull|Once a day, at bedtime|Time|false|false||QHSnull|Neuropathic pain|Finding|false|false||neuropathic pain
null|Neuralgia|Finding|false|false||neuropathic painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|lisinopril|Drug|false|false||Lisinopril
null|lisinopril|Drug|false|false||Lisinoprilnull|Daily|Time|false|false||DAILYnull|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitaminsnull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|Daily|Time|false|false||DAILYnull|nifedipine|Drug|false|false||NIFEdipine
null|nifedipine|Drug|false|false||NIFEdipinenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|nitroglycerin|Drug|false|false||Nitroglycerin
null|nitroglycerin|Drug|false|false||Nitroglycerinnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|pantoprazole|Drug|false|false||Pantoprazole
null|pantoprazole|Drug|false|false||Pantoprazolenull|Every twelve hours|Time|false|false||Q12Hnull|polyethylene glycols|Drug|false|false||Polyethylene Glycol
null|polyethylene glycols|Drug|false|false||Polyethylene Glycolnull|high-density polyethylene|Drug|false|false||Polyethylene
null|high-density polyethylene|Drug|false|false||Polyethylene
null|polyethylenes|Drug|false|false||Polyethylene
null|polyethylenes|Drug|false|false||Polyethylene
null|Polyethylene|Drug|false|false||Polyethylene
null|Polyethylene|Drug|false|false||Polyethylenenull|ethylene glycol|Drug|false|false||Glycol
null|Glycol|Drug|false|false||Glycol
null|ethylene glycol|Drug|false|false||Glycol
null|Glycols|Drug|false|false||Glycolnull|Daily|Time|false|false||DAILYnull|sennosides, USP|Drug|false|false||Senna
null|sennosides, USP|Drug|false|false||Sennanull|Senna alexandrina|Entity|false|false||Senna
null|Senna Plant|Entity|false|false||Sennanull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Constipation|Finding|false|false||constipationnull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|Storage Unit|Device|false|false||UNIT
null|Unit device|Device|false|false||UNITnull|Unit - NCI Thesaurus Property|LabModifier|false|false||UNIT
null|Unit of Measure|LabModifier|false|false||UNIT
null|Unit|LabModifier|false|false||UNIT
null|Enzyme Unit|LabModifier|false|false||UNITnull|Daily|Time|false|false||DAILYnull|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarinnull|allopurinol|Drug|false|false||Allopurinol
null|allopurinol|Drug|false|false||Allopurinolnull|Transaction counts and value totals - day|Finding|false|false||DAY
null|Precision - day|Finding|false|false||DAYnull|Land Dayak Languages|Entity|false|false||DAYnull|day|Time|false|false||DAY
null|Daily|Time|false|false||DAYnull|torsemide|Drug|false|false||Torsemide
null|torsemide|Drug|false|false||Torsemidenull|Daily|Time|false|false||DAILYnull|HumuLIN 70/30|Drug|false|false||HumuLIN 70/30
null|HumuLIN 70/30|Drug|false|false||HumuLIN 70/30
null|HumuLIN 70/30|Drug|false|false||HumuLIN 70/30null|Humulin insulin|Drug|false|false||HumuLIN
null|Humulin|Drug|false|false||HumuLIN
null|Humulin|Drug|false|false||HumuLIN
null|Humulin|Drug|false|false||HumuLIN
null|Humulin insulin|Drug|false|false||HumuLIN
null|Humulin insulin|Drug|false|false||HumuLIN
null|Humulin S|Drug|false|false||HumuLIN
null|Humulin S|Drug|false|false||HumuLIN
null|Humulin S|Drug|false|false||HumuLINnull|insulin isophane|Drug|false|false||insulin NPH
null|insulin isophane|Drug|false|false||insulin NPH
null|insulin isophane|Drug|false|false||insulin NPHnull|insulin, regular, human|Drug|false|false||insulin
null|Insulin [EPC]|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulinnull|INS gene|Finding|false|false||insulinnull|Insulin measurement|Procedure|false|false||insulinnull|Hydrocephalus, Normal Pressure|Disorder|false|false||NPHnull|Nasopharynx|Anatomy|false|false||NPHnull|Regular|Modifier|false|false||regularnull|Homo sapiens|Subject|false|false||humannull|Unit per Milliliter|LabModifier|false|false||unit/mLnull|Storage Unit|Device|false|false||unit
null|Unit device|Device|false|false||unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||unit
null|Unit of Measure|LabModifier|false|false||unit
null|Unit|LabModifier|false|false||unit
null|Enzyme Unit|LabModifier|false|false||unitnull|per milliliter|LabModifier|false|false||/mLnull|Subcutaneous Route of Administration|Finding|false|false||subcutaneousnull|subcutaneous|Modifier|false|false||subcutaneousnull|Unit - NCI Thesaurus Property|LabModifier|false|false||units
null|Unit of Measure|LabModifier|false|false||units
null|Unit|LabModifier|false|false||unitsnull|With dinner|Time|false|false||with dinnernull|Dinner|Finding|false|false||dinnernull|With dinner|Time|false|false||dinnernull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|HumuLIN 70/30|Drug|false|false||HumuLIN 70/30
null|HumuLIN 70/30|Drug|false|false||HumuLIN 70/30
null|HumuLIN 70/30|Drug|false|false||HumuLIN 70/30null|Humulin insulin|Drug|false|false||HumuLIN
null|Humulin|Drug|false|false||HumuLIN
null|Humulin|Drug|false|false||HumuLIN
null|Humulin|Drug|false|false||HumuLIN
null|Humulin insulin|Drug|false|false||HumuLIN
null|Humulin insulin|Drug|false|false||HumuLIN
null|Humulin S|Drug|false|false||HumuLIN
null|Humulin S|Drug|false|false||HumuLIN
null|Humulin S|Drug|false|false||HumuLINnull|insulin isophane|Drug|false|false||insulin NPH
null|insulin isophane|Drug|false|false||insulin NPH
null|insulin isophane|Drug|false|false||insulin NPHnull|insulin, regular, human|Drug|false|false||insulin
null|Insulin [EPC]|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulinnull|INS gene|Finding|false|false||insulinnull|Insulin measurement|Procedure|false|false||insulinnull|Hydrocephalus, Normal Pressure|Disorder|false|false||NPHnull|Nasopharynx|Anatomy|false|false||NPHnull|Regular|Modifier|false|false||regularnull|Homo sapiens|Subject|false|false||humannull|Unit per Milliliter|LabModifier|false|false||unit/mLnull|Storage Unit|Device|false|false||unit
null|Unit device|Device|false|false||unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||unit
null|Unit of Measure|LabModifier|false|false||unit
null|Unit|LabModifier|false|false||unit
null|Enzyme Unit|LabModifier|false|false||unitnull|per milliliter|LabModifier|false|false||/mLnull|Subcutaneous Route of Administration|Finding|false|false||subcutaneousnull|subcutaneous|Modifier|false|false||subcutaneousnull|Unit - NCI Thesaurus Property|LabModifier|false|false||units
null|Unit of Measure|LabModifier|false|false||units
null|Unit|LabModifier|false|false||unitsnull|With dinner|Time|false|false||with dinnernull|Dinner|Finding|false|false||dinnernull|With dinner|Time|false|false||dinnernull|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarinnull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|Storage Unit|Device|false|false||UNIT
null|Unit device|Device|false|false||UNITnull|Unit - NCI Thesaurus Property|LabModifier|false|false||UNIT
null|Unit of Measure|LabModifier|false|false||UNIT
null|Unit|LabModifier|false|false||UNIT
null|Enzyme Unit|LabModifier|false|false||UNITnull|Daily|Time|false|false||DAILYnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|allopurinol|Drug|false|false||Allopurinol
null|allopurinol|Drug|false|false||Allopurinolnull|Transaction counts and value totals - day|Finding|false|false||DAY
null|Precision - day|Finding|false|false||DAYnull|Land Dayak Languages|Entity|false|false||DAYnull|day|Time|false|false||DAY
null|Daily|Time|false|false||DAYnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||DAILYnull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|gabapentin|Drug|false|false||Gabapentin
null|gabapentin|Drug|false|false||Gabapentinnull|Once a day, at bedtime|Time|false|false||QHSnull|Neuropathic pain|Finding|false|false||neuropathic pain
null|Neuralgia|Finding|false|false||neuropathic painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|lisinopril|Drug|false|false||Lisinopril
null|lisinopril|Drug|false|false||Lisinoprilnull|Daily|Time|false|false||DAILYnull|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitaminsnull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|Daily|Time|false|false||DAILYnull|nitroglycerin|Drug|false|false||Nitroglycerin
null|nitroglycerin|Drug|false|false||Nitroglycerinnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|polyethylene glycols|Drug|false|false||Polyethylene Glycol
null|polyethylene glycols|Drug|false|false||Polyethylene Glycolnull|high-density polyethylene|Drug|false|false||Polyethylene
null|high-density polyethylene|Drug|false|false||Polyethylene
null|polyethylenes|Drug|false|false||Polyethylene
null|polyethylenes|Drug|false|false||Polyethylene
null|Polyethylene|Drug|false|false||Polyethylene
null|Polyethylene|Drug|false|false||Polyethylenenull|ethylene glycol|Drug|false|false||Glycol
null|Glycol|Drug|false|false||Glycol
null|ethylene glycol|Drug|false|false||Glycol
null|Glycols|Drug|false|false||Glycolnull|Daily|Time|false|false||DAILYnull|sennosides, USP|Drug|false|false||Senna
null|sennosides, USP|Drug|false|false||Sennanull|Senna alexandrina|Entity|false|false||Senna
null|Senna Plant|Entity|false|false||Sennanull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Constipation|Finding|false|false||constipationnull|torsemide|Drug|false|false||Torsemide
null|torsemide|Drug|false|false||Torsemidenull|Daily|Time|false|false||DAILYnull|torsemide|Drug|false|false||torsemide
null|torsemide|Drug|false|false||torsemidenull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Once daily|Time|false|false||once dailynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Daily|Time|false|false||dailynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|pantoprazole|Drug|false|false||Pantoprazole
null|pantoprazole|Drug|false|false||Pantoprazolenull|Every twelve hours|Time|false|false||Q12Hnull|carvedilol|Drug|false|false||Carvedilol
null|carvedilol|Drug|false|false||Carvedilolnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|nifedipine|Drug|false|false||NIFEdipine
null|nifedipine|Drug|false|false||NIFEdipinenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|nifedipine|Drug|false|false||nifedipine
null|nifedipine|Drug|false|false||nifedipinenull|capsule (pharmacologic)|Drug|false|false||capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||capsule
null|Structure of organ capsule|Anatomy|false|false||capsulenull|Capsule Shape|Modifier|false|false||capsulenull|Capsule (unit of presentation)|LabModifier|false|false||capsule
null|Capsule Dosing Unit|LabModifier|false|false||capsulenull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Twice a day|Time|false|false||twice dailynull|Daily|Time|false|false||dailynull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|refill|Finding|false|false||Refillsnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Acute-on-chronic|Time|false|false||Acute on chronicnull|Admission Level of Care Code - Acute|Finding|false|false||Acute
null|Acute - Triage Code|Finding|false|false||Acutenull|acute|Time|false|false||Acutenull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Decompensated|Modifier|false|false||decompensatednull|Congestive heart failure|Disorder|false|false||congestive Heart Failurenull|Congestive|Modifier|false|false||congestivenull|Congestive heart failure|Disorder|false|false||Heart Failure
null|Heart failure|Disorder|false|false||Heart Failurenull|Malignant neoplasm of heart|Disorder|false|false||Heart
null|benign neoplasm of heart|Disorder|false|false||Heartnull|HEART PROBLEM|Finding|false|false||Heartnull|Chest>Heart|Anatomy|false|false||Heart
null|Heart|Anatomy|false|false||Heartnull|Failure (biologic function)|Finding|false|false||Failure
null|Failure|Finding|false|false||Failure
null|Personal failure|Finding|false|false||Failurenull|Hypertensive disease|Disorder|false|false||Hypertensionnull|Neoplasm Metastasis|Disorder|false|false||Secondarynull|metastatic qualifier|Finding|false|false||Secondarynull|Secondary to|Modifier|false|false||Secondarynull|second (number)|LabModifier|false|false||Secondarynull|Diagnosis|Procedure|false|false||Diagnosesnull|Anemia|Disorder|false|false||Anemianull|Anemia <Anemiaceae>|Entity|false|false||Anemianull|Diabetes Mellitus|Disorder|false|false||Diabetes mellitusnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Diabetes
null|Diabetes|Disorder|false|false||Diabetes
null|Diabetes Mellitus|Disorder|false|false||Diabetesnull|null|Time|false|false||Priornull|Deep vein thrombosis of lower limb|Disorder|false|false||deep vein thrombosis
null|Deep Vein Thrombosis|Disorder|false|false||deep vein thrombosisnull|Structure of deep vein|Anatomy|false|false||deep veinnull|Deep Resection Margin|Attribute|false|false||deepnull|Deep (qualifier value)|Modifier|false|false||deepnull|Venous Thrombosis|Finding|false|false||vein thrombosisnull|Veins|Anatomy|false|false||veinnull|Thrombosis|Finding|false|false||thrombosisnull|Chronic Kidney Diseases|Disorder|false|false||Chronic Kidney Diseasenull|Chronic - Admission Level of Care Code|Finding|false|false||Chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||Chronicnull|chronic|Time|false|false||Chronicnull|Kidney Diseases|Disorder|false|false||Kidney Diseasenull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false||Kidney
null|Benign neoplasm of kidney|Disorder|false|false||Kidneynull|Kidney problem|Finding|false|false||Kidneynull|examination of kidney|Procedure|false|false||Kidney
null|Procedures on Kidney|Procedure|false|false||Kidneynull|Kidney|Anatomy|false|false||Kidney
null|Both kidneys|Anatomy|false|false||Kidneynull|Disease|Disorder|false|false||Diseasenull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|Congestive|Modifier|false|false||congestivenull|Congestive heart failure|Disorder|false|false||heart failure
null|Heart failure|Disorder|false|false||heart failurenull|Malignant neoplasm of heart|Disorder|false|false||heart
null|benign neoplasm of heart|Disorder|false|false||heartnull|HEART PROBLEM|Finding|false|false||heartnull|Chest>Heart|Anatomy|false|false||heart
null|Heart|Anatomy|false|false||heartnull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Hypertensive disease|Disorder|false|false||hypertensionnull|Diuretics|Drug|false|false||diureticsnull|Improvement|Finding|false|false||improvementnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Laboratory test finding|Lab|false|false||labsnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Blood pressure finding|Finding|false|false||blood pressure
null|Systemic arterial pressure|Finding|false|false||blood pressure
null|Blood Pressure|Finding|false|false||blood pressurenull|Blood pressure determination|Procedure|false|false||blood pressurenull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Pharmaceutical Preparations|Drug|false|false||medicinesnull|Production Class Code - Pleasure|Finding|false|false||pleasure
null|pleasurable emotion|Finding|false|false||pleasurenull|Pleasure - Animals raised for recreation|Entity|false|false||pleasurenull|care of - AddressPartType|Finding|false|false||care ofnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|NCK-Interacting Protein with SH3 Domain|Drug|false|false||wishnull|NCKIPSD wt Allele|Finding|false|false||wish
null|NCKIPSD gene|Finding|false|false||wishnull|Vitelliform Macular Dystrophy|Disorder|false|false||bestnull|BEST1 wt Allele|Finding|false|false||best
null|BEST1 gene|Finding|false|false||bestnull|best (quality)|Modifier|false|false||bestnull|Team|Subject|false|false||Teamnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions