 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|33,37
No|38,40
:|40,41
_|44,45
_|45,46
_|46,47
<EOL>|47,48
<EOL>|49,50
Admission|50,59
Date|60,64
:|64,65
_|67,68
_|68,69
_|69,70
Discharge|84,93
Date|94,98
:|98,99
_|102,103
_|103,104
_|104,105
<EOL>|105,106
<EOL>|107,108
Date|108,112
of|113,115
Birth|116,121
:|121,122
_|124,125
_|125,126
_|126,127
Sex|140,143
:|143,144
F|147,148
<EOL>|148,149
<EOL>|150,151
Service|151,158
:|158,159
MEDICINE|160,168
<EOL>|168,169
<EOL>|170,171
Allergies|171,180
:|180,181
<EOL>|182,183
Percocet|183,191
/|192,193
Vicodin|194,201
<EOL>|201,202
<EOL>|203,204
Attending|204,213
:|213,214
_|215,216
_|216,217
_|217,218
<EOL>|218,219
<EOL>|220,221
Chief|221,226
Complaint|227,236
:|236,237
<EOL>|237,238
altered|238,245
mental|246,252
status|253,259
<EOL>|259,260
<EOL>|261,262
Major|262,267
Surgical|268,276
or|277,279
Invasive|280,288
Procedure|289,298
:|298,299
<EOL>|299,300
none|300,304
<EOL>|304,305
<EOL>|306,307
History|307,314
of|315,317
Present|318,325
Illness|326,333
:|333,334
<EOL>|334,335
Mrs.|335,339
_|340,341
_|341,342
_|342,343
is|344,346
a|347,348
_|349,350
_|350,351
_|351,352
female|353,359
with|360,364
HIV|365,368
on|369,371
HAART|372,377
,|377,378
COPD|379,383
,|383,384
HCV|385,388
<EOL>|389,390
cirrhosis|390,399
complicated|400,411
by|412,414
ascites|415,422
and|423,426
hepatic|427,434
encephalopathy|435,449
who|450,453
<EOL>|454,455
initially|455,464
presented|465,474
to|475,477
the|478,481
ED|482,484
yesterday|485,494
with|495,499
hypotension|500,511
after|512,517
a|518,519
<EOL>|520,521
paracentesis|521,533
.|533,534
<EOL>|536,537
The|537,540
patient|541,548
has|549,552
had|553,556
accelerated|557,568
decompensation|569,583
of|584,586
her|587,590
cirrhosis|591,600
<EOL>|601,602
recently|602,610
with|611,615
worsening|616,625
ascites|626,633
,|633,634
and|635,638
she|639,642
is|643,645
maintained|646,656
on|657,659
twice|660,665
<EOL>|666,667
weekly|667,673
paracentesis|674,686
.|686,687
She|688,691
was|692,695
at|696,698
her|699,702
regular|703,710
session|711,718
yesterday|719,728
<EOL>|729,730
when|730,734
she|735,738
had|739,742
hypotension|743,754
to|755,757
SBP|758,761
_|762,763
_|763,764
_|764,765
and|766,769
felt|770,774
lightheadedness|775,790
.|790,791
<EOL>|792,793
Per|793,796
the|797,800
patient|801,808
,|808,809
that|810,814
's|814,816
when|817,821
her|822,825
memory|826,832
started|833,840
to|841,843
get|844,847
fuzzy|848,853
.|853,854
<EOL>|855,856
She|856,859
does|860,864
not|865,868
have|869,873
much|874,878
recollection|879,891
of|892,894
what|895,899
happened|900,908
since|909,914
then|915,919
.|919,920
<EOL>|921,922
Her|922,925
outpatient|926,936
hepatologist|937,949
saw|950,953
her|954,957
and|958,961
recommended|962,973
that|974,978
she|979,982
go|983,985
<EOL>|986,987
to|987,989
the|990,993
ED|994,996
.|996,997
In|998,1000
the|1001,1004
ED|1005,1007
,|1007,1008
she|1009,1012
was|1013,1016
evaluated|1017,1026
and|1027,1030
deemed|1031,1037
to|1038,1040
have|1041,1045
<EOL>|1046,1047
stable|1047,1053
blood|1054,1059
pressure|1060,1068
.|1068,1069
She|1070,1073
was|1074,1077
discharged|1078,1088
home|1089,1093
.|1093,1094
At|1095,1097
home|1098,1102
,|1102,1103
she|1104,1107
had|1108,1111
<EOL>|1112,1113
worsening|1113,1122
mental|1123,1129
status|1130,1136
with|1137,1141
her|1142,1145
daughter|1146,1154
getting|1155,1162
concerned|1163,1172
,|1172,1173
and|1174,1177
<EOL>|1178,1179
she|1179,1182
returned|1183,1191
to|1192,1194
the|1195,1198
ED|1199,1201
.|1201,1202
<EOL>|1204,1205
In|1205,1207
the|1208,1211
ED|1212,1214
,|1214,1215
initial|1216,1223
vitals|1224,1230
were|1231,1235
98.7|1236,1240
77|1241,1243
96|1244,1246
/|1246,1247
50|1247,1249
16|1250,1252
98|1253,1255
%|1255,1256
RA|1257,1259
.|1259,1260
The|1261,1264
<EOL>|1265,1266
patient|1266,1273
was|1274,1277
only|1278,1282
oriented|1283,1291
to|1292,1294
person|1295,1301
.|1301,1302
Her|1303,1306
labs|1307,1311
were|1312,1316
notable|1317,1324
for|1325,1328
<EOL>|1329,1330
Na|1330,1332
126|1333,1336
,|1336,1337
K|1338,1339
6.7|1340,1343
,|1343,1344
Cr|1345,1347
0.7|1348,1351
(|1352,1353
baseline|1353,1361
0.4|1362,1365
)|1365,1366
,|1366,1367
ALT|1368,1371
153|1372,1375
,|1375,1376
AST|1377,1380
275|1381,1384
,|1384,1385
TBili|1386,1391
<EOL>|1392,1393
1.9|1393,1396
,|1396,1397
Lip|1398,1401
66|1402,1404
,|1404,1405
INR|1406,1409
1.5|1410,1413
.|1413,1414
Initial|1415,1422
EKG|1423,1426
showed|1427,1433
sinus|1434,1439
rhythm|1440,1446
with|1447,1451
<EOL>|1452,1453
peaked|1453,1459
T|1460,1461
waves|1462,1467
.|1467,1468
Her|1469,1472
head|1473,1477
CT|1478,1480
was|1481,1484
negative|1485,1493
for|1494,1497
any|1498,1501
acute|1502,1507
<EOL>|1508,1509
processes|1509,1518
.|1518,1519
She|1520,1523
received|1524,1532
ceftriaxone|1533,1544
2gm|1545,1548
x1|1549,1551
,|1551,1552
regular|1553,1560
insulin|1561,1568
10U|1569,1572
,|1572,1573
<EOL>|1574,1575
calcium|1575,1582
gluconate|1583,1592
1g|1593,1595
,|1595,1596
lactulose|1597,1606
30|1607,1609
mL|1610,1612
x2|1613,1615
,|1615,1616
and|1617,1620
25g|1621,1624
5|1625,1626
%|1626,1627
albumin|1628,1635
.|1635,1636
<EOL>|1638,1639
On|1639,1641
transfer|1642,1650
,|1650,1651
vitals|1652,1658
were|1659,1663
99.0|1664,1668
93|1669,1671
84|1672,1674
/|1674,1675
40|1675,1677
16|1678,1680
95|1681,1683
%|1683,1684
NC|1685,1687
.|1687,1688
On|1689,1691
arrival|1692,1699
to|1700,1702
<EOL>|1703,1704
the|1704,1707
MICU|1708,1712
,|1712,1713
patient|1714,1721
was|1722,1725
more|1726,1730
alert|1731,1736
and|1737,1740
conversant|1741,1751
.|1751,1752
She|1753,1756
has|1757,1760
no|1761,1763
<EOL>|1764,1765
abdominal|1765,1774
pain|1775,1779
,|1779,1780
nausea|1781,1787
,|1787,1788
vomiting|1789,1797
,|1797,1798
chest|1799,1804
pain|1805,1809
,|1809,1810
or|1811,1813
difficulty|1814,1824
<EOL>|1825,1826
breathing|1826,1835
.|1835,1836
She|1837,1840
has|1841,1844
a|1845,1846
chronic|1847,1854
cough|1855,1860
that|1861,1865
is|1866,1868
not|1869,1872
much|1873,1877
changed|1878,1885
.|1885,1886
She|1887,1890
<EOL>|1891,1892
has|1892,1895
not|1896,1899
had|1900,1903
any|1904,1907
fever|1908,1913
or|1914,1916
chills|1917,1923
.|1923,1924
She|1925,1928
reports|1929,1936
taking|1937,1943
all|1944,1947
of|1948,1950
her|1951,1954
<EOL>|1955,1956
medications|1956,1967
except|1968,1974
for|1975,1978
lactulose|1979,1988
,|1988,1989
which|1990,1995
she|1996,1999
thinks|2000,2006
taste|2007,2012
<EOL>|2013,2014
disgusting|2014,2024
.|2024,2025
<EOL>|2027,2028
<EOL>|2029,2030
Past|2030,2034
Medical|2035,2042
History|2043,2050
:|2050,2051
<EOL>|2051,2052
-|2052,2053
HCV|2054,2057
Cirrhosis|2058,2067
:|2067,2068
genotype|2069,2077
3a|2078,2080
<EOL>|2082,2083
-|2083,2084
HIV|2085,2088
:|2088,2089
on|2090,2092
HAART|2093,2098
,|2098,2099
_|2100,2101
_|2101,2102
_|2102,2103
CD4|2104,2107
count|2108,2113
173|2114,2117
,|2117,2118
_|2119,2120
_|2120,2121
_|2121,2122
HIV|2123,2126
viral|2127,2132
load|2133,2137
<EOL>|2138,2139
undetectable|2139,2151
<EOL>|2153,2154
-|2154,2155
COPD|2156,2160
:|2160,2161
_|2162,2163
_|2163,2164
_|2164,2165
PFT|2166,2169
showed|2170,2176
FVC|2177,2180
1.95|2181,2185
(|2186,2187
65|2187,2189
%|2189,2190
)|2190,2191
,|2191,2192
FEV1|2193,2197
0.88|2198,2202
(|2203,2204
37|2204,2206
%|2206,2207
)|2207,2208
,|2208,2209
<EOL>|2210,2211
FEFmax|2211,2217
2.00|2218,2222
(|2223,2224
33|2224,2226
%|2226,2227
)|2227,2228
<EOL>|2230,2231
-|2231,2232
Bipolar|2233,2240
Affective|2241,2250
Disorder|2251,2259
<EOL>|2261,2262
-|2262,2263
PTSD|2264,2268
<EOL>|2270,2271
-|2271,2272
Hx|2273,2275
of|2276,2278
cocaine|2279,2286
and|2287,2290
heroin|2291,2297
abuse|2298,2303
<EOL>|2305,2306
-|2306,2307
Hx|2308,2310
of|2311,2313
skin|2314,2318
cancer|2319,2325
per|2326,2329
patient|2330,2337
report|2338,2344
<EOL>|2346,2347
<EOL>|2348,2349
Social|2349,2355
History|2356,2363
:|2363,2364
<EOL>|2364,2365
_|2365,2366
_|2366,2367
_|2367,2368
<EOL>|2368,2369
Family|2369,2375
History|2376,2383
:|2383,2384
<EOL>|2384,2385
She|2385,2388
a|2389,2390
total|2391,2396
of|2397,2399
five|2400,2404
siblings|2405,2413
,|2413,2414
but|2415,2418
she|2419,2422
is|2423,2425
not|2426,2429
talking|2431,2438
to|2439,2441
most|2442,2446
of|2447,2449
<EOL>|2450,2451
them|2451,2455
.|2455,2456
She|2457,2460
only|2461,2465
has|2466,2469
one|2470,2473
brother|2474,2481
that|2482,2486
she|2487,2490
is|2491,2493
in|2494,2496
touch|2498,2503
with|2504,2508
and|2509,2512
<EOL>|2513,2514
lives|2514,2519
in|2520,2522
_|2523,2524
_|2524,2525
_|2525,2526
.|2526,2527
She|2528,2531
is|2532,2534
not|2535,2538
aware|2539,2544
of|2545,2547
any|2548,2551
known|2552,2557
GI|2558,2560
or|2561,2563
liver|2564,2569
<EOL>|2570,2571
disease|2571,2578
in|2579,2581
her|2582,2585
family|2586,2592
.|2592,2593
<EOL>|2595,2596
<EOL>|2597,2598
Physical|2598,2606
Exam|2607,2611
:|2611,2612
<EOL>|2612,2613
ADMISSION|2613,2622
PHYSICAL|2623,2631
EXAM|2632,2636
:|2636,2637
<EOL>|2637,2638
Vitals|2638,2644
T|2645,2646
:|2646,2647
98.7|2648,2652
BP|2653,2655
:|2655,2656
84|2657,2659
/|2659,2660
48|2660,2662
P|2663,2664
:|2664,2665
91|2666,2668
R|2669,2670
:|2670,2671
24|2672,2674
O2|2675,2677
:|2677,2678
98|2679,2681
%|2681,2682
NC|2683,2685
on|2686,2688
2L|2689,2691
<EOL>|2693,2694
GENERAL|2694,2701
:|2701,2702
Alert|2703,2708
,|2708,2709
oriented|2710,2718
,|2718,2719
no|2720,2722
acute|2723,2728
distress|2729,2737
<EOL>|2739,2740
LUNGS|2740,2745
:|2745,2746
Decreased|2747,2756
air|2757,2760
movement|2761,2769
on|2770,2772
both|2773,2777
sides|2778,2783
,|2783,2784
scattered|2785,2794
<EOL>|2795,2796
expiratory|2796,2806
wheezes|2807,2814
<EOL>|2816,2817
CV|2817,2819
:|2819,2820
Regular|2821,2828
rate|2829,2833
and|2834,2837
rhythm|2838,2844
,|2844,2845
normal|2846,2852
S1|2853,2855
S2|2856,2858
,|2858,2859
no|2860,2862
murmurs|2863,2870
,|2870,2871
rubs|2872,2876
,|2876,2877
<EOL>|2878,2879
gallops|2879,2886
<EOL>|2888,2889
ABD|2889,2892
:|2892,2893
Soft|2894,2898
,|2898,2899
non-tender|2900,2910
,|2910,2911
distended|2912,2921
,|2921,2922
flank|2923,2928
dullness|2929,2937
bilaterally|2938,2949
,|2949,2950
<EOL>|2951,2952
bowel|2952,2957
sounds|2958,2964
present|2965,2972
<EOL>|2974,2975
EXT|2975,2978
:|2978,2979
Warm|2980,2984
,|2984,2985
well|2986,2990
perfused|2991,2999
,|2999,3000
2|3001,3002
+|3002,3003
pulses|3004,3010
,|3010,3011
no|3012,3014
cyanosis|3015,3023
or|3024,3026
edema|3027,3032
<EOL>|3034,3035
<EOL>|3035,3036
DISCHARGE|3036,3045
PHYSICAL|3046,3054
EXAM|3055,3059
:|3059,3060
<EOL>|3060,3061
Vitals|3061,3067
-|3067,3068
Tm|3069,3071
99.5|3072,3076
,|3076,3077
Tc|3078,3080
98.7|3081,3085
,|3085,3086
_|3087,3088
_|3088,3089
_|3089,3090
79|3091,3093
-|3093,3094
96|3094,3096
/|3096,3097
43|3097,3099
-|3099,3100
58|3100,3102
20|3103,3105
95|3106,3108
%|3108,3109
on|3110,3112
3L|3113,3115
NC|3116,3118
,|3118,3119
<EOL>|3120,3121
7BM|3121,3124
.|3124,3125
<EOL>|3127,3128
General|3128,3135
-|3135,3136
Cachectic|3137,3146
-|3146,3147
appearing|3147,3156
woman|3157,3162
,|3162,3163
alert|3164,3169
,|3169,3170
oriented|3171,3179
,|3179,3180
no|3181,3183
acute|3184,3189
<EOL>|3190,3191
distress|3191,3199
<EOL>|3201,3202
HEENT|3202,3207
-|3207,3208
Sclera|3209,3215
anicteric|3216,3225
,|3225,3226
MMM|3227,3230
,|3230,3231
oropharynx|3232,3242
clear|3243,3248
,|3248,3249
poor|3250,3254
dentition|3255,3264
<EOL>|3265,3266
with|3266,3270
partial|3271,3278
dentures|3279,3287
<EOL>|3289,3290
Neck|3290,3294
-|3294,3295
supple|3296,3302
,|3302,3303
JVP|3304,3307
not|3308,3311
elevated|3312,3320
,|3320,3321
no|3322,3324
LAD|3325,3328
<EOL>|3330,3331
Lungs|3331,3336
-|3336,3337
Clear|3338,3343
to|3344,3346
auscultation|3347,3359
bilaterally|3360,3371
,|3371,3372
no|3373,3375
wheezes|3376,3383
,|3383,3384
rales|3385,3390
,|3390,3391
<EOL>|3392,3393
ronchi|3393,3399
<EOL>|3401,3402
CV|3402,3404
-|3404,3405
Regular|3406,3413
rate|3414,3418
and|3419,3422
rhythm|3423,3429
,|3429,3430
normal|3431,3437
S1|3438,3440
+|3441,3442
S2|3443,3445
,|3445,3446
no|3447,3449
murmurs|3450,3457
,|3457,3458
rubs|3459,3463
,|3463,3464
<EOL>|3465,3466
gallops|3466,3473
<EOL>|3475,3476
Abdomen|3476,3483
-|3483,3484
Mildly|3485,3491
distended|3492,3501
and|3502,3505
firm|3506,3510
,|3510,3511
non-tender|3512,3522
,|3522,3523
bowel|3524,3529
sounds|3530,3536
<EOL>|3537,3538
present|3538,3545
,|3545,3546
no|3547,3549
rebound|3550,3557
tenderness|3558,3568
or|3569,3571
guarding|3572,3580
<EOL>|3582,3583
GU|3583,3585
-|3585,3586
no|3587,3589
foley|3590,3595
<EOL>|3597,3598
Ext|3598,3601
-|3601,3602
warm|3603,3607
,|3607,3608
well|3609,3613
perfused|3614,3622
,|3622,3623
2|3624,3625
+|3625,3626
pulses|3627,3633
,|3633,3634
no|3635,3637
clubbing|3638,3646
,|3646,3647
cyanosis|3648,3656
or|3657,3659
<EOL>|3660,3661
edema|3661,3666
<EOL>|3668,3669
Neuro|3669,3674
-|3674,3675
AOx3|3676,3680
,|3680,3681
No|3682,3684
asterixis|3685,3694
.|3694,3695
<EOL>|3697,3698
<EOL>|3699,3700
Pertinent|3700,3709
Results|3710,3717
:|3717,3718
<EOL>|3718,3719
ADMISSION|3719,3728
LABS|3729,3733
:|3733,3734
<EOL>|3734,3735
=|3735,3736
=|3736,3737
=|3737,3738
=|3738,3739
=|3739,3740
=|3740,3741
=|3741,3742
=|3742,3743
=|3743,3744
=|3744,3745
=|3745,3746
=|3746,3747
=|3747,3748
=|3748,3749
=|3749,3750
=|3750,3751
=|3751,3752
<EOL>|3752,3753
_|3753,3754
_|3754,3755
_|3755,3756
06|3757,3759
:|3759,3760
39AM|3760,3764
BLOOD|3765,3770
WBC|3771,3774
-|3774,3775
6.9|3775,3778
RBC|3779,3782
-|3782,3783
3|3783,3784
.|3784,3785
98|3785,3787
*|3787,3788
Hgb|3789,3792
-|3792,3793
14.1|3793,3797
Hct|3798,3801
-|3801,3802
41.1|3802,3806
<EOL>|3807,3808
MCV|3808,3811
-|3811,3812
103|3812,3815
*|3815,3816
MCH|3817,3820
-|3820,3821
35|3821,3823
.|3823,3824
4|3824,3825
*|3825,3826
MCHC|3827,3831
-|3831,3832
34.3|3832,3836
RDW|3837,3840
-|3840,3841
15|3841,3843
.|3843,3844
8|3844,3845
*|3845,3846
Plt|3847,3850
_|3851,3852
_|3852,3853
_|3853,3854
<EOL>|3854,3855
_|3855,3856
_|3856,3857
_|3857,3858
06|3859,3861
:|3861,3862
39AM|3862,3866
BLOOD|3867,3872
Neuts|3873,3878
-|3878,3879
72|3879,3881
.|3881,3882
7|3882,3883
*|3883,3884
Lymphs|3885,3891
-|3891,3892
14|3892,3894
.|3894,3895
7|3895,3896
*|3896,3897
Monos|3898,3903
-|3903,3904
9.8|3904,3907
<EOL>|3908,3909
Eos|3909,3912
-|3912,3913
2.5|3913,3916
Baso|3917,3921
-|3921,3922
0.3|3922,3925
<EOL>|3925,3926
_|3926,3927
_|3927,3928
_|3928,3929
06|3930,3932
:|3932,3933
39AM|3933,3937
BLOOD|3938,3943
_|3944,3945
_|3945,3946
_|3946,3947
PTT|3948,3951
-|3951,3952
32.4|3952,3956
_|3957,3958
_|3958,3959
_|3959,3960
<EOL>|3960,3961
_|3961,3962
_|3962,3963
_|3963,3964
06|3965,3967
:|3967,3968
39AM|3968,3972
BLOOD|3973,3978
Glucose|3979,3986
-|3986,3987
102|3987,3990
*|3990,3991
UreaN|3992,3997
-|3997,3998
49|3998,4000
*|4000,4001
Creat|4002,4007
-|4007,4008
0.7|4008,4011
Na|4012,4014
-|4014,4015
126|4015,4018
*|4018,4019
<EOL>|4020,4021
K|4021,4022
-|4022,4023
6|4023,4024
.|4024,4025
7|4025,4026
*|4026,4027
Cl|4028,4030
-|4030,4031
95|4031,4033
*|4033,4034
HCO3|4035,4039
-|4039,4040
25|4040,4042
AnGap|4043,4048
-|4048,4049
13|4049,4051
<EOL>|4051,4052
_|4052,4053
_|4053,4054
_|4054,4055
06|4056,4058
:|4058,4059
39AM|4059,4063
BLOOD|4064,4069
ALT|4070,4073
-|4073,4074
153|4074,4077
*|4077,4078
AST|4079,4082
-|4082,4083
275|4083,4086
*|4086,4087
AlkPhos|4088,4095
-|4095,4096
114|4096,4099
*|4099,4100
<EOL>|4101,4102
TotBili|4102,4109
-|4109,4110
1|4110,4111
.|4111,4112
9|4112,4113
*|4113,4114
<EOL>|4114,4115
_|4115,4116
_|4116,4117
_|4117,4118
06|4119,4121
:|4121,4122
39AM|4122,4126
BLOOD|4127,4132
Albumin|4133,4140
-|4140,4141
3.6|4141,4144
<EOL>|4144,4145
<EOL>|4145,4146
IMAGING|4146,4153
/|4153,4154
STUDIES|4154,4161
:|4161,4162
<EOL>|4162,4163
=|4163,4164
=|4164,4165
=|4165,4166
=|4166,4167
=|4167,4168
=|4168,4169
=|4169,4170
=|4170,4171
=|4171,4172
=|4172,4173
=|4173,4174
=|4174,4175
=|4175,4176
=|4176,4177
=|4177,4178
=|4178,4179
<EOL>|4179,4180
_|4180,4181
_|4181,4182
_|4182,4183
CT|4184,4186
HEAD|4187,4191
:|4191,4192
<EOL>|4192,4193
No|4193,4195
evidence|4196,4204
of|4205,4207
acute|4208,4213
intracranial|4214,4226
process|4227,4234
.|4234,4235
<EOL>|4235,4236
The|4236,4239
left|4240,4244
zygomatic|4245,4254
arch|4255,4259
deformity|4260,4269
is|4270,4272
probably|4273,4281
chronic|4282,4289
as|4290,4292
there|4293,4298
<EOL>|4299,4300
is|4300,4302
no|4303,4305
<EOL>|4305,4306
associated|4306,4316
soft|4317,4321
tissue|4322,4328
swelling|4329,4337
.|4337,4338
<EOL>|4338,4339
<EOL>|4339,4340
_|4340,4341
_|4341,4342
_|4342,4343
CXR|4344,4347
:|4347,4348
<EOL>|4348,4349
No|4349,4351
acute|4352,4357
intrathoracic|4358,4371
process|4372,4379
.|4379,4380
<EOL>|4380,4381
<EOL>|4381,4382
DISCHARGE|4382,4391
LABS|4392,4396
:|4396,4397
<EOL>|4397,4398
=|4398,4399
=|4399,4400
=|4400,4401
=|4401,4402
=|4402,4403
=|4403,4404
=|4404,4405
=|4405,4406
=|4406,4407
=|4407,4408
=|4408,4409
=|4409,4410
=|4410,4411
=|4411,4412
=|4412,4413
<EOL>|4413,4414
_|4414,4415
_|4415,4416
_|4416,4417
04|4418,4420
:|4420,4421
45AM|4421,4425
BLOOD|4426,4431
WBC|4432,4435
-|4435,4436
4.8|4436,4439
RBC|4440,4443
-|4443,4444
3|4444,4445
.|4445,4446
15|4446,4448
*|4448,4449
Hgb|4450,4453
-|4453,4454
11|4454,4456
.|4456,4457
2|4457,4458
*|4458,4459
Hct|4460,4463
-|4463,4464
32|4464,4466
.|4466,4467
1|4467,4468
*|4468,4469
<EOL>|4470,4471
MCV|4471,4474
-|4474,4475
102|4475,4478
*|4478,4479
MCH|4480,4483
-|4483,4484
35|4484,4486
.|4486,4487
4|4487,4488
*|4488,4489
MCHC|4490,4494
-|4494,4495
34.8|4495,4499
RDW|4500,4503
-|4503,4504
15|4504,4506
.|4506,4507
8|4507,4508
*|4508,4509
Plt|4510,4513
Ct|4514,4516
-|4516,4517
95|4517,4519
*|4519,4520
<EOL>|4520,4521
_|4521,4522
_|4522,4523
_|4523,4524
04|4525,4527
:|4527,4528
45AM|4528,4532
BLOOD|4533,4538
_|4539,4540
_|4540,4541
_|4541,4542
PTT|4543,4546
-|4546,4547
37|4547,4549
.|4549,4550
6|4550,4551
*|4551,4552
_|4553,4554
_|4554,4555
_|4555,4556
<EOL>|4556,4557
_|4557,4558
_|4558,4559
_|4559,4560
04|4561,4563
:|4563,4564
45AM|4564,4568
BLOOD|4569,4574
Glucose|4575,4582
-|4582,4583
121|4583,4586
*|4586,4587
UreaN|4588,4593
-|4593,4594
35|4594,4596
*|4596,4597
Creat|4598,4603
-|4603,4604
0.4|4604,4607
Na|4608,4610
-|4610,4611
130|4611,4614
*|4614,4615
<EOL>|4616,4617
K|4617,4618
-|4618,4619
5|4619,4620
.|4620,4621
2|4621,4622
*|4622,4623
Cl|4624,4626
-|4626,4627
97|4627,4629
HCO3|4630,4634
-|4634,4635
27|4635,4637
AnGap|4638,4643
-|4643,4644
11|4644,4646
<EOL>|4646,4647
_|4647,4648
_|4648,4649
_|4649,4650
04|4651,4653
:|4653,4654
45AM|4654,4658
BLOOD|4659,4664
ALT|4665,4668
-|4668,4669
96|4669,4671
*|4671,4672
AST|4673,4676
-|4676,4677
168|4677,4680
*|4680,4681
AlkPhos|4682,4689
-|4689,4690
69|4690,4692
TotBili|4693,4700
-|4700,4701
1|4701,4702
.|4702,4703
7|4703,4704
*|4704,4705
<EOL>|4705,4706
_|4706,4707
_|4707,4708
_|4708,4709
04|4710,4712
:|4712,4713
45AM|4713,4717
BLOOD|4718,4723
Calcium|4724,4731
-|4731,4732
8.6|4732,4735
Phos|4736,4740
-|4740,4741
2|4741,4742
.|4742,4743
4|4743,4744
*|4744,4745
Mg|4746,4748
-|4748,4749
2.|4749,4751
_|4751,4752
_|4752,4753
_|4753,4754
w|4755,4756
/|4756,4757
HIV|4758,4761
on|4762,4764
HAART|4765,4770
,|4770,4771
COPD|4772,4776
on|4777,4779
3L|4780,4782
home|4783,4787
O2|4788,4790
,|4790,4791
HCV|4792,4795
cirrhosis|4796,4805
<EOL>|4806,4807
decompensated|4807,4820
(|4821,4822
ascites|4822,4829
requiring|4830,4839
biweekly|4840,4848
therapeutic|4849,4860
<EOL>|4861,4862
paracenteses|4862,4874
,|4874,4875
hepatic|4876,4883
encephalopathy|4884,4898
;|4898,4899
not|4900,4903
on|4904,4906
transplant|4907,4917
list|4918,4922
_|4923,4924
_|4924,4925
_|4925,4926
<EOL>|4927,4928
comorbidities|4928,4941
)|4941,4942
w|4943,4944
/|4944,4945
AMS|4946,4949
,|4949,4950
hypotension|4951,4962
,|4962,4963
_|4964,4965
_|4965,4966
_|4966,4967
,|4967,4968
and|4969,4972
hyperkalemia|4973,4985
.|4985,4986
<EOL>|4987,4988
Altered|4988,4995
mental|4996,5002
status|5003,5009
improved|5010,5018
with|5019,5023
lactulose|5024,5033
.|5033,5034
Hypotension|5035,5046
was|5047,5050
<EOL>|5051,5052
felt|5052,5056
to|5057,5059
be|5060,5062
due|5063,5066
to|5067,5069
fluid|5070,5075
shifts|5076,5082
from|5083,5087
paracentesis|5088,5100
on|5101,5103
the|5104,5107
day|5108,5111
<EOL>|5112,5113
prior|5113,5118
to|5119,5121
admission|5122,5131
as|5132,5134
well|5135,5139
as|5140,5142
low|5143,5146
PO|5147,5149
intake|5150,5156
in|5157,5159
the|5160,5163
setting|5164,5171
of|5172,5174
<EOL>|5175,5176
AMS|5176,5179
.|5179,5180
Hypotension|5181,5192
and|5193,5196
_|5197,5198
_|5198,5199
_|5199,5200
resolved|5201,5209
with|5210,5214
IV|5215,5217
albumin|5218,5225
.|5225,5226
Hyperkalemia|5227,5239
<EOL>|5240,5241
resolved|5241,5249
with|5250,5254
insulin|5255,5262
and|5263,5266
kayexalate|5267,5277
.|5277,5278
<EOL>|5278,5279
<EOL>|5279,5280
#|5280,5281
Hypotension|5282,5293
:|5293,5294
Patient|5295,5302
presented|5303,5312
with|5313,5317
SBP|5318,5321
in|5322,5324
_|5325,5326
_|5326,5327
_|5327,5328
and|5329,5332
improved|5333,5341
<EOL>|5342,5343
with|5343,5347
albumin|5348,5355
in|5356,5358
the|5359,5362
ED|5363,5365
to|5366,5368
_|5369,5370
_|5370,5371
_|5371,5372
.|5372,5373
It|5374,5376
was|5377,5380
felt|5381,5385
to|5386,5388
be|5389,5391
due|5392,5395
to|5396,5398
<EOL>|5399,5400
fluid|5400,5405
shifts|5406,5412
from|5413,5417
paracentesis|5418,5430
on|5431,5433
_|5434,5435
_|5435,5436
_|5436,5437
,|5437,5438
as|5439,5441
well|5442,5446
as|5447,5449
likely|5450,5456
<EOL>|5457,5458
hypovolemia|5458,5469
given|5470,5475
AMS|5476,5479
and|5480,5483
decreased|5484,5493
PO|5494,5496
intake|5497,5503
.|5503,5504
No|5505,5507
concern|5508,5515
for|5516,5519
<EOL>|5520,5521
bleeding|5521,5529
or|5530,5532
sepsis|5533,5539
with|5540,5544
baseline|5545,5553
CBC|5554,5557
and|5558,5561
lack|5562,5566
of|5567,5569
fever|5570,5575
.|5575,5576
She|5577,5580
<EOL>|5581,5582
continued|5582,5591
to|5592,5594
received|5595,5603
IV|5604,5606
albumin|5607,5614
during|5615,5621
her|5622,5625
hospital|5626,5634
course|5635,5641
,|5641,5642
<EOL>|5643,5644
with|5644,5648
which|5649,5654
her|5655,5658
SBP|5659,5662
improved|5663,5671
to|5672,5674
_|5675,5676
_|5676,5677
_|5677,5678
and|5679,5682
patient|5683,5690
remained|5691,5699
<EOL>|5700,5701
asymptomatic|5701,5713
.|5713,5714
<EOL>|5716,5717
<EOL>|5717,5718
#|5718,5719
Hyperkalemia|5720,5732
:|5732,5733
Patient|5734,5741
presented|5742,5751
with|5752,5756
K|5757,5758
6.7|5759,5762
with|5763,5767
EKG|5768,5771
changes|5772,5779
.|5779,5780
<EOL>|5781,5782
Given|5782,5787
low|5788,5791
Na|5792,5794
,|5794,5795
likely|5796,5802
the|5803,5806
result|5807,5813
of|5814,5816
low|5817,5820
effective|5821,5830
arterial|5831,5839
volume|5840,5846
<EOL>|5847,5848
leading|5848,5855
to|5856,5858
poor|5859,5863
K|5864,5865
excretion|5866,5875
,|5875,5876
with|5877,5881
likely|5882,5888
exacerbation|5889,5901
from|5902,5906
_|5907,5908
_|5908,5909
_|5909,5910
.|5910,5911
<EOL>|5912,5913
AM|5913,5915
cortisol|5916,5924
was|5925,5928
normal|5929,5935
.|5935,5936
K|5937,5938
improved|5939,5947
with|5948,5952
insulin|5953,5960
and|5961,5964
kayexalate|5965,5975
<EOL>|5976,5977
and|5977,5980
K|5981,5982
was|5983,5986
5.2|5987,5990
on|5991,5993
day|5994,5997
of|5998,6000
discharge|6001,6010
.|6010,6011
Bactrim|6012,6019
was|6020,6023
held|6024,6028
during|6029,6035
<EOL>|6036,6037
hospital|6037,6045
course|6046,6052
.|6052,6053
<EOL>|6054,6055
<EOL>|6055,6056
#|6056,6057
_|6058,6059
_|6059,6060
_|6060,6061
:|6061,6062
Patient|6063,6070
presented|6071,6080
with|6081,6085
Cr|6086,6088
0.7|6089,6092
from|6093,6097
baseline|6098,6106
Cr|6107,6109
is|6110,6112
<EOL>|6113,6114
0.3|6114,6117
-|6117,6118
0.4|6118,6121
.|6121,6122
It|6123,6125
was|6126,6129
felt|6130,6134
to|6135,6137
be|6138,6140
likely|6141,6147
due|6148,6151
to|6152,6154
volume|6155,6161
shift|6162,6167
from|6168,6172
her|6173,6176
<EOL>|6177,6178
paracentesis|6178,6190
on|6191,6193
the|6194,6197
day|6198,6201
prior|6202,6207
to|6208,6210
admission|6211,6220
as|6221,6223
well|6224,6228
as|6229,6231
now|6232,6235
low|6236,6239
<EOL>|6240,6241
effective|6241,6250
arterial|6251,6259
volume|6260,6266
,|6266,6267
likely|6268,6274
_|6275,6276
_|6276,6277
_|6277,6278
poor|6279,6283
PO|6284,6286
intake|6287,6293
_|6294,6295
_|6295,6296
_|6296,6297
AMS|6298,6301
.|6301,6302
Cr|6303,6305
<EOL>|6306,6307
improved|6307,6315
to|6316,6318
0.4|6319,6322
with|6323,6327
albumin|6328,6335
administration|6336,6350
.|6350,6351
Furosemide|6352,6362
and|6363,6366
<EOL>|6367,6368
Bactrim|6368,6375
were|6376,6380
held|6381,6385
during|6386,6392
hospital|6393,6401
course|6402,6408
.|6408,6409
<EOL>|6412,6413
<EOL>|6413,6414
#|6414,6415
GOC|6415,6418
:|6418,6419
The|6420,6423
_|6424,6425
_|6425,6426
_|6426,6427
son|6428,6431
(|6432,6433
HCP|6433,6436
)|6436,6437
met|6438,6441
with|6442,6446
Dr.|6447,6450
_|6451,6452
_|6452,6453
_|6453,6454
<EOL>|6455,6456
outpatient|6456,6466
hepatologist|6467,6479
)|6479,6480
during|6481,6487
_|6488,6489
_|6489,6490
_|6490,6491
hospital|6492,6500
course|6501,6507
.|6507,6508
They|6509,6513
<EOL>|6514,6515
discussed|6515,6524
that|6525,6529
the|6530,6533
patient|6534,6541
is|6542,6544
not|6545,6548
a|6549,6550
transplant|6551,6561
candidate|6562,6571
<EOL>|6572,6573
givenevere|6573,6583
underlying|6584,6594
lung|6595,6599
disease|6600,6607
(|6608,6609
FEV1|6609,6613
~|6614,6615
0.8|6615,6618
)|6618,6619
,|6619,6620
hypoxia|6621,6628
,|6628,6629
RV|6630,6632
<EOL>|6633,6634
dilation|6634,6642
and|6643,6646
very|6647,6651
low|6652,6655
BMI|6656,6659
.|6659,6660
A|6661,6662
more|6663,6667
conservative|6668,6680
approach|6681,6689
was|6690,6693
<EOL>|6694,6695
recommended|6695,6706
and|6707,6710
the|6711,6714
patient|6715,6722
was|6723,6726
transitioned|6727,6739
to|6740,6742
DNR|6743,6746
/|6746,6747
DNI|6747,6750
.|6750,6751
The|6752,6755
<EOL>|6756,6757
patient|6757,6764
agreed|6765,6771
with|6772,6776
this|6777,6781
plan|6782,6786
.|6786,6787
She|6788,6791
was|6792,6795
treated|6796,6803
with|6804,6808
the|6809,6812
goal|6813,6817
of|6818,6820
<EOL>|6821,6822
treating|6822,6830
any|6831,6834
any|6835,6838
correctable|6839,6850
issues|6851,6857
.|6857,6858
Social|6859,6865
work|6866,6870
met|6871,6874
with|6875,6879
the|6880,6883
<EOL>|6884,6885
patient|6885,6892
prior|6893,6898
to|6899,6901
discharge|6902,6911
.|6911,6912
The|6913,6916
patient|6917,6924
was|6925,6928
interested|6929,6939
in|6940,6942
<EOL>|6943,6944
following|6944,6953
up|6954,6956
with|6957,6961
palliative|6962,6972
care|6973,6977
,|6977,6978
for|6979,6982
which|6983,6988
an|6989,6991
outpatient|6992,7002
<EOL>|7003,7004
referral|7004,7012
was|7013,7016
made|7017,7021
.|7021,7022
<EOL>|7023,7024
<EOL>|7025,7026
#|7026,7027
Altered|7028,7035
Mental|7036,7042
Status|7043,7049
:|7049,7050
Patient|7051,7058
presented|7059,7068
with|7069,7073
confusion|7074,7083
that|7084,7088
<EOL>|7089,7090
was|7090,7093
most|7094,7098
likely|7099,7105
secondary|7106,7115
to|7116,7118
hepatic|7119,7126
encephalopathy|7127,7141
.|7141,7142
Based|7143,7148
on|7149,7151
<EOL>|7152,7153
outpatient|7153,7163
records|7164,7171
,|7171,7172
patient|7173,7180
has|7181,7184
had|7185,7188
steady|7189,7195
decline|7196,7203
in|7204,7206
<EOL>|7207,7208
decompensated|7208,7221
cirrhosis|7222,7231
and|7232,7235
mental|7236,7242
status|7243,7249
.|7249,7250
No|7251,7253
signs|7254,7259
of|7260,7262
infection|7263,7272
<EOL>|7273,7274
and|7274,7277
head|7278,7282
CT|7283,7285
was|7286,7289
negative|7290,7298
as|7299,7301
well|7302,7306
.|7306,7307
Mental|7308,7314
status|7315,7321
improved|7322,7330
with|7331,7335
<EOL>|7336,7337
lactulose|7337,7346
in|7347,7349
the|7350,7353
ED|7354,7356
and|7357,7360
patient|7361,7368
reports|7369,7376
that|7377,7381
she|7382,7385
has|7386,7389
not|7390,7393
been|7394,7398
<EOL>|7399,7400
taking|7400,7406
lactulose|7407,7416
regularly|7417,7426
at|7427,7429
home|7430,7434
.|7434,7435
Patient|7436,7443
was|7444,7447
also|7448,7452
continued|7453,7462
<EOL>|7463,7464
on|7464,7466
rifaximin|7467,7476
.|7476,7477
<EOL>|7480,7481
<EOL>|7481,7482
#|7482,7483
HCV|7484,7487
Cirrhosis|7488,7497
:|7497,7498
Genotype|7499,7507
3a|7508,7510
.|7510,7511
Patient|7512,7519
is|7520,7522
decompensated|7523,7536
with|7537,7541
<EOL>|7542,7543
increasing|7543,7553
ascites|7554,7561
and|7562,7565
worsening|7566,7575
hepatic|7576,7583
encephalopathy|7584,7598
.|7598,7599
She|7600,7603
is|7604,7606
<EOL>|7607,7608
dependent|7608,7617
on|7618,7620
twice|7621,7626
weekly|7627,7633
paracentesis|7634,7646
.|7646,7647
Spironolactone|7648,7662
was|7663,7666
<EOL>|7667,7668
recently|7668,7676
stopped|7677,7684
due|7685,7688
to|7689,7691
hyperkalemia|7692,7704
.|7704,7705
Patient|7706,7713
is|7714,7716
not|7717,7720
a|7721,7722
<EOL>|7723,7724
transplant|7724,7734
candidate|7735,7744
given|7745,7750
her|7751,7754
comorbidities|7755,7768
COPD|7769,7773
per|7774,7777
outpatient|7778,7788
<EOL>|7789,7790
hepatologist|7790,7802
.|7802,7803
The|7804,7807
patient|7808,7815
would|7816,7821
like|7822,7826
to|7827,7829
continue|7830,7838
biweekly|7839,7847
<EOL>|7848,7849
paracenteses|7849,7861
as|7862,7864
an|7865,7867
outpatient|7868,7878
.|7878,7879
<EOL>|7879,7880
<EOL>|7880,7881
#|7881,7882
HIV|7883,7886
:|7886,7887
Most|7888,7892
recent|7893,7899
CD4|7900,7903
count|7904,7909
173|7910,7913
on|7914,7916
_|7917,7918
_|7918,7919
_|7919,7920
.|7920,7921
HIV|7922,7925
viral|7926,7931
load|7932,7936
on|7937,7939
<EOL>|7940,7941
_|7941,7942
_|7942,7943
_|7943,7944
was|7945,7948
undetectable|7949,7961
.|7961,7962
She|7963,7966
was|7967,7970
continued|7971,7980
on|7981,7983
her|7984,7987
home|7988,7992
regimen|7993,8000
<EOL>|8001,8002
of|8002,8004
raltegravir|8005,8016
,|8016,8017
emtricitabine|8018,8031
,|8031,8032
and|8033,8036
tenofovir|8037,8046
.|8046,8047
Bactrim|8048,8055
<EOL>|8056,8057
prophylaxis|8057,8068
was|8069,8072
held|8073,8077
during|8078,8084
admission|8085,8094
because|8095,8102
of|8103,8105
hyperkalemia|8106,8118
.|8118,8119
<EOL>|8122,8123
<EOL>|8123,8124
<EOL>|8124,8125
#|8125,8126
COPD|8127,8131
:|8131,8132
Patient|8133,8140
on|8141,8143
3L|8144,8146
NC|8147,8149
at|8150,8152
home|8153,8157
.|8157,8158
She|8159,8162
was|8163,8166
continued|8167,8176
on|8177,8179
her|8180,8183
home|8184,8188
<EOL>|8189,8190
regimen|8190,8197
.|8197,8198
<EOL>|8198,8199
<EOL>|8199,8200
TRANSITIONAL|8200,8212
ISSUES|8213,8219
:|8219,8220
<EOL>|8220,8221
-|8221,8222
Follow|8222,8228
up|8229,8231
with|8232,8236
Palliative|8237,8247
Care|8248,8252
as|8253,8255
outpatient|8256,8266
<EOL>|8266,8267
-|8267,8268
Bactrim|8268,8275
prophylaxis|8276,8287
(|8288,8289
HIV|8289,8292
+|8292,8293
)|8293,8294
was|8295,8298
held|8299,8303
during|8304,8310
hospital|8311,8319
course|8320,8326
due|8327,8330
<EOL>|8331,8332
to|8332,8334
_|8335,8336
_|8336,8337
_|8337,8338
.|8338,8339
Consider|8340,8348
restarting|8349,8359
as|8360,8362
outpatient|8363,8373
.|8373,8374
<EOL>|8374,8375
-|8375,8376
Furosemide|8376,8386
was|8387,8390
held|8391,8395
due|8396,8399
to|8400,8402
_|8403,8404
_|8404,8405
_|8405,8406
,|8406,8407
consider|8408,8416
restarting|8417,8427
as|8428,8430
<EOL>|8431,8432
outpatient|8432,8442
<EOL>|8442,8443
-|8443,8444
Follow|8444,8450
up|8451,8453
with|8454,8458
hepatology|8459,8469
<EOL>|8469,8470
-|8470,8471
Continue|8471,8479
biweekly|8480,8488
therapeurtic|8489,8501
paracenteses|8502,8514
<EOL>|8514,8515
-|8515,8516
Code|8516,8520
status|8521,8527
:|8527,8528
DNR|8529,8532
/|8532,8533
DNI|8533,8536
<EOL>|8536,8537
<EOL>|8538,8539
Medications|8539,8550
on|8551,8553
Admission|8554,8563
:|8563,8564
<EOL>|8564,8565
The|8565,8568
Preadmission|8569,8581
Medication|8582,8592
list|8593,8597
is|8598,8600
accurate|8601,8609
and|8610,8613
complete|8614,8622
.|8622,8623
<EOL>|8623,8624
1.|8624,8626
Lactulose|8627,8636
15|8637,8639
mL|8640,8642
PO|8643,8645
TID|8646,8649
<EOL>|8650,8651
2.|8651,8653
Tiotropium|8654,8664
Bromide|8665,8672
1|8673,8674
CAP|8675,8678
IH|8679,8681
DAILY|8682,8687
<EOL>|8688,8689
3.|8689,8691
Raltegravir|8692,8703
400|8704,8707
mg|8708,8710
PO|8711,8713
BID|8714,8717
<EOL>|8718,8719
4.|8719,8721
Emtricitabine|8722,8735
-|8735,8736
Tenofovir|8736,8745
(|8746,8747
Truvada|8747,8754
)|8754,8755
1|8756,8757
TAB|8758,8761
PO|8762,8764
DAILY|8765,8770
<EOL>|8771,8772
5.|8772,8774
Furosemide|8775,8785
40|8786,8788
mg|8789,8791
PO|8792,8794
DAILY|8795,8800
<EOL>|8801,8802
6.|8802,8804
TraMADOL|8805,8813
(|8814,8815
Ultram|8815,8821
)|8821,8822
50|8823,8825
mg|8826,8828
PO|8829,8831
Q8H|8832,8835
:|8835,8836
PRN|8836,8839
Pain|8840,8844
<EOL>|8845,8846
7.|8846,8848
Fluticasone|8849,8860
Propionate|8861,8871
110mcg|8872,8878
1|8879,8880
PUFF|8881,8885
IH|8886,8888
BID|8889,8892
<EOL>|8893,8894
8.|8894,8896
Calcium|8897,8904
Carbonate|8905,8914
500|8915,8918
mg|8919,8921
PO|8922,8924
BID|8925,8928
<EOL>|8929,8930
9.|8930,8932
Rifaximin|8933,8942
550|8943,8946
mg|8947,8949
PO|8950,8952
BID|8953,8956
<EOL>|8957,8958
10.|8958,8961
albuterol|8962,8971
sulfate|8972,8979
90|8980,8982
mcg|8983,8986
/|8986,8987
actuation|8987,8996
inhalation|8997,9007
Q6H|9008,9011
:|9011,9012
PRN|9012,9015
<EOL>|9016,9017
Wheezing|9017,9025
<EOL>|9026,9027
11.|9027,9030
Sulfameth|9031,9040
/|9040,9041
Trimethoprim|9041,9053
DS|9054,9056
1|9057,9058
TAB|9059,9062
PO|9063,9065
DAILY|9066,9071
<EOL>|9072,9073
<EOL>|9073,9074
<EOL>|9075,9076
Discharge|9076,9085
Medications|9086,9097
:|9097,9098
<EOL>|9098,9099
1|9099,9100
.|9100,9101
Calcium|9102,9109
Carbonate|9110,9119
500|9120,9123
mg|9124,9126
PO|9127,9129
BID|9130,9133
<EOL>|9134,9135
2.|9135,9137
Emtricitabine|9138,9151
-|9151,9152
Tenofovir|9152,9161
(|9162,9163
Truvada|9163,9170
)|9170,9171
1|9172,9173
TAB|9174,9177
PO|9178,9180
DAILY|9181,9186
<EOL>|9187,9188
3.|9188,9190
Fluticasone|9191,9202
Propionate|9203,9213
110mcg|9214,9220
1|9221,9222
PUFF|9223,9227
IH|9228,9230
BID|9231,9234
<EOL>|9235,9236
4.|9236,9238
Lactulose|9239,9248
30|9249,9251
mL|9252,9254
PO|9255,9257
TID|9258,9261
<EOL>|9262,9263
5.|9263,9265
Raltegravir|9266,9277
400|9278,9281
mg|9282,9284
PO|9285,9287
BID|9288,9291
<EOL>|9292,9293
6.|9293,9295
Rifaximin|9296,9305
550|9306,9309
mg|9310,9312
PO|9313,9315
BID|9316,9319
<EOL>|9320,9321
7.|9321,9323
TraMADOL|9324,9332
(|9333,9334
Ultram|9334,9340
)|9340,9341
_|9342,9343
_|9343,9344
_|9344,9345
mg|9346,9348
PO|9349,9351
Q6H|9352,9355
:|9355,9356
PRN|9356,9359
pain|9360,9364
<EOL>|9365,9366
8.|9366,9368
albuterol|9369,9378
sulfate|9379,9386
90|9387,9389
mcg|9390,9393
/|9393,9394
actuation|9394,9403
inhalation|9404,9414
Q6H|9415,9418
:|9418,9419
PRN|9419,9422
<EOL>|9423,9424
Wheezing|9424,9432
<EOL>|9433,9434
9.|9434,9436
Tiotropium|9437,9447
Bromide|9448,9455
1|9456,9457
CAP|9458,9461
IH|9462,9464
DAILY|9465,9470
<EOL>|9471,9472
<EOL>|9472,9473
<EOL>|9474,9475
Discharge|9475,9484
Disposition|9485,9496
:|9496,9497
<EOL>|9497,9498
Home|9498,9502
<EOL>|9502,9503
<EOL>|9504,9505
Discharge|9505,9514
Diagnosis|9515,9524
:|9524,9525
<EOL>|9525,9526
Primary|9526,9533
:|9533,9534
<EOL>|9534,9535
Hypotension|9535,9546
<EOL>|9546,9547
Hyperkalemia|9547,9559
<EOL>|9559,9560
Acute|9560,9565
Kidney|9566,9572
Injury|9573,9579
<EOL>|9579,9580
<EOL>|9580,9581
Secondary|9581,9590
:|9590,9591
<EOL>|9591,9592
HIV|9592,9595
<EOL>|9595,9596
Cirrhosis|9596,9605
<EOL>|9605,9606
COPD|9606,9610
<EOL>|9610,9611
<EOL>|9612,9613
Discharge|9613,9622
Condition|9623,9632
:|9632,9633
<EOL>|9633,9634
Mental|9634,9640
Status|9641,9647
:|9647,9648
Clear|9649,9654
and|9655,9658
coherent|9659,9667
.|9667,9668
<EOL>|9668,9669
Level|9669,9674
of|9675,9677
Consciousness|9678,9691
:|9691,9692
Alert|9693,9698
and|9699,9702
interactive|9703,9714
.|9714,9715
<EOL>|9715,9716
Activity|9716,9724
Status|9725,9731
:|9731,9732
Ambulatory|9733,9743
-|9744,9745
Independent|9746,9757
.|9757,9758
<EOL>|9758,9759
<EOL>|9760,9761
Discharge|9761,9770
Instructions|9771,9783
:|9783,9784
<EOL>|9784,9785
Dear|9785,9789
Ms.|9790,9793
_|9794,9795
_|9795,9796
_|9796,9797
,|9797,9798
<EOL>|9798,9799
<EOL>|9799,9800
You|9800,9803
were|9804,9808
admitted|9809,9817
to|9818,9820
_|9821,9822
_|9822,9823
_|9823,9824
because|9825,9832
of|9833,9835
confusion|9836,9845
,|9845,9846
low|9847,9850
blood|9851,9856
<EOL>|9857,9858
pressure|9858,9866
,|9866,9867
and|9868,9871
a|9872,9873
high|9874,9878
potassium|9879,9888
value|9889,9894
.|9894,9895
Your|9896,9900
confusion|9901,9910
improved|9911,9919
<EOL>|9920,9921
with|9921,9925
lactulose|9926,9935
.|9935,9936
Your|9937,9941
blood|9942,9947
pressure|9948,9956
improved|9957,9965
with|9966,9970
extra|9971,9976
fluids|9977,9983
<EOL>|9984,9985
and|9985,9988
your|9989,9993
potassium|9994,10003
improved|10004,10012
as|10013,10015
well|10016,10020
.|10020,10021
You|10022,10025
also|10026,10030
had|10031,10034
small|10035,10040
degree|10041,10047
<EOL>|10048,10049
of|10049,10051
kidney|10052,10058
injury|10059,10065
when|10066,10070
you|10071,10074
came|10075,10079
to|10080,10082
the|10083,10086
hospital|10087,10095
,|10095,10096
and|10097,10100
this|10101,10105
also|10106,10110
<EOL>|10111,10112
improved|10112,10120
with|10121,10125
fluids|10126,10132
.|10132,10133
While|10134,10139
you|10140,10143
were|10144,10148
here|10149,10153
,|10153,10154
you|10155,10158
discussed|10159,10168
<EOL>|10169,10170
changing|10170,10178
your|10179,10183
goals|10184,10189
of|10190,10192
care|10193,10197
to|10198,10200
focusing|10201,10209
on|10210,10212
symptom|10213,10220
management|10221,10231
<EOL>|10232,10233
and|10233,10236
treatment|10237,10246
of|10247,10249
reversible|10250,10260
processes|10261,10270
,|10270,10271
such|10272,10276
as|10277,10279
an|10280,10282
infection|10283,10292
.|10292,10293
<EOL>|10294,10295
While|10295,10300
you|10301,10304
were|10305,10309
in|10310,10312
the|10313,10316
hospital|10317,10325
,|10325,10326
you|10327,10330
were|10331,10335
seen|10336,10340
by|10341,10343
one|10344,10347
of|10348,10350
our|10351,10354
<EOL>|10355,10356
social|10356,10362
workers|10363,10370
.|10370,10371
You|10372,10375
will|10376,10380
also|10381,10385
follow|10386,10392
up|10393,10395
with|10396,10400
Palliative|10401,10411
Care|10412,10416
in|10417,10419
<EOL>|10420,10421
their|10421,10426
clinic|10427,10433
and|10434,10437
will|10438,10442
continue|10443,10451
to|10452,10454
have|10455,10459
therapeutic|10460,10471
paracenteses|10472,10484
.|10484,10485
<EOL>|10485,10486
<EOL>|10486,10487
It|10487,10489
has|10490,10493
been|10494,10498
a|10499,10500
pleasure|10501,10509
taking|10510,10516
care|10517,10521
of|10522,10524
you|10525,10528
and|10529,10532
we|10533,10535
wish|10536,10540
you|10541,10544
all|10545,10548
<EOL>|10549,10550
the|10550,10553
best|10554,10558
,|10558,10559
<EOL>|10559,10560
Your|10560,10564
_|10565,10566
_|10566,10567
_|10567,10568
Care|10569,10573
team|10574,10578
<EOL>|10578,10579
<EOL>|10580,10581
Followup|10581,10589
Instructions|10590,10602
:|10602,10603
<EOL>|10603,10604
_|10604,10605
_|10605,10606
_|10606,10607
<EOL>|10607,10608

