 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|47,56|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|47,56|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|47,61|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|81,90|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|81,90|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|81,90|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|81,90|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|81,90|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|81,95|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|113,118|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|113,118|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|113,118|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|137,140|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|137,140|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|137,140|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|137,140|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|137,140|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|148,155|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|148,155|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|SIMPLE_SEGMENT|157,164|false|false|false|||SURGERY
Finding|Finding|SIMPLE_SEGMENT|157,164|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Finding|Functional Concept|SIMPLE_SEGMENT|157,164|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Finding|Idea or Concept|SIMPLE_SEGMENT|157,164|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|157,164|false|false|false|C0543467|Operative Surgical Procedures|SURGERY
Attribute|Clinical Attribute|Allergies|188,197|false|false|false|C1717415||Allergies
Event|Event|Allergies|188,197|false|false|false|||Allergies
Finding|Pathologic Function|Allergies|188,197|false|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|Allergies|200,222|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|Allergies|208,212|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|Allergies|208,212|false|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|Allergies|208,222|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Event|Event|Allergies|213,222|false|false|false|||Reactions
Event|Event|Allergies|225,234|false|false|false|||Attending
Finding|Functional Concept|Allergies|225,234|false|false|false|C1999232|Attending (action)|Attending
Disorder|Neoplastic Process|Chief Complaint|260,294|false|false|false|C5206813|Locally Advanced Gastric Carcinoma|Locally advanced gastric carcinoma
Anatomy|Body Part, Organ, or Organ Component|Chief Complaint|277,284|false|false|false|C0038351|Stomach|gastric
Disorder|Neoplastic Process|Chief Complaint|277,294|false|false|false|C0699791|Stomach Carcinoma|gastric carcinoma
Disorder|Neoplastic Process|Chief Complaint|285,294|false|false|false|C0007097|Carcinoma|carcinoma
Event|Event|Chief Complaint|285,294|false|false|false|||carcinoma
Finding|Classification|Chief Complaint|297,302|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|303,311|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|303,311|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|315,333|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|324,333|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|324,333|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|324,333|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|324,333|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|324,333|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|Chief Complaint|335,345|false|false|false|||Cystoscopy
Procedure|Diagnostic Procedure|Chief Complaint|335,345|false|false|false|C0010702|Cystoscopy|Cystoscopy
Event|Event|Chief Complaint|356,364|false|false|false|||catheter
Finding|Intellectual Product|Chief Complaint|356,364|false|true|false|C1546572||catheter
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|356,374|false|true|false|C0883301|Catheter placement|catheter placement
Event|Event|Chief Complaint|365,374|false|false|false|||placement
Procedure|Health Care Activity|Chief Complaint|365,374|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|365,374|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Event|Event|Chief Complaint|376,387|false|false|false|||Laparoscopy
Procedure|Diagnostic Procedure|Chief Complaint|376,387|false|false|false|C0031150;C1883297|Laparoscopy;Therapeutic Laparoscopy|Laparoscopy
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|376,387|false|false|false|C0031150;C1883297|Laparoscopy;Therapeutic Laparoscopy|Laparoscopy
Event|Event|Chief Complaint|394,400|false|false|false|||biopsy
Finding|Finding|Chief Complaint|394,400|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Finding|Intellectual Product|Chief Complaint|394,400|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Procedure|Diagnostic Procedure|Chief Complaint|394,400|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Procedure|Health Care Activity|Chief Complaint|394,400|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Event|Event|Chief Complaint|402,413|false|false|false|||Gastroscopy
Procedure|Diagnostic Procedure|Chief Complaint|402,413|false|false|false|C0017195|Endoscopy of stomach|Gastroscopy
Finding|Idea or Concept|History of Present Illness|462,466|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|History of Present Illness|462,466|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|History of Present Illness|467,470|false|false|false|||old
Finding|Finding|History of Present Illness|471,475|false|false|false|C1706180|Male Gender|male
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|498,505|false|false|false|C0038351|Stomach|gastric
Disorder|Neoplastic Process|History of Present Illness|507,513|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|History of Present Illness|507,513|false|false|false|||cancer
Attribute|Clinical Attribute|History of Present Illness|515,520|false|false|false|C1300072|Tumor stage|stage
Event|Event|History of Present Illness|536,543|false|false|false|||arrives
Event|Event|History of Present Illness|556,564|false|false|false|||curative
Finding|Conceptual Entity|History of Present Illness|556,564|false|false|false|C1880198|Cure (remedy)|curative
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|556,564|false|false|false|C1276305|Curative - procedure intent|curative
Finding|Idea or Concept|History of Present Illness|565,571|false|false|false|C0162425;C1550453|Act Mood - intent|intent
Finding|Mental Process|History of Present Illness|565,571|false|false|false|C0162425;C1550453|Act Mood - intent|intent
Procedure|Health Care Activity|History of Present Illness|572,580|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|572,580|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|572,590|false|false|false|C0015252;C0728940|Excision;removal technique|surgical resection
Event|Event|History of Present Illness|581,590|false|false|false|||resection
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|581,590|false|false|false|C0015252;C0728940|Excision;removal technique|resection
Event|Event|History of Present Illness|597,607|false|false|false|||completion
Event|Event|History of Present Illness|611,620|false|false|false|||induction
Finding|Functional Concept|History of Present Illness|611,620|false|false|false|C0205263|Induce (action)|induction
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|611,620|false|false|false|C0857127|Induction procedure|induction
Event|Event|History of Present Illness|622,634|false|false|false|||chemotherapy
Finding|Functional Concept|History of Present Illness|622,634|false|false|false|C0013217|pharmacotherapeutic|chemotherapy
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|622,634|false|false|false|C0013216;C0392920;C3665472|Chemotherapy;Chemotherapy Regimen;Pharmacotherapy|chemotherapy
Event|Event|History of Present Illness|645,652|false|false|false|||started
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|656,667|false|false|false|C0600558|Neoadjuvant Therapy|neoadjuvant
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|656,680|false|false|false|C5392214|Neoadjuvant Chemotherapy|neoadjuvant chemotherapy
Event|Event|History of Present Illness|668,680|false|false|false|||chemotherapy
Finding|Functional Concept|History of Present Illness|668,680|false|false|false|C0013217|pharmacotherapeutic|chemotherapy
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|668,680|false|false|false|C0013216;C0392920;C3665472|Chemotherapy;Chemotherapy Regimen;Pharmacotherapy|chemotherapy
Finding|Intellectual Product|History of Present Illness|700,707|false|false|false|C0282416|Overall Publication Type|Overall
Event|Event|History of Present Illness|711,720|false|false|false|||tolerated
Event|Event|History of Present Illness|725,737|false|false|false|||chemotherapy
Finding|Functional Concept|History of Present Illness|725,737|false|false|false|C0013217|pharmacotherapeutic|chemotherapy
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|725,737|false|false|false|C0013216;C0392920;C3665472|Chemotherapy;Chemotherapy Regimen;Pharmacotherapy|chemotherapy
Finding|Finding|History of Present Illness|738,742|false|false|false|C5575035|Well (answer to question)|well
Finding|Idea or Concept|History of Present Illness|756,767|false|false|false|C0750502|Significant|significant
Finding|Functional Concept|History of Present Illness|768,780|false|false|false|C0001688;C0879626|Adverse effects;aspects of adverse effects|side effects
Finding|Pathologic Function|History of Present Illness|768,780|false|false|false|C0001688;C0879626|Adverse effects;aspects of adverse effects|side effects
Event|Event|History of Present Illness|773,780|false|false|false|||effects
Finding|Idea or Concept|History of Present Illness|796,801|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|History of Present Illness|796,801|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Event|Event|History of Present Illness|805,814|false|false|false|||developed
Finding|Functional Concept|History of Present Illness|815,820|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|815,836|false|false|false|C0230329|Right upper extremity|right upper extremity
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|821,836|false|false|false|C1140618|Upper Extremity|upper extremity
Finding|Pathologic Function|History of Present Illness|821,842|false|false|false|C0522035|Edema of the upper extremity|upper extremity edema
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|827,836|false|false|false|C0015385|Limb structure|extremity
Finding|Pathologic Function|History of Present Illness|827,842|false|false|false|C0085649|Peripheral edema|extremity edema
Attribute|Clinical Attribute|History of Present Illness|837,842|false|false|false|C1717255||edema
Event|Event|History of Present Illness|837,842|false|false|false|||edema
Finding|Pathologic Function|History of Present Illness|837,842|false|false|false|C0013604|Edema|edema
Event|Event|History of Present Illness|851,856|false|false|false|||noted
Event|Event|History of Present Illness|867,877|false|false|false|||thrombosis
Finding|Pathologic Function|History of Present Illness|867,877|false|false|false|C0040053|Thrombosis|thrombosis
Event|Event|History of Present Illness|899,906|false|false|false|||started
Drug|Organic Chemical|History of Present Illness|910,917|false|false|false|C0728963|Lovenox|Lovenox
Drug|Pharmacologic Substance|History of Present Illness|910,917|false|false|false|C0728963|Lovenox|Lovenox
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|927,930|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|927,930|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|History of Present Illness|927,930|false|false|false|C1530795|BID protein, human|BID
Event|Event|History of Present Illness|927,930|false|false|false|||BID
Finding|Gene or Genome|History of Present Illness|927,930|false|false|false|C1332410|BID gene|BID
Event|Event|History of Present Illness|944,953|false|false|false|||compliant
Finding|Individual Behavior|History of Present Illness|944,953|false|false|false|C1321605|Compliance behavior|compliant
Event|Event|History of Present Illness|960,966|false|false|false|||Denies
Event|Event|History of Present Illness|971,976|false|false|false|||fever
Finding|Finding|History of Present Illness|971,976|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|History of Present Illness|971,976|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Attribute|Clinical Attribute|History of Present Illness|978,984|true|false|false|C4255480||nausea
Event|Event|History of Present Illness|978,984|false|false|false|||nausea
Finding|Sign or Symptom|History of Present Illness|978,984|true|false|false|C0027497|Nausea|nausea
Event|Event|History of Present Illness|986,992|false|false|false|||emesis
Finding|Body Substance|History of Present Illness|986,992|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Physiologic Function|History of Present Illness|986,992|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Sign or Symptom|History of Present Illness|986,992|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Event|Event|History of Present Illness|994,1000|false|false|false|||chills
Finding|Sign or Symptom|History of Present Illness|994,1000|false|false|false|C0085593|Chills|chills
Attribute|Clinical Attribute|History of Present Illness|1002,1008|false|false|false|C0944911||weight
Event|Event|History of Present Illness|1002,1008|false|false|false|||weight
Finding|Finding|History of Present Illness|1002,1008|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|History of Present Illness|1002,1008|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|History of Present Illness|1002,1008|false|false|false|C1305866|Weighing patient|weight
Finding|Finding|History of Present Illness|1002,1013|false|false|false|C1262477;C3540682|Losing Weight (question);Weight Loss|weight loss
Finding|Intellectual Product|History of Present Illness|1002,1013|false|false|false|C1262477;C3540682|Losing Weight (question);Weight Loss|weight loss
Event|Event|History of Present Illness|1009,1013|false|false|false|||loss
Finding|Finding|History of Present Illness|1009,1013|false|false|false|C5890125|Loss (adaptation)|loss
Event|Event|History of Present Illness|1015,1021|false|false|false|||melena
Finding|Pathologic Function|History of Present Illness|1015,1021|false|false|false|C0025222|Melena|melena
Disorder|Disease or Syndrome|History of Present Illness|1023,1035|false|false|false|C0018932|Hematochezia|hematochezia
Event|Event|History of Present Illness|1023,1035|false|false|false|||hematochezia
Finding|Sign or Symptom|History of Present Illness|1023,1035|false|false|false|C1321898|Blood in stool|hematochezia
Disorder|Disease or Syndrome|History of Present Illness|1039,1048|false|false|false|C0018965|Hematuria|hematuria
Event|Event|History of Present Illness|1039,1048|false|false|false|||hematuria
Event|Event|History of Present Illness|1055,1060|false|false|false|||comes
Finding|Functional Concept|History of Present Illness|1074,1080|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Event|Event|History of Present Illness|1081,1088|false|false|false|||staging
Finding|Functional Concept|History of Present Illness|1081,1088|false|false|false|C0332305|With staging|staging
Event|Event|History of Present Illness|1106,1108|false|false|false|||CT
Event|Event|History of Present Illness|1109,1113|false|false|false|||scan
Procedure|Diagnostic Procedure|History of Present Illness|1109,1113|false|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Event|Event|History of Present Illness|1114,1127|false|false|false|||demonstrating
Event|Event|History of Present Illness|1131,1139|false|false|false|||evidence
Finding|Idea or Concept|History of Present Illness|1131,1139|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|History of Present Illness|1131,1142|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Disease or Syndrome|History of Present Illness|1143,1150|true|false|false|C0012634|Disease|disease
Event|Event|History of Present Illness|1143,1150|false|false|false|||disease
Event|Event|History of Present Illness|1166,1171|false|false|false|||taken
Finding|Finding|History of Present Illness|1179,1188|false|false|false|C4738506|Operating|operating
Finding|Finding|History of Present Illness|1221,1229|false|false|false|C0332149|Possible|possibly
Drug|Chemical Viewed Structurally|History of Present Illness|1235,1242|false|false|false|C0302912|Radicals (chemistry)|radical
Event|Event|History of Present Illness|1235,1242|false|false|false|||radical
Attribute|Clinical Attribute|History of Present Illness|1243,1249|false|false|false|C4522154|Distal Resection Margin|distal
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1243,1261|false|false|false|C0176758;C0192440|Billroth I Procedure;Partial gastrectomy with anastomosis to duodenum|distal gastrectomy
Event|Event|History of Present Illness|1250,1261|false|false|false|||gastrectomy
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1250,1261|false|false|false|C0017118|Gastrectomy|gastrectomy
Event|Event|History of Present Illness|1267,1282|false|false|false|||lymphadenectomy
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1267,1282|false|false|false|C0024203|Lymph node excision|lymphadenectomy
Event|Event|History of Present Illness|1289,1294|false|false|false|||risks
Finding|Idea or Concept|History of Present Illness|1289,1294|false|false|false|C0035647|Risk|risks
Event|Event|History of Present Illness|1299,1307|false|false|false|||benefits
Event|Event|History of Present Illness|1311,1318|false|false|false|||surgery
Finding|Finding|History of Present Illness|1311,1318|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|History of Present Illness|1311,1318|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|History of Present Illness|1311,1318|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1311,1318|false|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Event|History of Present Illness|1329,1338|false|false|false|||described
Finding|Body Substance|History of Present Illness|1348,1355|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1348,1355|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1348,1355|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|History of Present Illness|1359,1365|false|false|false|C1561567|detail - Response Level|detail
Event|Event|History of Present Illness|1374,1384|false|false|false|||documented
Event|Event|History of Present Illness|1410,1414|false|false|false|||note
Finding|Finding|Past Medical History|1440,1460|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|Past Medical History|1445,1452|false|false|false|||Medical
Finding|Functional Concept|Past Medical History|1445,1452|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|Past Medical History|1445,1452|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|Past Medical History|1445,1452|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|Past Medical History|1445,1452|false|false|false|C0199168|Medical service|Medical
Finding|Finding|Past Medical History|1445,1460|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|Past Medical History|1453,1460|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|Past Medical History|1453,1460|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|Past Medical History|1453,1460|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1462,1470|false|false|false|C0033572;C4266527|Prostate;Structure of prostate (body structure)|Prostate
Disorder|Disease or Syndrome|Past Medical History|1462,1470|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|Prostate
Disorder|Neoplastic Process|Past Medical History|1462,1470|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|Prostate
Disorder|Neoplastic Process|Past Medical History|1462,1477|false|false|false|C0376358;C0600139|Malignant neoplasm of prostate;Prostate carcinoma|Prostate cancer
Disorder|Neoplastic Process|Past Medical History|1471,1477|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Past Medical History|1471,1477|false|false|false|||cancer
Disorder|Neoplastic Process|Past Medical History|1471,1486|false|false|false|C0549473|Thyroid carcinoma|cancer, Thyroid
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1479,1486|false|false|false|C0040132|Thyroid Gland|Thyroid
Disorder|Disease or Syndrome|Past Medical History|1479,1486|false|false|false|C0040128|Thyroid Diseases|Thyroid
Drug|Amino Acid, Peptide, or Protein|Past Medical History|1479,1486|false|false|false|C0040134;C3540038;C5781115|THYROID;THYROID DIAGNOSTIC RADIOPHARMACEUTICALS;thyroid (USP)|Thyroid
Drug|Hormone|Past Medical History|1479,1486|false|false|false|C0040134;C3540038;C5781115|THYROID;THYROID DIAGNOSTIC RADIOPHARMACEUTICALS;thyroid (USP)|Thyroid
Drug|Indicator, Reagent, or Diagnostic Aid|Past Medical History|1479,1486|false|false|false|C0040134;C3540038;C5781115|THYROID;THYROID DIAGNOSTIC RADIOPHARMACEUTICALS;thyroid (USP)|Thyroid
Drug|Organic Chemical|Past Medical History|1479,1486|false|false|false|C0040134;C3540038;C5781115|THYROID;THYROID DIAGNOSTIC RADIOPHARMACEUTICALS;thyroid (USP)|Thyroid
Drug|Pharmacologic Substance|Past Medical History|1479,1486|false|false|false|C0040134;C3540038;C5781115|THYROID;THYROID DIAGNOSTIC RADIOPHARMACEUTICALS;thyroid (USP)|Thyroid
Event|Event|Past Medical History|1479,1486|false|false|false|||Thyroid
Procedure|Health Care Activity|Past Medical History|1479,1486|false|false|false|C2228489|examination of thyroid|Thyroid
Disorder|Neoplastic Process|Past Medical History|1479,1493|false|false|false|C0040137|Thyroid Nodule|Thyroid nodule
Finding|Finding|Past Medical History|1479,1493|false|false|false|C2116082||Thyroid nodule
Event|Event|Past Medical History|1487,1493|false|false|false|||nodule
Disorder|Disease or Syndrome|Past Medical History|1495,1506|false|false|false|C0020676|Hypothyroidism|Hypothyroid
Event|Event|Past Medical History|1495,1506|false|false|false|||Hypothyroid
Disorder|Disease or Syndrome|Past Medical History|1508,1512|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|Past Medical History|1508,1512|false|false|false|||GERD
Finding|Intellectual Product|Past Medical History|1513,1517|false|false|false|C1547225|Mild Severity of Illness Code|mild
Disorder|Disease or Syndrome|Past Medical History|1519,1533|false|false|false|C1510475|Diverticulosis|Diverticulosis
Event|Event|Past Medical History|1519,1533|false|false|false|||Diverticulosis
Event|Event|Past Medical History|1537,1548|false|false|false|||colonoscopy
Procedure|Diagnostic Procedure|Past Medical History|1537,1548|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Procedure|Health Care Activity|Past Medical History|1537,1548|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Disorder|Disease or Syndrome|Past Medical History|1553,1559|false|false|false|C0002871|Anemia|anemia
Event|Event|Past Medical History|1553,1559|false|false|false|||anemia
Drug|Biologically Active Substance|Past Medical History|1560,1564|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|Past Medical History|1560,1564|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|Past Medical History|1560,1564|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Event|Event|Past Medical History|1560,1564|false|false|false|||iron
Procedure|Laboratory Procedure|Past Medical History|1560,1564|false|false|false|C0337439|Iron measurement|iron
Drug|Hazardous or Poisonous Substance|Past Medical History|1565,1568|false|false|false|C0054282|butyl phosphorotrithioate|def
Drug|Organic Chemical|Past Medical History|1565,1568|false|false|false|C0054282|butyl phosphorotrithioate|def
Event|Event|Past Medical History|1565,1568|false|false|false|||def
Finding|Gene or Genome|Past Medical History|1565,1568|false|false|false|C1823727|UTP25 gene|def
Disorder|Disease or Syndrome|Past Medical History|1570,1576|false|false|false|C0002871|Anemia|anemia
Event|Event|Past Medical History|1570,1576|false|false|false|||anemia
Event|Event|Past Medical History|1583,1591|false|false|false|||resolved
Event|Event|Past Medical History|1599,1605|false|false|false|||workup
Finding|Finding|Past Medical History|1607,1628|false|false|false|C0455610|History of surgery|Past Surgical History
Procedure|Health Care Activity|Past Medical History|1612,1620|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1612,1620|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Finding|Finding|Past Medical History|1612,1628|false|false|false|C0744961|history of prior surgery|Surgical History
Event|Event|Past Medical History|1621,1628|false|false|false|||History
Finding|Conceptual Entity|Past Medical History|1621,1628|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|Past Medical History|1621,1628|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|Past Medical History|1621,1628|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1630,1638|false|false|false|C0033572;C4266527|Prostate;Structure of prostate (body structure)|Prostate
Disorder|Disease or Syndrome|Past Medical History|1630,1638|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|Prostate
Disorder|Neoplastic Process|Past Medical History|1630,1638|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|Prostate
Disorder|Neoplastic Process|Past Medical History|1630,1645|false|false|false|C0376358;C0600139|Malignant neoplasm of prostate;Prostate carcinoma|Prostate cancer
Disorder|Neoplastic Process|Past Medical History|1639,1645|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Past Medical History|1639,1645|false|false|false|||cancer
Anatomy|Body Location or Region|Past Medical History|1646,1654|false|false|false|C1548801|Body Site Modifier - External|external
Finding|Functional Concept|Past Medical History|1646,1654|false|false|false|C0521134|External route|external
Drug|Organic Chemical|Past Medical History|1655,1659|false|false|false|C4521565|Beam -- chemical|beam
Drug|Pharmacologic Substance|Past Medical History|1655,1659|false|false|false|C4521565|Beam -- chemical|beam
Event|Event|Past Medical History|1655,1659|false|false|false|||beam
Phenomenon|Phenomenon or Process|Past Medical History|1655,1659|false|false|false|C2347880|Beam - rays of radiation or stream of particles|beam
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1655,1659|false|false|false|C0338248|carmustine/cytarabine/etoposide/melphalan regimen|beam
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1665,1673|false|false|false|C0001074|Structure of achilles tendon|Achilles
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1665,1680|false|false|false|C0001074;C1305378|Structure of achilles tendon|Achilles tendon
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1665,1687|false|false|false|C0407029|Repair of Achilles tendon|Achilles tendon repair
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1674,1680|false|false|false|C0039508|Tendon structure|tendon
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1674,1687|false|false|false|C0565350|Plastic repair of tendon|tendon repair
Event|Event|Past Medical History|1681,1687|false|false|false|||repair
Finding|Functional Concept|Past Medical History|1681,1687|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Finding|Organism Function|Past Medical History|1681,1687|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Procedure|Health Care Activity|Past Medical History|1681,1687|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1681,1687|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Finding|Functional Concept|Past Medical History|1703,1708|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1703,1714|false|false|false|C0817321|Right tibia|right tibia
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1709,1714|false|false|false|C0040184|Bone structure of tibia|tibia
Anatomy|Body Location or Region|Past Medical History|1709,1725|false|false|false|C0947635|tibia and fibula|tibia and fibula
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1719,1725|false|false|false|C0016068|Fibula|fibula
Event|Event|Past Medical History|1727,1740|false|false|false|||Tonsillectomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1727,1740|false|false|false|C0040423|Tonsillectomy|Tonsillectomy
Attribute|Clinical Attribute|Past Medical History|1741,1744|false|false|false|C1114365||age
Drug|Biologically Active Substance|Past Medical History|1741,1744|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|Past Medical History|1741,1744|false|false|false|C0162574|Glycation End Products, Advanced|age
Event|Event|Past Medical History|1741,1744|false|false|false|||age
Finding|Conceptual Entity|Family Medical History|1788,1794|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|Family Medical History|1788,1794|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Event|Event|Family Medical History|1795,1799|false|false|false|||died
Disorder|Neoplastic Process|Family Medical History|1812,1820|false|false|false|C0024299|Lymphoma|Lymphoma
Event|Event|Family Medical History|1812,1820|false|false|false|||Lymphoma
Finding|Idea or Concept|Family Medical History|1822,1828|false|false|false|C1546508|Relationship - Mother|Mother
Event|Event|Family Medical History|1829,1833|false|false|false|||died
Finding|Gene or Genome|Family Medical History|1846,1850|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Intellectual Product|Family Medical History|1846,1850|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Disorder|Mental or Behavioral Dysfunction|Family Medical History|1859,1867|false|false|false|C0011265;C0497327|Dementia;Presenile dementia|Dementia
Event|Event|Family Medical History|1859,1867|false|false|false|||Dementia
Event|Event|General Exam|1898,1902|false|false|false|||Data
Finding|Idea or Concept|General Exam|1898,1902|false|false|false|C1511726|Data|Data
Event|Event|General Exam|1909,1916|false|false|false|||updated
Event|Event|General Exam|1933,1937|false|false|false|||Temp
Finding|Gene or Genome|General Exam|1933,1937|false|false|false|C1823816|C1orf210 gene|Temp
Procedure|Therapeutic or Preventive Procedure|General Exam|1933,1937|false|false|false|C0279848|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Temp
Event|Event|General Exam|1983,1985|false|false|false|||HR
Event|Event|General Exam|2038,2046|false|false|false|||delivery
Finding|Finding|General Exam|2038,2046|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Finding|Functional Concept|General Exam|2038,2046|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Finding|Organism Function|General Exam|2038,2046|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Procedure|Therapeutic or Preventive Procedure|General Exam|2038,2046|false|false|false|C0011209|Obstetric Delivery|delivery
Event|Event|General Exam|2053,2056|false|false|false|||GEN
Finding|Classification|General Exam|2053,2056|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|GEN
Finding|Gene or Genome|General Exam|2053,2056|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|GEN
Event|Event|General Exam|2060,2063|false|false|false|||Ox3
Disorder|Disease or Syndrome|General Exam|2065,2068|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|2065,2068|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|2065,2068|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|2065,2068|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|2065,2068|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|General Exam|2065,2068|false|false|false|||NAD
Finding|Finding|General Exam|2065,2068|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Event|Event|General Exam|2070,2077|false|false|false|||resting
Anatomy|Body Location or Region|General Exam|2091,2096|false|false|false|C1512338|HEENT|HEENT
Event|Event|General Exam|2098,2102|false|false|false|||NCAT
Event|Event|General Exam|2104,2108|false|false|false|||EOMI
Anatomy|Body Part, Organ, or Organ Component|General Exam|2110,2116|false|false|false|C0036410|Sclera|sclera
Disorder|Disease or Syndrome|General Exam|2110,2116|false|false|false|C0036412|Scleral Diseases|sclera
Event|Event|General Exam|2110,2116|false|false|false|||sclera
Procedure|Health Care Activity|General Exam|2110,2116|false|false|false|C2228481|examination of sclera|sclera
Event|Event|General Exam|2117,2126|false|false|false|||anicteric
Finding|Finding|General Exam|2117,2126|false|false|false|C0205180|Anicteric|anicteric
Event|Event|General Exam|2131,2134|false|false|false|||RRR
Event|Event|General Exam|2135,2139|false|false|false|||PULM
Procedure|Health Care Activity|General Exam|2135,2139|false|false|false|C1315068|Pulmonary ventilator management|PULM
Attribute|Clinical Attribute|General Exam|2144,2155|true|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|General Exam|2144,2155|true|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|General Exam|2144,2155|true|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|General Exam|2144,2155|true|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Sign or Symptom|General Exam|2144,2164|true|false|false|C0476273|Respiratory distress|respiratory distress
Event|Event|General Exam|2156,2164|false|false|false|||distress
Finding|Finding|General Exam|2156,2164|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|General Exam|2156,2164|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|General Exam|2165,2168|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|ABD
Disorder|Cell or Molecular Dysfunction|General Exam|2165,2168|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|ABD
Event|Event|General Exam|2165,2168|false|false|false|||ABD
Disorder|Disease or Syndrome|General Exam|2170,2174|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|General Exam|2170,2174|false|false|false|||soft
Event|Event|General Exam|2187,2194|false|false|false|||rebound
Event|Event|General Exam|2198,2206|false|false|false|||guarding
Finding|Finding|General Exam|2198,2206|true|false|false|C0427198|Protective muscle spasm|guarding
Disorder|Congenital Abnormality|General Exam|2208,2211|false|false|false|C0015306|Hereditary Multiple Exostoses|EXT
Event|Event|General Exam|2208,2211|false|false|false|||EXT
Finding|Gene or Genome|General Exam|2208,2211|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|EXT
Event|Event|General Exam|2213,2217|false|false|false|||warm
Finding|Finding|General Exam|2213,2217|false|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|General Exam|2213,2217|false|false|false|C0687712|warming process|warm
Finding|Finding|General Exam|2219,2223|false|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|2224,2232|false|false|false|||perfused
Attribute|Clinical Attribute|General Exam|2237,2242|true|false|false|C1717255||edema
Event|Event|General Exam|2237,2242|false|false|false|||edema
Finding|Pathologic Function|General Exam|2237,2242|true|false|false|C0013604|Edema|edema
Disorder|Mental or Behavioral Dysfunction|General Exam|2244,2249|false|false|false|C0004936;C1306597|Mental disorders;Psychiatric problem|PSYCH
Event|Event|General Exam|2244,2249|false|false|false|||PSYCH
Event|Event|General Exam|2258,2265|false|false|false|||insight
Finding|Mental Process|General Exam|2258,2265|false|false|false|C0233820|Insight|insight
Event|Event|General Exam|2267,2273|false|false|false|||memory
Finding|Finding|General Exam|2267,2273|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Intellectual Product|General Exam|2267,2273|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Mental Process|General Exam|2267,2273|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Attribute|Clinical Attribute|General Exam|2279,2283|false|false|false|C2713234||mood
Event|Event|General Exam|2279,2283|false|false|false|||mood
Finding|Conceptual Entity|General Exam|2279,2283|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|mood
Finding|Finding|General Exam|2279,2283|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|mood
Finding|Mental Process|General Exam|2279,2283|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|mood
Disorder|Injury or Poisoning|General Exam|2284,2289|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|WOUND
Event|Event|General Exam|2284,2289|false|false|false|||WOUND
Finding|Body Substance|General Exam|2284,2289|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|WOUND
Finding|Functional Concept|General Exam|2284,2289|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|WOUND
Finding|Intellectual Product|General Exam|2284,2289|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|WOUND
Anatomy|Body Location or Region|General Exam|2294,2302|false|false|false|C2338258|Cranial incision point|Incision
Disorder|Injury or Poisoning|General Exam|2294,2302|false|false|false|C0332803|Surgical wound|Incision
Procedure|Therapeutic or Preventive Procedure|General Exam|2294,2302|false|false|false|C0184898|Surgical incisions|Incision
Finding|Idea or Concept|Hospital Course|2351,2355|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|Hospital Course|2351,2355|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|Hospital Course|2360,2364|false|false|false|||Male
Finding|Finding|Hospital Course|2360,2364|false|false|false|C1706180|Male Gender|Male
Event|Event|Hospital Course|2369,2378|false|false|false|||presented
Event|Event|Hospital Course|2393,2400|false|false|false|||planned
Finding|Finding|Hospital Course|2424,2432|false|false|false|C0332149|Possible|possibly
Drug|Chemical Viewed Structurally|Hospital Course|2438,2445|false|false|false|C0302912|Radicals (chemistry)|radical
Attribute|Clinical Attribute|Hospital Course|2446,2452|false|false|false|C4522154|Distal Resection Margin|distal
Event|Event|Hospital Course|2454,2465|false|false|false|||gastrectomy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2454,2465|false|false|false|C0017118|Gastrectomy|gastrectomy
Event|Event|Hospital Course|2471,2486|false|false|false|||lymphadenectomy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2471,2486|false|false|false|C0024203|Lymph node excision|lymphadenectomy
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|2508,2515|false|false|false|C0038351|Stomach|gastric
Disorder|Neoplastic Process|Hospital Course|2517,2526|false|false|false|C0007097|Carcinoma|carcinoma
Event|Event|Hospital Course|2517,2526|false|false|false|||carcinoma
Event|Event|Hospital Course|2533,2545|false|false|false|||chemotherapy
Finding|Functional Concept|Hospital Course|2533,2545|false|false|false|C0013217|pharmacotherapeutic|chemotherapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2533,2545|false|false|false|C0013216;C0392920;C3665472|Chemotherapy;Chemotherapy Regimen;Pharmacotherapy|chemotherapy
Event|Event|Hospital Course|2553,2562|false|false|false|||placement
Procedure|Health Care Activity|Hospital Course|2553,2562|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2553,2562|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Finding|Functional Concept|Hospital Course|2570,2575|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Drug|Food|Hospital Course|2592,2596|false|false|false|C0452253|Port - alcoholic beverage|port
Event|Event|Hospital Course|2592,2596|false|false|false|||port
Event|Event|Hospital Course|2598,2610|false|false|false|||insufflation
Finding|Functional Concept|Hospital Course|2598,2610|false|false|false|C4281791|Insufflation route|insufflation
Procedure|Health Care Activity|Hospital Course|2598,2610|false|false|false|C0021634|Insufflation|insufflation
Event|Event|Hospital Course|2611,2619|false|false|false|||revealed
Finding|Functional Concept|Hospital Course|2624,2629|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|Hospital Course|2624,2644|false|false|false|C0230177|Structure of right upper quadrant of abdomen|right upper quadrant
Drug|Food|Hospital Course|2646,2650|false|false|false|C0452253|Port - alcoholic beverage|port
Event|Event|Hospital Course|2646,2650|false|false|false|||port
Event|Event|Hospital Course|2657,2668|false|false|false|||penetrating
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|2673,2680|false|false|false|C0028977|Omentum|omentum
Event|Event|Hospital Course|2685,2693|false|false|false|||appeared
Event|Event|Hospital Course|2697,2701|false|false|false|||miss
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|2707,2727|false|false|false|C0230254|Structure of transverse mesocolon|transverse mesocolon
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|2718,2727|false|false|false|C0025483|Mesocolon|mesocolon
Finding|Finding|Hospital Course|2731,2735|false|false|false|C5575035|Well (answer to question)|well
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|2743,2748|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|Hospital Course|2743,2748|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|Hospital Course|2743,2748|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Finding|Finding|Hospital Course|2743,2748|false|false|false|C0750873|COLON PROBLEM|colon
Event|Event|Hospital Course|2749,2755|false|false|false|||itself
Event|Event|Hospital Course|2769,2776|false|false|false|||surgery
Finding|Finding|Hospital Course|2769,2776|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Hospital Course|2769,2776|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Hospital Course|2769,2776|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2769,2776|false|false|false|C0543467|Operative Surgical Procedures|surgery
Anatomy|Body Location or Region|Hospital Course|2806,2816|false|false|false|C0031153;C0442034|Peritoneum;peritoneal|peritoneal
Anatomy|Tissue|Hospital Course|2806,2816|false|false|false|C0031153;C0442034|Peritoneum;peritoneal|peritoneal
Event|Event|Hospital Course|2817,2825|false|false|false|||deposits
Finding|Functional Concept|Hospital Course|2817,2825|false|false|false|C0333562|Deposition (morphologic abnormality)|deposits
Anatomy|Body Location or Region|Hospital Course|2834,2844|false|false|false|C0031153;C0442034|Peritoneum;peritoneal|peritoneal
Anatomy|Tissue|Hospital Course|2834,2844|false|false|false|C0031153;C0442034|Peritoneum;peritoneal|peritoneal
Event|Event|Hospital Course|2845,2853|false|false|false|||surfaces
Event|Event|Hospital Course|2883,2895|false|false|false|||demonstrated
Disorder|Neoplastic Process|Hospital Course|2908,2922|false|false|false|C0205699;C2007060|Carcinomatosis;carcinomatosis of unspecified behavior|carcinomatosis
Event|Event|Hospital Course|2908,2922|false|false|false|||carcinomatosis
Disorder|Neoplastic Process|Hospital Course|2947,2961|false|false|false|C0001418;C5551397|Adenocarcinoma;Malignant adenomatous neoplasm|adenocarcinoma
Event|Event|Hospital Course|2947,2961|false|false|false|||adenocarcinoma
Event|Event|Hospital Course|2963,2972|false|false|false|||involving
Anatomy|Tissue|Hospital Course|2977,2987|false|false|false|C0031153;C0230198;C4482223|Abdomen>Peritoneum;Peritoneum;Serous layer of peritoneum|peritoneum
Disorder|Neoplastic Process|Hospital Course|2977,2987|false|false|false|C0496874;C0496954|Benign neoplasm of peritoneum;Neoplasm of uncertain or unknown behavior of peritoneum|peritoneum
Event|Event|Hospital Course|2998,3004|false|false|false|||reason
Finding|Idea or Concept|Hospital Course|2998,3004|false|false|false|C0392360|Indication of (contextual qualifier)|reason
Attribute|Clinical Attribute|Hospital Course|3010,3019|false|false|false|C0945766||procedure
Event|Event|Hospital Course|3010,3019|false|false|false|||procedure
Event|Occupational Activity|Hospital Course|3010,3019|false|false|false|C1546467|Act Class - procedure|procedure
Finding|Functional Concept|Hospital Course|3010,3019|false|false|false|C2700391|Procedure (set of actions)|procedure
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3010,3019|false|false|false|C0184661|Interventional procedure|procedure
Finding|Intellectual Product|Hospital Course|3025,3029|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|Hospital Course|3030,3037|false|false|false|||aborted
Finding|Body Substance|Hospital Course|3060,3067|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|3060,3067|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|3060,3067|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|3072,3077|false|false|false|||taken
Event|Event|Hospital Course|3085,3089|false|false|false|||PACU
Event|Event|Hospital Course|3097,3103|false|false|false|||stable
Finding|Intellectual Product|Hospital Course|3097,3103|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Intellectual Product|Hospital Course|3108,3112|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|Hospital Course|3113,3124|false|false|false|||transferred
Event|Event|Hospital Course|3144,3150|false|false|false|||stable
Finding|Intellectual Product|Hospital Course|3144,3150|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|Hospital Course|3158,3162|false|false|false|||home
Finding|Idea or Concept|Hospital Course|3158,3162|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|3158,3162|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|3158,3162|false|false|false|C1553498|home health encounter|home
Finding|Body Substance|Hospital Course|3178,3185|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|3178,3185|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|3178,3185|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Attribute|Clinical Attribute|Hospital Course|3190,3195|false|false|false|C5890168||alert
Drug|Organic Chemical|Hospital Course|3190,3195|false|false|false|C0718338|Alert brand of caffeine|alert
Drug|Pharmacologic Substance|Hospital Course|3190,3195|false|false|false|C0718338|Alert brand of caffeine|alert
Event|Event|Hospital Course|3190,3195|false|false|false|||alert
Finding|Finding|Hospital Course|3190,3195|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Functional Concept|Hospital Course|3190,3195|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Intellectual Product|Hospital Course|3190,3195|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Event|Event|Hospital Course|3200,3208|false|false|false|||oriented
Finding|Finding|Hospital Course|3200,3208|false|false|false|C1961028|Oriented to place|oriented
Event|Event|Hospital Course|3221,3236|false|false|false|||hospitalization
Procedure|Health Care Activity|Hospital Course|3221,3236|false|false|false|C0019993|Hospitalization|hospitalization
Attribute|Clinical Attribute|Hospital Course|3238,3242|false|false|false|C2598155||pain
Event|Event|Hospital Course|3238,3242|false|false|false|||pain
Finding|Functional Concept|Hospital Course|3238,3242|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|3238,3242|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|3257,3264|false|false|false|||managed
Drug|Organic Chemical|Hospital Course|3270,3278|false|false|false|C0728755|Dilaudid|dilaudid
Drug|Pharmacologic Substance|Hospital Course|3270,3278|false|false|false|C0728755|Dilaudid|dilaudid
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|3279,3282|false|false|false|C0149576|Structure of posterior cerebral artery|PCA
Disorder|Disease or Syndrome|Hospital Course|3279,3282|false|false|false|C0268398;C4275079|Familial lichen amyloidosis;Posterior cortical atrophy syndrome|PCA
Drug|Amino Acid, Peptide, or Protein|Hospital Course|3279,3282|false|false|false|C0030131;C0034330|p-Chloroamphetamine;pyrrolidonecarboxylic acid|PCA
Drug|Biologically Active Substance|Hospital Course|3279,3282|false|false|false|C0030131;C0034330|p-Chloroamphetamine;pyrrolidonecarboxylic acid|PCA
Drug|Indicator, Reagent, or Diagnostic Aid|Hospital Course|3279,3282|false|false|false|C0030131;C0034330|p-Chloroamphetamine;pyrrolidonecarboxylic acid|PCA
Drug|Organic Chemical|Hospital Course|3279,3282|false|false|false|C0030131;C0034330|p-Chloroamphetamine;pyrrolidonecarboxylic acid|PCA
Drug|Pharmacologic Substance|Hospital Course|3279,3282|false|false|false|C0030131;C0034330|p-Chloroamphetamine;pyrrolidonecarboxylic acid|PCA
Event|Event|Hospital Course|3279,3282|false|false|false|||PCA
Finding|Finding|Hospital Course|3279,3282|false|false|false|C0220723;C1549860;C1836722|CHOANAL ATRESIA, POSTERIOR;FLVCR1 gene;PCA Message Structure|PCA
Finding|Gene or Genome|Hospital Course|3279,3282|false|false|false|C0220723;C1549860;C1836722|CHOANAL ATRESIA, POSTERIOR;FLVCR1 gene;PCA Message Structure|PCA
Finding|Intellectual Product|Hospital Course|3279,3282|false|false|false|C0220723;C1549860;C1836722|CHOANAL ATRESIA, POSTERIOR;FLVCR1 gene;PCA Message Structure|PCA
Procedure|Laboratory Procedure|Hospital Course|3279,3282|false|false|false|C0030625;C0078944;C5968782|Passive Cutaneous Anaphylaxis;Patient controlled intravenous analgesia;Patient-Controlled Analgesia|PCA
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3279,3282|false|false|false|C0030625;C0078944;C5968782|Passive Cutaneous Anaphylaxis;Patient controlled intravenous analgesia;Patient-Controlled Analgesia|PCA
Event|Event|Hospital Course|3301,3306|false|false|false|||using
Finding|Intellectual Product|Hospital Course|3311,3315|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|Hospital Course|3316,3328|false|false|false|||transitioned
Drug|Organic Chemical|Hospital Course|3332,3340|false|false|false|C0040610|tramadol|tramadol
Drug|Pharmacologic Substance|Hospital Course|3332,3340|false|false|false|C0040610|tramadol|tramadol
Event|Event|Hospital Course|3332,3340|false|false|false|||tramadol
Procedure|Laboratory Procedure|Hospital Course|3332,3340|false|false|false|C1266765|Tramadol measurement (procedure)|tramadol
Attribute|Clinical Attribute|Hospital Course|3370,3374|false|false|false|C2598155||Pain
Event|Event|Hospital Course|3370,3374|false|false|false|||Pain
Finding|Functional Concept|Hospital Course|3370,3374|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Hospital Course|3370,3374|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Finding|Hospital Course|3379,3388|false|false|false|C5202951;C5202952;C5202953|Can Do Very Well;Describes Very Well;Very Well|very well
Finding|Finding|Hospital Course|3384,3388|false|false|false|C5575035|Well (answer to question)|well
Event|Event|Hospital Course|3389,3399|false|false|false|||controlled
Finding|Body Substance|Hospital Course|3411,3418|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|3411,3418|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|3411,3418|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|3419,3427|false|false|false|||remained
Event|Event|Hospital Course|3428,3434|false|false|false|||stable
Finding|Intellectual Product|Hospital Course|3428,3434|false|false|false|C1547311|Patient Condition Code - Stable|stable
Anatomy|Body System|Hospital Course|3442,3456|false|false|false|C0007226;C3887460|Cardiovascular;Cardiovascular system|cardiovascular
Drug|Food|Hospital Course|3470,3475|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|vital
Attribute|Clinical Attribute|Hospital Course|3470,3481|false|false|false|C0488614;C0518766|Vital signs|vital signs
Procedure|Health Care Activity|Hospital Course|3470,3481|false|false|false|C0150404|Taking vital signs|vital signs
Event|Event|Hospital Course|3476,3481|false|false|false|||signs
Finding|Finding|Hospital Course|3476,3481|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Hospital Course|3476,3481|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Event|Event|Hospital Course|3497,3506|false|false|false|||monitored
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|3512,3521|false|false|false|C0024109|Lung|PULMONARY
Attribute|Clinical Attribute|Hospital Course|3512,3521|false|false|false|C2707265||PULMONARY
Finding|Finding|Hospital Course|3512,3521|false|false|false|C4522268|Pulmonary (intended site)|PULMONARY
Finding|Body Substance|Hospital Course|3527,3534|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|3527,3534|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|3527,3534|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|3535,3543|false|false|false|||remained
Event|Event|Hospital Course|3544,3550|false|false|false|||stable
Finding|Intellectual Product|Hospital Course|3544,3550|false|false|false|C1547311|Patient Condition Code - Stable|stable
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|3558,3567|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Hospital Course|3558,3567|false|false|false|C2707265||pulmonary
Finding|Finding|Hospital Course|3558,3567|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Drug|Food|Hospital Course|3581,3586|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|vital
Attribute|Clinical Attribute|Hospital Course|3581,3592|false|false|false|C0488614;C0518766|Vital signs|vital signs
Procedure|Health Care Activity|Hospital Course|3581,3592|false|false|false|C0150404|Taking vital signs|vital signs
Event|Event|Hospital Course|3587,3592|false|false|false|||signs
Finding|Finding|Hospital Course|3587,3592|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Hospital Course|3587,3592|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Event|Event|Hospital Course|3608,3617|false|false|false|||monitored
Finding|Idea or Concept|Hospital Course|3619,3623|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|Good
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|3624,3633|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Hospital Course|3624,3633|false|false|false|C2707265||pulmonary
Finding|Finding|Hospital Course|3624,3633|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Event|Event|Hospital Course|3635,3641|false|false|false|||toilet
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3635,3641|false|false|false|C0184958|Toilet procedure|toilet
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3643,3659|false|false|false|C0013457|Early Ambulation|early ambulation
Event|Event|Hospital Course|3649,3659|false|false|false|||ambulation
Finding|Daily or Recreational Activity|Hospital Course|3649,3659|false|false|false|C0080331;C0945826|Ambulation;Walking (function)|ambulation
Finding|Functional Concept|Hospital Course|3649,3659|false|false|false|C0080331;C0945826|Ambulation;Walking (function)|ambulation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3664,3684|false|false|false|C0454512|Incentive spirometry|incentive spirometry
Event|Event|Hospital Course|3674,3684|false|false|false|||spirometry
Procedure|Diagnostic Procedure|Hospital Course|3674,3684|false|false|false|C0037981|Spirometry|spirometry
Event|Event|Hospital Course|3691,3701|false|false|false|||encouraged
Event|Event|Hospital Course|3713,3728|false|false|false|||hospitalization
Procedure|Health Care Activity|Hospital Course|3713,3728|false|false|false|C0019993|Hospitalization|hospitalization
Attribute|Clinical Attribute|Hospital Course|3756,3765|false|false|false|C0945766||procedure
Event|Event|Hospital Course|3756,3765|false|false|false|||procedure
Event|Occupational Activity|Hospital Course|3756,3765|false|false|false|C1546467|Act Class - procedure|procedure
Finding|Functional Concept|Hospital Course|3756,3765|false|false|false|C2700391|Procedure (set of actions)|procedure
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3756,3765|false|false|false|C0184661|Interventional procedure|procedure
Event|Event|Hospital Course|3766,3773|false|false|false|||started
Event|Event|Hospital Course|3788,3794|false|false|false|||unable
Finding|Finding|Hospital Course|3788,3794|false|false|false|C1299582|Unable|unable
Event|Event|Hospital Course|3799,3803|false|false|false|||pass
Finding|Finding|Hospital Course|3799,3803|false|false|false|C2828386|Pass (indicator)|pass
Event|Event|Hospital Course|3816,3823|false|false|false|||attempt
Event|Event|Hospital Course|3816,3823|false|false|false|C1516084|Attempt|attempt
Event|Event|Hospital Course|3829,3837|false|false|false|||standard
Finding|Idea or Concept|Hospital Course|3829,3837|false|false|false|C1548173;C2828392|Standard (document);Type of Agreement - Standard|standard
Finding|Intellectual Product|Hospital Course|3829,3837|false|false|false|C1548173;C2828392|Standard (document);Type of Agreement - Standard|standard
Procedure|Laboratory Procedure|Hospital Course|3829,3837|false|false|false|C3873211|Standard base excess calculation technique|standard
Event|Event|Hospital Course|3848,3852|false|false|false|||type
Finding|Gene or Genome|Hospital Course|3848,3852|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Intellectual Product|Hospital Course|3848,3852|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Finding|Hospital Course|3874,3881|false|false|false|C0021359;C4074771|Infertility;Sterility, Reproductive|sterile
Finding|Pathologic Function|Hospital Course|3874,3881|false|false|false|C0021359;C4074771|Infertility;Sterility, Reproductive|sterile
Event|Event|Hospital Course|3882,3891|false|false|false|||technique
Finding|Functional Concept|Hospital Course|3882,3891|false|false|false|C0449851|Techniques|technique
Event|Event|Hospital Course|3906,3911|false|false|false|||foley
Event|Event|Hospital Course|3913,3922|false|false|false|||placement
Procedure|Health Care Activity|Hospital Course|3913,3922|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3913,3922|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Event|Event|Hospital Course|3941,3952|false|false|false|||application
Finding|Functional Concept|Hospital Course|3941,3952|false|false|false|C0870325;C1547755;C1947919;C2347934;C4048755|Application Document;Apply;Computer Application;HL7 Version 2.5 - Application;Regulatory Application|application
Finding|Idea or Concept|Hospital Course|3941,3952|false|false|false|C0870325;C1547755;C1947919;C2347934;C4048755|Application Document;Apply;Computer Application;HL7 Version 2.5 - Application;Regulatory Application|application
Finding|Intellectual Product|Hospital Course|3941,3952|false|false|false|C0870325;C1547755;C1947919;C2347934;C4048755|Application Document;Apply;Computer Application;HL7 Version 2.5 - Application;Regulatory Application|application
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3941,3952|false|false|false|C0185125|Application procedure|application
Finding|Gene or Genome|Hospital Course|3977,3981|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Intellectual Product|Hospital Course|3977,3981|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Event|Event|Hospital Course|3982,3991|false|false|false|||catheters
Event|Event|Hospital Course|4005,4011|false|false|false|||unable
Finding|Finding|Hospital Course|4005,4011|false|false|false|C1299582|Unable|unable
Event|Event|Hospital Course|4019,4025|false|false|false|||passed
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4031,4039|false|false|false|C0033572;C4266527|Prostate;Structure of prostate (body structure)|prostate
Disorder|Disease or Syndrome|Hospital Course|4031,4039|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|prostate
Disorder|Neoplastic Process|Hospital Course|4031,4039|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|prostate
Event|Event|Hospital Course|4031,4039|false|false|false|||prostate
Event|Event|Hospital Course|4053,4062|false|false|false|||consulted
Event|Event|Hospital Course|4105,4118|false|false|false|||demonstrating
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4128,4135|false|false|false|C0041967|Urethra|urethra
Disorder|Disease or Syndrome|Hospital Course|4128,4135|false|false|false|C0041969;C0153620;C0154019;C0496929|Benign neoplasm of urethra;Malignant neoplasm of urethra;Neoplasm of uncertain or unknown behavior of urethra;Urethral Diseases|urethra
Disorder|Neoplastic Process|Hospital Course|4128,4135|false|false|false|C0041969;C0153620;C0154019;C0496929|Benign neoplasm of urethra;Malignant neoplasm of urethra;Neoplasm of uncertain or unknown behavior of urethra;Urethral Diseases|urethra
Event|Event|Hospital Course|4128,4135|false|false|false|||urethra
Finding|Body Substance|Hospital Course|4128,4135|false|false|false|C1547951;C1550675|Urethra specimen;Urethra specimen code|urethra
Finding|Intellectual Product|Hospital Course|4128,4135|false|false|false|C1547951;C1550675|Urethra specimen;Urethra specimen code|urethra
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4128,4135|false|false|false|C0810170|Procedure on urethra|urethra
Event|Event|Hospital Course|4145,4153|false|false|false|||flexible
Event|Event|Hospital Course|4155,4164|false|false|false|||guidewire
Event|Event|Hospital Course|4166,4176|false|false|false|||cystoscope
Event|Event|Hospital Course|4181,4189|false|false|false|||advanced
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4199,4206|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|Hospital Course|4199,4206|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4199,4206|false|false|false|C0872388|Procedures on bladder|bladder
Finding|Conceptual Entity|Hospital Course|4212,4217|false|false|false|C1710028|Scope|scope
Event|Event|Hospital Course|4223,4232|false|false|false|||withdrawn
Event|Event|Hospital Course|4243,4250|false|false|false|||council
Event|Event|Hospital Course|4255,4263|false|false|false|||advanced
Finding|Gene or Genome|Hospital Course|4273,4277|false|false|false|C1823858|WIPF2 gene|wire
Event|Event|Hospital Course|4280,4286|false|false|false|||passed
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4291,4299|false|false|false|C0033572;C4266527|Prostate;Structure of prostate (body structure)|prostate
Disorder|Disease or Syndrome|Hospital Course|4291,4299|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|prostate
Disorder|Neoplastic Process|Hospital Course|4291,4299|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|prostate
Event|Event|Hospital Course|4291,4299|false|false|false|||prostate
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4313,4320|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|Hospital Course|4313,4320|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Event|Event|Hospital Course|4313,4320|false|false|false|||bladder
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4313,4320|false|false|false|C0872388|Procedures on bladder|bladder
Finding|Body Substance|Hospital Course|4326,4333|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|4326,4333|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|4326,4333|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|4339,4349|false|false|false|||discharged
Event|Activity|Hospital Course|4368,4373|false|false|false|C1882509|put - instruction imperative|place
Event|Event|Hospital Course|4368,4373|false|false|false|||place
Finding|Functional Concept|Hospital Course|4368,4373|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|Hospital Course|4368,4373|false|false|false|C1533810||place
Attribute|Clinical Attribute|Hospital Course|4379,4391|false|false|false|C3263700||instructions
Event|Event|Hospital Course|4379,4391|false|false|false|||instructions
Finding|Intellectual Product|Hospital Course|4379,4391|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|instructions
Event|Event|Hospital Course|4396,4402|false|false|false|||follow
Event|Event|Hospital Course|4422,4432|false|false|false|||outpatient
Finding|Classification|Hospital Course|4422,4432|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|4422,4432|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Functional Concept|Hospital Course|4455,4462|false|false|false|C0042034;C4067975|Urination;Voids|voiding
Finding|Organism Function|Hospital Course|4455,4462|false|false|false|C0042034;C4067975|Urination;Voids|voiding
Event|Event|Hospital Course|4463,4468|false|false|false|||trial
Procedure|Research Activity|Hospital Course|4463,4468|false|false|false|C0008976|Clinical Trials|trial
Drug|Antibiotic|Hospital Course|4473,4484|true|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|Hospital Course|4473,4484|false|false|false|||antibiotics
Event|Event|Hospital Course|4490,4502|false|false|false|||administered
Finding|Body Substance|Hospital Course|4508,4515|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|4508,4515|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|4508,4515|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|4521,4531|false|false|false|||tolerating
Finding|Daily or Recreational Activity|Hospital Course|4534,4546|false|false|false|C0184625||regular diet
Drug|Food|Hospital Course|4542,4546|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|Hospital Course|4542,4546|false|false|false|||diet
Finding|Functional Concept|Hospital Course|4542,4546|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|Hospital Course|4542,4546|false|false|false|C0012159|Diet therapy|diet
Event|Event|Hospital Course|4556,4565|false|false|false|||discharge
Finding|Body Substance|Hospital Course|4556,4565|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|4556,4565|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|4556,4565|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|4556,4565|false|false|false|C0030685|Patient Discharge|discharge
Finding|Body Substance|Hospital Course|4578,4585|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|4578,4585|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|4578,4585|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|Hospital Course|4588,4593|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|Hospital Course|4588,4593|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|Hospital Course|4594,4600|false|false|false|||curves
Event|Event|Hospital Course|4614,4621|false|false|false|||watched
Event|Event|Hospital Course|4626,4631|false|false|false|||signs
Finding|Finding|Hospital Course|4626,4631|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Hospital Course|4626,4631|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Disorder|Disease or Syndrome|Hospital Course|4636,4645|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|Hospital Course|4636,4645|false|false|false|||infection
Finding|Pathologic Function|Hospital Course|4636,4645|false|false|false|C3714514|Infection|infection
Event|Event|Hospital Course|4667,4671|false|false|false|||none
Drug|Biologically Active Substance|Hospital Course|4677,4681|false|false|false|C0018966|Heme|HEME
Drug|Organic Chemical|Hospital Course|4677,4681|false|false|false|C0018966|Heme|HEME
Event|Event|Hospital Course|4677,4681|false|false|false|||HEME
Finding|Body Substance|Hospital Course|4683,4690|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|4683,4690|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|4683,4690|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|4691,4699|false|false|false|||received
Disorder|Mental or Behavioral Dysfunction|Hospital Course|4700,4703|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4700,4703|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|4700,4703|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|4700,4703|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|4700,4703|false|false|false|C1332410|BID gene|BID
Event|Event|Hospital Course|4704,4707|false|false|false|||SQH
Anatomy|Body Location or Region|Hospital Course|4712,4715|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Hospital Course|4712,4715|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Hospital Course|4712,4715|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4712,4727|false|false|false|C0853245|DVT prophylaxis|DVT prophylaxis
Event|Event|Hospital Course|4716,4727|false|false|false|||prophylaxis
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4716,4727|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Event|Event|Hospital Course|4732,4740|false|false|false|||addition
Finding|Functional Concept|Hospital Course|4732,4740|false|false|false|C0332287;C1883712|Add - instruction imperative;In addition to|addition
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4757,4773|false|false|false|C0013457|Early Ambulation|early ambulation
Event|Event|Hospital Course|4763,4773|false|false|false|||ambulation
Finding|Daily or Recreational Activity|Hospital Course|4763,4773|false|false|false|C0080331;C0945826|Ambulation;Walking (function)|ambulation
Finding|Functional Concept|Hospital Course|4763,4773|false|false|false|C0080331;C0945826|Ambulation;Walking (function)|ambulation
Event|Event|Hospital Course|4787,4798|false|false|false|||compression
Finding|Functional Concept|Hospital Course|4787,4798|false|false|false|C0332459;C4551657|Compressed structure|compression
Phenomenon|Natural Phenomenon or Process|Hospital Course|4787,4798|false|false|false|C0728907|Compression|compression
Procedure|Machine Activity|Hospital Course|4787,4798|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4787,4798|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Event|Event|Hospital Course|4800,4807|false|false|false|||devices
Finding|Gene or Genome|Hospital Course|4812,4816|false|false|false|C1420638;C1539127;C1710283|CORO7 gene;TCF21 gene;TCF21 wt Allele|POD1
Finding|Body Substance|Hospital Course|4821,4828|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|4821,4828|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|4821,4828|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|4833,4842|false|false|false|||restarted
Event|Event|Hospital Course|4850,4854|false|false|false|||home
Finding|Idea or Concept|Hospital Course|4850,4854|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|4850,4854|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|4850,4854|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|4856,4866|false|false|false|C0206460|enoxaparin|enoxaparin
Drug|Pharmacologic Substance|Hospital Course|4856,4866|false|false|false|C0206460|enoxaparin|enoxaparin
Event|Event|Hospital Course|4856,4866|false|false|false|||enoxaparin
Event|Event|Hospital Course|4874,4883|false|false|false|||discharge
Finding|Body Substance|Hospital Course|4874,4883|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|4874,4883|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|4874,4883|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|4874,4883|false|false|false|C0030685|Patient Discharge|discharge
Finding|Idea or Concept|Hospital Course|4887,4899|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Event|Event|Hospital Course|4900,4906|false|false|false|||ISSUES
Finding|Finding|Hospital Course|4936,4940|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Hospital Course|4936,4940|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Hospital Course|4936,4940|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|Hospital Course|4944,4953|false|false|false|||discharge
Finding|Body Substance|Hospital Course|4944,4953|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|4944,4953|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|4944,4953|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|4944,4953|false|false|false|C0030685|Patient Discharge|discharge
Finding|Body Substance|Hospital Course|4959,4966|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|4959,4966|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|4959,4966|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|4977,4981|false|false|false|||well
Finding|Finding|Hospital Course|4977,4981|false|false|false|C5575035|Well (answer to question)|well
Event|Event|Hospital Course|4983,4991|false|false|false|||afebrile
Finding|Finding|Hospital Course|4983,4991|false|false|false|C0277797|Apyrexial|afebrile
Event|Event|Hospital Course|4998,5004|false|false|false|||stable
Finding|Intellectual Product|Hospital Course|4998,5004|false|false|false|C1547311|Patient Condition Code - Stable|stable
Drug|Food|Hospital Course|5005,5010|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|vital
Attribute|Clinical Attribute|Hospital Course|5005,5016|false|false|false|C0488614;C0518766|Vital signs|vital signs
Procedure|Health Care Activity|Hospital Course|5005,5016|false|false|false|C0150404|Taking vital signs|vital signs
Event|Event|Hospital Course|5011,5016|false|false|false|||signs
Finding|Finding|Hospital Course|5011,5016|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Hospital Course|5011,5016|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Body Substance|Hospital Course|5022,5029|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|5022,5029|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|5022,5029|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|5034,5044|false|false|false|||tolerating
Drug|Food|Hospital Course|5045,5049|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|Hospital Course|5045,5049|false|false|false|||diet
Finding|Functional Concept|Hospital Course|5045,5049|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|Hospital Course|5045,5049|false|false|false|C0012159|Diet therapy|diet
Anatomy|Body Space or Junction|Hospital Course|5064,5068|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|5064,5068|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|5064,5068|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|5064,5068|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|Hospital Course|5070,5080|false|false|false|||ambulating
Attribute|Clinical Attribute|Hospital Course|5086,5090|false|false|false|C2598155||pain
Event|Event|Hospital Course|5086,5090|false|false|false|||pain
Finding|Functional Concept|Hospital Course|5086,5090|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|5086,5090|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Hospital Course|5095,5099|false|false|false|C5575035|Well (answer to question)|well
Event|Event|Hospital Course|5100,5110|false|false|false|||controlled
Finding|Body Substance|Hospital Course|5117,5124|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|5117,5124|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|5117,5124|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|5129,5139|false|false|false|||discharged
Event|Event|Hospital Course|5140,5144|false|false|false|||home
Finding|Idea or Concept|Hospital Course|5140,5144|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|5140,5144|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|5140,5144|false|false|false|C1553498|home health encounter|home
Event|Event|Hospital Course|5160,5168|false|false|false|||catheter
Finding|Intellectual Product|Hospital Course|5160,5168|false|false|false|C1546572||catheter
Event|Event|Hospital Course|5187,5195|false|false|false|||teaching
Finding|Intellectual Product|Hospital Course|5187,5195|false|false|false|C1548344|Visit User Code - Teaching|teaching
Procedure|Educational Activity|Hospital Course|5187,5195|false|false|false|C0039401;C0220924|Education (procedure);Teaching aspects|teaching
Event|Activity|Hospital Course|5200,5204|false|false|false|C1947933|care activity|care
Event|Event|Hospital Course|5200,5204|false|false|false|||care
Finding|Finding|Hospital Course|5200,5204|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Hospital Course|5200,5204|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Body Substance|Hospital Course|5210,5217|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|5210,5217|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|5210,5217|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|5227,5236|false|false|false|||discharge
Finding|Body Substance|Hospital Course|5227,5236|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|5227,5236|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|5227,5236|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|5227,5236|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|Hospital Course|5238,5246|false|false|false|||teaching
Finding|Intellectual Product|Hospital Course|5238,5246|false|false|false|C1548344|Visit User Code - Teaching|teaching
Procedure|Educational Activity|Hospital Course|5238,5246|false|false|false|C0039401;C0220924|Education (procedure);Teaching aspects|teaching
Event|Event|Hospital Course|5251,5257|false|false|false|||follow
Attribute|Clinical Attribute|Hospital Course|5261,5273|false|false|false|C3263700||instructions
Event|Event|Hospital Course|5261,5273|false|false|false|||instructions
Finding|Intellectual Product|Hospital Course|5261,5273|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|instructions
Event|Event|Hospital Course|5279,5292|false|false|false|||understanding
Finding|Mental Process|Hospital Course|5279,5292|false|false|false|C0162340|Comprehension|understanding
Event|Event|Hospital Course|5294,5304|false|false|false|||verbalized
Attribute|Clinical Attribute|Hospital Course|5309,5318|false|false|false|C4255433||agreement
Event|Event|Hospital Course|5309,5318|false|false|false|||agreement
Finding|Intellectual Product|Hospital Course|5309,5318|false|false|false|C0680240;C4255373|Agreement;Agreement (document)|agreement
Finding|Social Behavior|Hospital Course|5309,5318|false|false|false|C0680240;C4255373|Agreement;Agreement (document)|agreement
Event|Event|Hospital Course|5328,5337|false|false|false|||discharge
Finding|Body Substance|Hospital Course|5328,5337|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|5328,5337|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|5328,5337|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|5328,5337|false|false|false|C0030685|Patient Discharge|discharge
Attribute|Clinical Attribute|Hospital Course|5328,5342|false|false|false|C2745873||discharge plan
Finding|Intellectual Product|Hospital Course|5328,5342|false|false|false|C2735970|Discharge plan|discharge plan
Procedure|Health Care Activity|Hospital Course|5328,5342|false|false|false|C0012622|Discharge Planning|discharge plan
Disorder|Disease or Syndrome|Hospital Course|5338,5342|false|false|false|C0270724|Infantile Neuroaxonal Dystrophy|plan
Event|Event|Hospital Course|5338,5342|false|false|false|||plan
Finding|Functional Concept|Hospital Course|5338,5342|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Intellectual Product|Hospital Course|5338,5342|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Mental Process|Hospital Course|5338,5342|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Attribute|Clinical Attribute|Hospital Course|5346,5357|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|5346,5357|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|5346,5357|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|5346,5357|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|5346,5370|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|5361,5370|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|5361,5370|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|Hospital Course|5372,5383|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|5372,5383|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|5372,5383|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|5372,5383|false|false|false|C4284232|Medications|Medications
Attribute|Clinical Attribute|Hospital Course|5386,5398|false|false|false|C5886759|Prescription (attribute)|Prescription
Event|Event|Hospital Course|5386,5398|false|false|false|||Prescription
Finding|Intellectual Product|Hospital Course|5386,5398|false|false|false|C1521941|prescription document|Prescription
Procedure|Health Care Activity|Hospital Course|5386,5398|false|false|false|C0033080|Prescription (procedure)|Prescription
Drug|Hormone|Hospital Course|5399,5409|false|false|false|C1878933|Bio-Throid|BIO-THROID
Drug|Organic Chemical|Hospital Course|5399,5409|false|false|false|C1878933|Bio-Throid|BIO-THROID
Drug|Pharmacologic Substance|Hospital Course|5399,5409|false|false|false|C1878933|Bio-Throid|BIO-THROID
Drug|Hormone|Hospital Course|5412,5422|false|false|false|C1878933|Bio-Throid|Bio-Throid
Drug|Organic Chemical|Hospital Course|5412,5422|false|false|false|C1878933|Bio-Throid|Bio-Throid
Drug|Pharmacologic Substance|Hospital Course|5412,5422|false|false|false|C1878933|Bio-Throid|Bio-Throid
Event|Event|Hospital Course|5412,5422|false|false|false|||Bio-Throid
Finding|Intellectual Product|Hospital Course|5433,5437|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|5433,5443|false|false|false|C3537736|Once A Day|once a day
Event|Event|Hospital Course|5440,5443|false|false|false|||day
Finding|Idea or Concept|Hospital Course|5440,5443|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|5440,5443|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|5448,5458|false|false|false|||Prescribed
Finding|Functional Concept|Hospital Course|5469,5477|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|Provider
Finding|Intellectual Product|Hospital Course|5469,5477|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|Provider
Drug|Organic Chemical|Hospital Course|5479,5489|false|false|false|C0206460|enoxaparin|ENOXAPARIN
Drug|Pharmacologic Substance|Hospital Course|5479,5489|false|false|false|C0206460|enoxaparin|ENOXAPARIN
Event|Event|Hospital Course|5479,5489|false|false|false|||ENOXAPARIN
Drug|Organic Chemical|Hospital Course|5492,5502|false|false|false|C0206460|enoxaparin|enoxaparin
Drug|Pharmacologic Substance|Hospital Course|5492,5502|false|false|false|C0206460|enoxaparin|enoxaparin
Event|Event|Hospital Course|5492,5502|false|false|false|||enoxaparin
Finding|Functional Concept|Hospital Course|5517,5529|false|false|false|C1522438|Subcutaneous Route of Administration|subcutaneous
Event|Event|Hospital Course|5530,5537|false|false|false|||syringe
Drug|Organic Chemical|Hospital Course|5556,5566|false|false|false|C0028978|omeprazole|OMEPRAZOLE
Drug|Pharmacologic Substance|Hospital Course|5556,5566|false|false|false|C0028978|omeprazole|OMEPRAZOLE
Drug|Organic Chemical|Hospital Course|5569,5579|false|false|false|C0028978|omeprazole|omeprazole
Drug|Pharmacologic Substance|Hospital Course|5569,5579|false|false|false|C0028978|omeprazole|omeprazole
Event|Event|Hospital Course|5569,5579|false|false|false|||omeprazole
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5586,5593|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|Hospital Course|5586,5593|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|Hospital Course|5586,5593|false|false|false|C0006935|capsule (pharmacologic)|capsule
Event|Event|Hospital Course|5594,5601|false|false|false|||delayed
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5614,5621|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|Hospital Course|5614,5621|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|Hospital Course|5614,5621|false|false|false|C0006935|capsule (pharmacologic)|capsule
Finding|Functional Concept|Hospital Course|5625,5633|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|5628,5633|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|5628,5633|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Organic Chemical|Hospital Course|5646,5655|false|false|false|C0077656|ubiquinol|UBIQUINOL
Drug|Pharmacologic Substance|Hospital Course|5646,5655|false|false|false|C0077656|ubiquinol|UBIQUINOL
Drug|Organic Chemical|Hospital Course|5658,5667|false|false|false|C0077656|ubiquinol|ubiquinol
Drug|Pharmacologic Substance|Hospital Course|5658,5667|false|false|false|C0077656|ubiquinol|ubiquinol
Event|Event|Hospital Course|5658,5667|false|false|false|||ubiquinol
Anatomy|Body Location or Region|Hospital Course|5687,5692|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|5687,5692|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|Hospital Course|5701,5704|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|5701,5704|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|5710,5720|false|false|false|||Prescribed
Finding|Functional Concept|Hospital Course|5730,5738|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|Provider
Finding|Intellectual Product|Hospital Course|5730,5738|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|Provider
Attribute|Clinical Attribute|Hospital Course|5742,5753|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|5742,5753|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|5742,5753|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|5742,5753|false|false|false|C4284232|Medications|Medications
Drug|Pharmacologic Substance|Hospital Course|5756,5759|false|false|false|C0013231|Drugs, Non-Prescription|OTC
Event|Event|Hospital Course|5756,5759|false|false|false|||OTC
Finding|Gene or Genome|Hospital Course|5756,5759|false|false|false|C1418193|OTC gene|OTC
Drug|Element, Ion, or Isotope|Hospital Course|5760,5767|false|false|false|C2346592|Ferrous|FERROUS
Drug|Inorganic Chemical|Hospital Course|5760,5775|false|false|false|C0060282|ferrous sulfate|FERROUS SULFATE
Drug|Pharmacologic Substance|Hospital Course|5760,5775|false|false|false|C0060282|ferrous sulfate|FERROUS SULFATE
Drug|Element, Ion, or Isotope|Hospital Course|5768,5775|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|SULFATE
Drug|Inorganic Chemical|Hospital Course|5768,5775|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|SULFATE
Drug|Pharmacologic Substance|Hospital Course|5768,5775|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|SULFATE
Drug|Element, Ion, or Isotope|Hospital Course|5778,5785|false|false|false|C2346592|Ferrous|ferrous
Drug|Inorganic Chemical|Hospital Course|5778,5793|false|false|false|C0060282|ferrous sulfate|ferrous sulfate
Drug|Pharmacologic Substance|Hospital Course|5778,5793|false|false|false|C0060282|ferrous sulfate|ferrous sulfate
Drug|Element, Ion, or Isotope|Hospital Course|5786,5793|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|Hospital Course|5786,5793|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|Hospital Course|5786,5793|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Event|Event|Hospital Course|5786,5793|false|false|false|||sulfate
Drug|Biologically Active Substance|Hospital Course|5808,5812|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|Hospital Course|5808,5812|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|Hospital Course|5808,5812|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Procedure|Laboratory Procedure|Hospital Course|5808,5812|false|false|false|C0337439|Iron measurement|iron
Drug|Biomedical or Dental Material|Hospital Course|5825,5831|false|false|false|C0039225|Tablet Dosage Form|tablet
Event|Event|Hospital Course|5825,5831|false|false|false|||tablet
Finding|Functional Concept|Hospital Course|5835,5843|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|5838,5843|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|5838,5843|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|Hospital Course|5852,5855|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|5852,5855|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|5860,5870|false|false|false|||Prescribed
Finding|Functional Concept|Hospital Course|5880,5888|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|Provider
Finding|Intellectual Product|Hospital Course|5880,5888|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|Provider
Event|Event|Hospital Course|5904,5915|false|false|false|||COMBINATION
Finding|Finding|Hospital Course|5904,5915|false|false|false|C3811910|combination - answer to question|COMBINATION
Event|Event|Hospital Course|5942,5951|false|false|false|||uncertain
Finding|Finding|Hospital Course|5942,5951|false|false|false|C0087130|Uncertainty|uncertain
Event|Event|Hospital Course|5957,5967|false|false|false|||Prescribed
Finding|Functional Concept|Hospital Course|5977,5985|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|Provider
Finding|Intellectual Product|Hospital Course|5977,5985|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|Provider
Event|Event|Hospital Course|5996,6005|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|5996,6005|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|5996,6005|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|5996,6005|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|5996,6005|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|5996,6017|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|6006,6017|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|6006,6017|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|6006,6017|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|6006,6017|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|6023,6036|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|6023,6036|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Hospital Course|6023,6036|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|6023,6036|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Event|Event|Hospital Course|6048,6051|false|false|false|||TID
Drug|Organic Chemical|Hospital Course|6058,6066|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|6058,6066|false|false|false|C1692318|docusate|Docusate
Event|Event|Hospital Course|6058,6066|false|false|false|||Docusate
Drug|Organic Chemical|Hospital Course|6058,6073|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|Hospital Course|6058,6073|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|Hospital Course|6067,6073|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|6067,6073|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|6067,6073|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|6067,6073|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|6067,6073|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|6067,6073|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6084,6087|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6084,6087|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|6084,6087|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|6084,6087|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|6084,6087|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|6094,6099|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|Hospital Course|6094,6099|false|false|false|C3489575|sennosides, USP|Senna
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6110,6113|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6110,6113|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|6110,6113|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|6110,6113|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|6110,6113|false|false|false|C1332410|BID gene|BID
Finding|Gene or Genome|Hospital Course|6114,6117|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Sign or Symptom|Hospital Course|6118,6130|false|false|false|C0009806|Constipation|Constipation
Drug|Biologically Active Substance|Hospital Course|6139,6143|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Hospital Course|6139,6143|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Drug|Substance|Hospital Course|6139,6143|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Event|Event|Hospital Course|6139,6143|false|false|false|||Line
Finding|Intellectual Product|Hospital Course|6139,6143|false|false|false|C1546701|line source specimen code|Line
Drug|Organic Chemical|Hospital Course|6150,6158|false|false|false|C0040610|tramadol|TraMADol
Drug|Pharmacologic Substance|Hospital Course|6150,6158|false|false|false|C0040610|tramadol|TraMADol
Event|Event|Hospital Course|6150,6158|false|false|false|||TraMADol
Procedure|Laboratory Procedure|Hospital Course|6150,6158|false|false|false|C1266765|Tramadol measurement (procedure)|TraMADol
Finding|Gene or Genome|Hospital Course|6172,6175|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|6176,6180|false|false|false|C2598155||Pain
Event|Event|Hospital Course|6176,6180|false|false|false|||Pain
Finding|Functional Concept|Hospital Course|6176,6180|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Hospital Course|6176,6180|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Finding|Hospital Course|6183,6191|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|Hospital Course|6183,6191|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Drug|Pharmacologic Substance|Hospital Course|6198,6208|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Hospital Course|6198,6208|false|false|false|||medication
Finding|Intellectual Product|Hospital Course|6198,6208|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Finding|Finding|Hospital Course|6214,6217|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Hospital Course|6214,6217|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Drug|Hazardous or Poisonous Substance|Hospital Course|6223,6231|false|false|false|C0027415|Narcotics|narcotic
Drug|Pharmacologic Substance|Hospital Course|6223,6231|false|false|false|C0027415|Narcotics|narcotic
Event|Event|Hospital Course|6223,6231|false|false|false|||narcotic
Event|Event|Hospital Course|6240,6245|false|false|false|||cause
Finding|Conceptual Entity|Hospital Course|6240,6245|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Finding|Functional Concept|Hospital Course|6240,6245|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Event|Event|Hospital Course|6247,6259|false|false|false|||constipation
Finding|Sign or Symptom|Hospital Course|6247,6259|false|false|false|C0009806|Constipation|constipation
Drug|Organic Chemical|Hospital Course|6266,6274|false|false|false|C0040610|tramadol|tramadol
Drug|Pharmacologic Substance|Hospital Course|6266,6274|false|false|false|C0040610|tramadol|tramadol
Event|Event|Hospital Course|6266,6274|false|false|false|||tramadol
Procedure|Laboratory Procedure|Hospital Course|6266,6274|false|false|false|C1266765|Tramadol measurement (procedure)|tramadol
Drug|Biomedical or Dental Material|Hospital Course|6289,6295|false|false|false|C0039225|Tablet Dosage Form|tablet
Event|Event|Hospital Course|6289,6295|false|false|false|||tablet
Finding|Functional Concept|Hospital Course|6299,6307|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|6302,6307|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|6302,6307|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Biomedical or Dental Material|Hospital Course|6339,6345|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|6346,6353|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|6346,6353|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|6362,6372|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Pharmacologic Substance|Hospital Course|6362,6372|false|false|false|C0206460|enoxaparin|Enoxaparin
Event|Event|Hospital Course|6362,6372|false|false|false|||Enoxaparin
Drug|Organic Chemical|Hospital Course|6362,6379|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Pharmacologic Substance|Hospital Course|6362,6379|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Biologically Active Substance|Hospital Course|6373,6379|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|6373,6379|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|6373,6379|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|6373,6379|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|6373,6379|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|6373,6379|false|false|false|C0337443|Sodium measurement|Sodium
Event|Event|Hospital Course|6401,6410|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|6401,6410|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|6401,6410|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|6401,6410|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|6401,6410|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|6401,6422|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|6401,6422|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|6411,6422|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|6411,6422|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|6411,6422|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|Hospital Course|6424,6428|false|false|false|||Home
Finding|Idea or Concept|Hospital Course|6424,6428|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|6424,6428|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|6424,6428|false|false|false|C1553498|home health encounter|Home
Event|Event|Hospital Course|6431,6440|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|6431,6440|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|6431,6440|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|6431,6440|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|6431,6440|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|6431,6450|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|6441,6450|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|6441,6450|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|6441,6450|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|6441,6450|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|6441,6450|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Functional Concept|Hospital Course|6452,6462|false|false|false|C0036525;C1522484|Metastatic to;metastatic qualifier|Metastatic
Disorder|Neoplastic Process|Hospital Course|6452,6477|false|false|false|C0278498|Malignant neoplasm of stomach stage IV|Metastatic gastric cancer
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6463,6470|false|false|false|C0038351|Stomach|gastric
Disorder|Neoplastic Process|Hospital Course|6463,6477|false|false|false|C0024623;C0699791|Malignant neoplasm of stomach;Stomach Carcinoma|gastric cancer
Disorder|Neoplastic Process|Hospital Course|6471,6477|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Hospital Course|6471,6477|false|false|false|||cancer
Attribute|Clinical Attribute|Hospital Course|6479,6484|false|false|false|C1300072|Tumor stage|stage
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6498,6506|false|false|false|C0041967|Urethra|Urethral
Drug|Biomedical or Dental Material|Hospital Course|6498,6506|false|false|false|C2349082|Urethral Dosage Form|Urethral
Finding|Functional Concept|Hospital Course|6498,6506|false|false|false|C1522518|Intraurethral Route of Administration|Urethral
Disorder|Disease or Syndrome|Hospital Course|6498,6516|false|false|false|C0041974|Urethral Stenosis|Urethral stricture
Finding|Pathologic Function|Hospital Course|6498,6516|false|false|false|C4551691|Urethral stricture|Urethral stricture
Event|Event|Hospital Course|6507,6516|false|false|false|||stricture
Finding|Pathologic Function|Hospital Course|6507,6516|false|false|false|C1261287|Stenosis|stricture
Finding|Mental Process|Discharge Condition|6540,6546|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|6540,6553|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|6540,6553|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|6547,6553|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|6547,6553|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|6555,6560|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|6555,6560|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|6565,6573|false|false|false|||coherent
Finding|Finding|Discharge Condition|6565,6573|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|6575,6580|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|6575,6597|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|6575,6597|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|6584,6597|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|6584,6597|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|6584,6597|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|6599,6604|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|6599,6604|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|6599,6604|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|6599,6604|false|false|false|||Alert
Finding|Finding|Discharge Condition|6599,6604|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|6599,6604|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|6599,6604|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|6609,6620|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|6609,6620|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|6622,6630|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|6622,6630|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|6622,6630|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|6631,6637|false|false|false|C5889824||Status
Event|Event|Discharge Condition|6631,6637|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|6631,6637|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|6639,6649|false|false|false|||Ambulatory
Finding|Functional Concept|Discharge Condition|6639,6649|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|6639,6649|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|6639,6649|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|6639,6649|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|6652,6663|false|false|false|||Independent
Finding|Finding|Discharge Condition|6652,6663|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Condition|6652,6663|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Gene or Genome|Discharge Instructions|6692,6696|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|Discharge Instructions|6716,6724|false|false|false|||pleasure
Finding|Intellectual Product|Discharge Instructions|6716,6724|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|Discharge Instructions|6716,6724|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|Discharge Instructions|6732,6736|false|false|false|C1947933|care activity|care
Event|Event|Discharge Instructions|6732,6736|false|false|false|||care
Finding|Finding|Discharge Instructions|6732,6736|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|6732,6736|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|6732,6739|false|false|false|C1555558|care of - AddressPartType|care of
Event|Event|Discharge Instructions|6771,6779|false|false|false|||admitted
Finding|Idea or Concept|Discharge Instructions|6787,6795|false|false|false|C1547192|Organization unit type - Hospital|hospital
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|6801,6808|false|false|false|C0038351|Stomach|gastric
Disorder|Neoplastic Process|Discharge Instructions|6801,6815|false|false|false|C0024623;C0699791|Malignant neoplasm of stomach;Stomach Carcinoma|gastric cancer
Disorder|Neoplastic Process|Discharge Instructions|6809,6815|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Discharge Instructions|6809,6815|false|false|false|||cancer
Event|Event|Discharge Instructions|6828,6837|false|false|false|||attempted
Event|Event|Discharge Instructions|6853,6865|false|false|false|||laparoscopic
Procedure|Diagnostic Procedure|Discharge Instructions|6853,6865|false|false|false|C0031150|Laparoscopy|laparoscopic
Finding|Idea or Concept|Discharge Instructions|6867,6874|false|false|false|C1550516|Target Awareness - partial|partial
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|6867,6886|false|false|false|C0030600|Subtotal gastrectomy|partial gastrectomy
Event|Event|Discharge Instructions|6875,6886|false|false|false|||gastrectomy
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|6875,6886|false|false|false|C0017118|Gastrectomy|gastrectomy
Event|Event|Discharge Instructions|6891,6902|false|false|false|||gastroscopy
Procedure|Diagnostic Procedure|Discharge Instructions|6891,6902|false|false|false|C0017195|Endoscopy of stomach|gastroscopy
Attribute|Clinical Attribute|Discharge Instructions|6919,6932|true|false|false|C0802632||complications
Event|Event|Discharge Instructions|6919,6932|false|false|false|||complications
Finding|Functional Concept|Discharge Instructions|6919,6932|true|false|false|C0009566;C1171258|Complication;complication aspects|complications
Finding|Pathologic Function|Discharge Instructions|6919,6932|true|false|false|C0009566;C1171258|Complication;complication aspects|complications
Event|Event|Discharge Instructions|6938,6947|false|false|false|||tolerated
Attribute|Clinical Attribute|Discharge Instructions|6952,6961|false|false|false|C0945766||procedure
Event|Event|Discharge Instructions|6952,6961|false|false|false|||procedure
Event|Occupational Activity|Discharge Instructions|6952,6961|false|false|false|C1546467|Act Class - procedure|procedure
Finding|Functional Concept|Discharge Instructions|6952,6961|false|false|false|C2700391|Procedure (set of actions)|procedure
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|6952,6961|false|false|false|C0184661|Interventional procedure|procedure
Finding|Finding|Discharge Instructions|6962,6966|false|false|false|C5575035|Well (answer to question)|well
Event|Event|Discharge Instructions|6976,6986|false|false|false|||ambulating
Event|Event|Discharge Instructions|6988,6996|false|false|false|||stooling
Finding|Body Substance|Discharge Instructions|6988,6996|false|false|false|C0015733|Feces|stooling
Event|Event|Discharge Instructions|6998,7008|false|false|false|||tolerating
Finding|Daily or Recreational Activity|Discharge Instructions|7011,7023|false|false|false|C0184625||regular diet
Drug|Food|Discharge Instructions|7019,7023|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|Discharge Instructions|7019,7023|false|false|false|||diet
Finding|Functional Concept|Discharge Instructions|7019,7023|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|Discharge Instructions|7019,7023|false|false|false|C0012159|Diet therapy|diet
Attribute|Clinical Attribute|Discharge Instructions|7034,7038|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|7034,7038|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|7034,7038|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|7034,7038|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Discharge Instructions|7043,7053|false|false|false|||controlled
Attribute|Clinical Attribute|Discharge Instructions|7057,7061|false|false|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|7057,7061|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|7057,7061|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|Discharge Instructions|7062,7073|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|7062,7073|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|7062,7073|false|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|7062,7073|false|false|false|C4284232|Medications|medications
Finding|Functional Concept|Discharge Instructions|7074,7082|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Discharge Instructions|7077,7082|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Discharge Instructions|7077,7082|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Event|Discharge Instructions|7096,7101|false|false|false|||ready
Event|Event|Discharge Instructions|7109,7119|false|false|false|||discharged
Event|Event|Discharge Instructions|7123,7127|false|false|false|||home
Finding|Idea or Concept|Discharge Instructions|7123,7127|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Discharge Instructions|7123,7127|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Discharge Instructions|7123,7127|false|false|false|C1553498|home health encounter|home
Event|Event|Discharge Instructions|7147,7162|false|false|false|||recommendations
Finding|Idea or Concept|Discharge Instructions|7147,7162|false|false|false|C0034866|Recommendation|recommendations
Event|Event|Discharge Instructions|7173,7179|false|false|false|||ensure
Event|Event|Discharge Instructions|7182,7188|false|false|false|||speedy
Finding|Finding|Discharge Instructions|7193,7203|false|false|false|C5453124|Uneventful|uneventful
Event|Activity|Discharge Instructions|7204,7212|false|false|false|C0237820||recovery
Event|Event|Discharge Instructions|7204,7212|false|false|false|||recovery
Finding|Organism Function|Discharge Instructions|7204,7212|false|false|false|C2004454|Recovery - healing process|recovery
Event|Activity|Discharge Instructions|7216,7224|false|false|false|C0441655|Activities|ACTIVITY
Event|Event|Discharge Instructions|7216,7224|false|false|false|||ACTIVITY
Finding|Daily or Recreational Activity|Discharge Instructions|7216,7224|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|ACTIVITY
Finding|Finding|Discharge Instructions|7216,7224|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|ACTIVITY
Event|Event|Discharge Instructions|7235,7240|false|false|false|||drive
Event|Event|Discharge Instructions|7264,7270|false|false|false|||taking
Attribute|Clinical Attribute|Discharge Instructions|7271,7275|false|false|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|7271,7275|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|7271,7275|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Hazardous or Poisonous Substance|Discharge Instructions|7271,7284|false|false|false|C0002771|Analgesics|pain medicine
Drug|Organic Chemical|Discharge Instructions|7271,7284|false|false|false|C0002771|Analgesics|pain medicine
Drug|Pharmacologic Substance|Discharge Instructions|7271,7284|false|false|false|C0002771|Analgesics|pain medicine
Drug|Pharmacologic Substance|Discharge Instructions|7276,7284|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Event|Event|Discharge Instructions|7276,7284|false|false|false|||medicine
Event|Event|Discharge Instructions|7305,7312|false|false|false|||respond
Event|Event|Discharge Instructions|7319,7328|false|false|false|||emergency
Finding|Finding|Discharge Instructions|7319,7328|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Idea or Concept|Discharge Instructions|7319,7328|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Intellectual Product|Discharge Instructions|7319,7328|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Pathologic Function|Discharge Instructions|7319,7328|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Phenomenon|Phenomenon or Process|Discharge Instructions|7319,7328|false|false|false|C0013956|Emergency Situation|emergency
Procedure|Health Care Activity|Discharge Instructions|7319,7328|false|false|false|C1553500|emergency encounter|emergency
Event|Event|Discharge Instructions|7346,7352|false|false|false|||stairs
Finding|Finding|Discharge Instructions|7346,7352|false|false|false|C4300351|Prior functioning.stairs|stairs
Event|Event|Discharge Instructions|7365,7373|false|false|false|||continue
Event|Event|Discharge Instructions|7377,7381|false|false|false|||walk
Event|Event|Discharge Instructions|7382,7389|false|false|false|||several
Disorder|Disease or Syndrome|Discharge Instructions|7391,7396|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Event|Event|Discharge Instructions|7391,7396|false|false|false|||times
Finding|Idea or Concept|Discharge Instructions|7399,7402|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Discharge Instructions|7399,7402|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Discharge Instructions|7431,7436|false|false|false|||avoid
Event|Event|Discharge Instructions|7437,7446|false|false|false|||traveling
Event|Event|Discharge Instructions|7452,7461|false|false|false|||distances
Event|Event|Discharge Instructions|7473,7476|false|false|false|||see
Attribute|Clinical Attribute|Discharge Instructions|7482,7489|false|false|false|C5444295||surgeon
Finding|Idea or Concept|Discharge Instructions|7498,7502|false|false|false|C1552851|next - HtmlLinkType|next
Event|Event|Discharge Instructions|7503,7508|false|false|false|||visit
Finding|Social Behavior|Discharge Instructions|7503,7508|false|false|false|C0545082|Visit|visit
Event|Event|Discharge Instructions|7521,7526|false|false|false|||start
Drug|Amino Acid, Peptide, or Protein|Discharge Instructions|7532,7537|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|Discharge Instructions|7532,7537|false|false|false|C1570446|TNFSF14 protein, human|light
Finding|Finding|Discharge Instructions|7532,7537|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|Discharge Instructions|7532,7537|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|Discharge Instructions|7532,7537|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|Discharge Instructions|7532,7537|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|7532,7537|false|false|false|C0031765|Phototherapy|light
Finding|Daily or Recreational Activity|Discharge Instructions|7532,7546|false|false|false|C1517883|Light Exercise|light exercise
Event|Event|Discharge Instructions|7538,7546|false|false|false|||exercise
Finding|Daily or Recreational Activity|Discharge Instructions|7538,7546|false|false|false|C0015259|Exercise|exercise
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|7538,7546|false|false|false|C1522704|Exercise Pain Management|exercise
Event|Event|Discharge Instructions|7561,7572|false|false|false|||comfortable
Finding|Finding|Discharge Instructions|7561,7572|false|false|false|C5546696|Feeling comfortable|comfortable
Event|Event|Discharge Instructions|7582,7590|false|false|false|||increase
Event|Activity|Discharge Instructions|7596,7604|false|false|false|C0441655|Activities|activity
Event|Event|Discharge Instructions|7596,7604|false|false|false|||activity
Finding|Daily or Recreational Activity|Discharge Instructions|7596,7604|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Finding|Finding|Discharge Instructions|7596,7604|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Event|Event|Discharge Instructions|7605,7609|false|false|false|||back
Drug|Biomedical or Dental Material|Discharge Instructions|7618,7626|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|Discharge Instructions|7618,7626|false|false|false|||baseline
Finding|Idea or Concept|Discharge Instructions|7618,7626|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|Discharge Instructions|7631,7640|false|false|false|||tolerated
Event|Event|Discharge Instructions|7650,7658|false|false|false|||exercise
Finding|Daily or Recreational Activity|Discharge Instructions|7650,7658|false|false|false|C0015259|Exercise|exercise
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|7650,7658|false|false|false|C1522704|Exercise Pain Management|exercise
Event|Event|Discharge Instructions|7666,7673|false|false|false|||started
Event|Event|Discharge Instructions|7693,7696|false|false|false|||use
Event|Event|Discharge Instructions|7697,7703|false|false|false|||common
Finding|Functional Concept|Discharge Instructions|7697,7703|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Finding|Intellectual Product|Discharge Instructions|7697,7703|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Event|Event|Discharge Instructions|7705,7710|false|false|false|||sense
Finding|Organ or Tissue Function|Discharge Instructions|7705,7710|false|false|false|C0036658|Sensory perception|sense
Event|Event|Discharge Instructions|7715,7717|false|false|false|||go
Event|Activity|Discharge Instructions|7747,7754|true|false|false|C0206244|Lifting|lifting
Event|Event|Discharge Instructions|7747,7754|false|false|false|||lifting
Finding|Finding|Discharge Instructions|7756,7765|true|false|false|C3845310|10 pounds|10 pounds
Event|Event|Discharge Instructions|7781,7788|false|false|false|||cleared
Attribute|Clinical Attribute|Discharge Instructions|7798,7805|false|false|false|C5444295||surgeon
Finding|Finding|Discharge Instructions|7807,7814|false|false|false|C3888388|Usually|usually
Event|Event|Discharge Instructions|7841,7847|false|false|false|||resume
Finding|Behavior|Discharge Instructions|7848,7854|false|false|false|C0036864|Sex Behavior|sexual
Finding|Behavior|Discharge Instructions|7848,7863|false|false|false|C0036864;C5575036|Sex Behavior;Sexual Activity|sexual activity
Finding|Individual Behavior|Discharge Instructions|7848,7863|false|false|false|C0036864;C5575036|Sex Behavior;Sexual Activity|sexual activity
Event|Activity|Discharge Instructions|7855,7863|false|false|false|C0441655|Activities|activity
Event|Event|Discharge Instructions|7855,7863|false|false|false|||activity
Finding|Daily or Recreational Activity|Discharge Instructions|7855,7863|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Finding|Finding|Discharge Instructions|7855,7863|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Event|Event|Discharge Instructions|7876,7882|false|false|false|||doctor
Finding|Intellectual Product|Discharge Instructions|7876,7882|false|false|false|C2348314|Doctor - Title|doctor
Event|Event|Discharge Instructions|7921,7925|false|false|false|||FEEL
Finding|Mental Process|Discharge Instructions|7921,7925|false|false|false|C1527305|Feelings|FEEL
Event|Event|Discharge Instructions|7938,7942|false|false|false|||feel
Finding|Intellectual Product|Discharge Instructions|7938,7947|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|feel weak
Finding|Sign or Symptom|Discharge Instructions|7938,7947|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|feel weak
Event|Event|Discharge Instructions|7943,7947|false|false|false|||weak
Finding|Intellectual Product|Discharge Instructions|7943,7947|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|weak
Finding|Sign or Symptom|Discharge Instructions|7943,7947|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|weak
Event|Event|Discharge Instructions|7952,7958|false|false|false|||washed
Event|Event|Discharge Instructions|7987,7991|false|false|false|||want
Drug|Indicator, Reagent, or Diagnostic Aid|Discharge Instructions|7996,7999|false|false|false|C4283878|Neutrophil Activation Probe Imaging Agent|nap
Event|Event|Discharge Instructions|7996,7999|false|false|false|||nap
Finding|Gene or Genome|Discharge Instructions|7996,7999|false|false|false|C0870935;C1423800|CTNNBL1 gene;Napping|nap
Finding|Physiologic Function|Discharge Instructions|7996,7999|false|false|false|C0870935;C1423800|CTNNBL1 gene;Napping|nap
Finding|Intellectual Product|Discharge Instructions|8000,8005|false|false|false|C4050225|Often - answer to question|often
Finding|Gene or Genome|Discharge Instructions|8007,8013|false|false|false|C1424587|LITAF gene|Simple
Drug|Hazardous or Poisonous Substance|Discharge Instructions|8024,8031|false|false|false|C0178629|exhaust|exhaust
Finding|Sign or Symptom|Discharge Instructions|8054,8058|false|false|false|C0234233;C1442877|Sore skin;Sore to touch|sore
Disorder|Disease or Syndrome|Discharge Instructions|8054,8065|false|false|false|C0031350|Pharyngitis|sore throat
Drug|Organic Chemical|Discharge Instructions|8054,8065|false|false|false|C0723402;C3244654|Sore Throat brand of Phenol;Sore Throat brand of benzocaine & menthol|sore throat
Drug|Pharmacologic Substance|Discharge Instructions|8054,8065|false|false|false|C0723402;C3244654|Sore Throat brand of Phenol;Sore Throat brand of benzocaine & menthol|sore throat
Finding|Sign or Symptom|Discharge Instructions|8054,8065|false|false|false|C0242429|Sore Throat|sore throat
Anatomy|Body Location or Region|Discharge Instructions|8059,8065|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|8059,8065|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Drug|Pharmacologic Substance|Discharge Instructions|8059,8065|false|false|false|C1950455|Throat Homeopathic Medication|throat
Event|Event|Discharge Instructions|8059,8065|false|false|false|||throat
Finding|Body Substance|Discharge Instructions|8059,8065|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Finding|Intellectual Product|Discharge Instructions|8059,8065|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Event|Event|Discharge Instructions|8079,8083|false|false|false|||tube
Finding|Functional Concept|Discharge Instructions|8079,8083|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Finding|Gene or Genome|Discharge Instructions|8079,8083|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Anatomy|Body Location or Region|Discharge Instructions|8102,8108|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|8102,8108|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Drug|Pharmacologic Substance|Discharge Instructions|8102,8108|false|false|false|C1950455|Throat Homeopathic Medication|throat
Event|Event|Discharge Instructions|8102,8108|false|false|false|||throat
Finding|Body Substance|Discharge Instructions|8102,8108|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Finding|Intellectual Product|Discharge Instructions|8102,8108|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Event|Event|Discharge Instructions|8120,8127|false|false|false|||surgery
Finding|Finding|Discharge Instructions|8120,8127|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Discharge Instructions|8120,8127|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Discharge Instructions|8120,8127|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|8120,8127|false|false|false|C0543467|Operative Surgical Procedures|surgery
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|8135,8141|false|false|false|C0021853|Intestines|BOWELS
Event|Event|Discharge Instructions|8145,8157|false|false|false|||Constipation
Finding|Sign or Symptom|Discharge Instructions|8145,8157|false|false|false|C0009806|Constipation|Constipation
Finding|Functional Concept|Discharge Instructions|8163,8169|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Finding|Intellectual Product|Discharge Instructions|8163,8169|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Finding|Pathologic Function|Discharge Instructions|8170,8181|false|false|false|C0879626|Adverse effects|side effect
Event|Event|Discharge Instructions|8175,8181|false|false|false|||effect
Drug|Hazardous or Poisonous Substance|Discharge Instructions|8185,8193|false|false|false|C0027415|Narcotics|narcotic
Drug|Pharmacologic Substance|Discharge Instructions|8185,8193|false|false|false|C0027415|Narcotics|narcotic
Event|Event|Discharge Instructions|8185,8193|false|false|false|||narcotic
Attribute|Clinical Attribute|Discharge Instructions|8194,8198|false|false|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|8194,8198|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|8194,8198|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Hazardous or Poisonous Substance|Discharge Instructions|8194,8207|false|false|false|C0002771|Analgesics|pain medicine
Drug|Organic Chemical|Discharge Instructions|8194,8207|false|false|false|C0002771|Analgesics|pain medicine
Drug|Pharmacologic Substance|Discharge Instructions|8194,8207|false|false|false|C0002771|Analgesics|pain medicine
Drug|Pharmacologic Substance|Discharge Instructions|8199,8207|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Event|Event|Discharge Instructions|8199,8207|false|false|false|||medicine
Drug|Organic Chemical|Discharge Instructions|8217,8226|false|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|Discharge Instructions|8217,8226|false|false|false|C0030049|oxycodone|oxycodone
Event|Event|Discharge Instructions|8217,8226|false|false|false|||oxycodone
Procedure|Laboratory Procedure|Discharge Instructions|8217,8226|false|false|false|C0524222|Oxycodone measurement|oxycodone
Event|Event|Discharge Instructions|8231,8237|false|false|false|||needed
Event|Event|Discharge Instructions|8247,8251|false|false|false|||take
Finding|Body Substance|Discharge Instructions|8254,8259|false|false|false|C0015733|Feces|stool
Drug|Organic Chemical|Discharge Instructions|8254,8268|false|false|false|C0301470;C1154263|Stool Softener;Stool Softener brand of docusate sodium|stool softener
Drug|Pharmacologic Substance|Discharge Instructions|8254,8268|false|false|false|C0301470;C1154263|Stool Softener;Stool Softener brand of docusate sodium|stool softener
Event|Event|Discharge Instructions|8260,8268|false|false|false|||softener
Drug|Organic Chemical|Discharge Instructions|8279,8285|false|false|false|C0282139|Colace|Colace
Drug|Pharmacologic Substance|Discharge Instructions|8279,8285|false|false|false|C0282139|Colace|Colace
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|8291,8298|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|Discharge Instructions|8291,8298|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|Discharge Instructions|8291,8298|false|false|false|C0006935|capsule (pharmacologic)|capsule
Drug|Organic Chemical|Discharge Instructions|8303,8309|false|false|false|C0720654|Gentle|gentle
Drug|Pharmacologic Substance|Discharge Instructions|8303,8309|false|false|false|C0720654|Gentle|gentle
Drug|Organic Chemical|Discharge Instructions|8303,8318|false|false|false|C0720655|Gentle Laxative|gentle laxative
Drug|Pharmacologic Substance|Discharge Instructions|8303,8318|false|false|false|C0720655|Gentle Laxative|gentle laxative
Drug|Pharmacologic Substance|Discharge Instructions|8310,8318|false|false|false|C0282090|Laxatives|laxative
Event|Event|Discharge Instructions|8310,8318|false|false|false|||laxative
Drug|Food|Discharge Instructions|8328,8332|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|milk
Drug|Immunologic Factor|Discharge Instructions|8328,8332|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|milk
Drug|Pharmacologic Substance|Discharge Instructions|8328,8332|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|milk
Drug|Substance|Discharge Instructions|8328,8332|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|milk
Event|Event|Discharge Instructions|8328,8332|false|false|false|||milk
Finding|Body Substance|Discharge Instructions|8328,8332|false|false|false|C0026131;C1546713|Milk (body substance);Milk Specimen Code|milk
Finding|Intellectual Product|Discharge Instructions|8328,8332|false|false|false|C0026131;C1546713|Milk (body substance);Milk Specimen Code|milk
Drug|Inorganic Chemical|Discharge Instructions|8337,8345|false|false|false|C0024477|magnesium oxide|magnesia
Drug|Pharmacologic Substance|Discharge Instructions|8337,8345|false|false|false|C0024477|magnesium oxide|magnesia
Event|Event|Discharge Instructions|8337,8345|false|false|false|||magnesia
Disorder|Disease or Syndrome|Discharge Instructions|8349,8352|false|false|false|C0265246|Townes syndrome|tbs
Event|Event|Discharge Instructions|8349,8352|false|false|false|||tbs
Finding|Finding|Discharge Instructions|8349,8352|false|false|false|C1419808;C5780809;C5958753|SALL1 gene;SALL1 wt Allele;Toxicity Burden Score|tbs
Finding|Gene or Genome|Discharge Instructions|8349,8352|false|false|false|C1419808;C5780809;C5958753|SALL1 gene;SALL1 wt Allele;Toxicity Burden Score|tbs
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|8349,8352|false|false|false|C5889868|theta-burst stimulation|tbs
Finding|Idea or Concept|Discharge Instructions|8362,8365|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Discharge Instructions|8362,8365|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Discharge Instructions|8379,8383|false|false|false|||both
Drug|Pharmacologic Substance|Discharge Instructions|8394,8403|false|false|false|C0013227|Pharmaceutical Preparations|medicines
Event|Event|Discharge Instructions|8394,8403|false|false|false|||medicines
Attribute|Clinical Attribute|Discharge Instructions|8414,8426|true|false|false|C5886759|Prescription (attribute)|prescription
Event|Event|Discharge Instructions|8414,8426|false|false|false|||prescription
Finding|Intellectual Product|Discharge Instructions|8414,8426|true|false|false|C1521941|prescription document|prescription
Procedure|Health Care Activity|Discharge Instructions|8414,8426|true|false|false|C0033080|Prescription (procedure)|prescription
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|8459,8464|false|false|false|C0021853|Intestines|bowel
Finding|Organism Function|Discharge Instructions|8459,8473|true|false|false|C0011135|Defecation|bowel movement
Event|Event|Discharge Instructions|8465,8473|false|false|false|||movement
Finding|Organism Function|Discharge Instructions|8465,8473|true|false|false|C0026649|Movement|movement
Finding|Intellectual Product|Discharge Instructions|8478,8487|false|false|false|C2984058|Have Pain|have pain
Attribute|Clinical Attribute|Discharge Instructions|8483,8487|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|8483,8487|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|8483,8487|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|8483,8487|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Discharge Instructions|8489,8495|false|false|false|||moving
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|8500,8506|false|false|false|C0021853|Intestines|bowels
Event|Event|Discharge Instructions|8508,8512|false|false|false|||call
Attribute|Clinical Attribute|Discharge Instructions|8518,8525|false|false|false|C5444295||surgeon
Event|Activity|Discharge Instructions|8540,8550|false|false|false|C3241922|Operation Activity|operations
Event|Event|Discharge Instructions|8540,8550|false|false|false|||operations
Finding|Functional Concept|Discharge Instructions|8540,8550|false|false|false|C0038895;C3244305;C3244306|ActInformationPrivacyReason - operations;HL7PublishingSubSection - operations;Surgical aspects|operations
Finding|Intellectual Product|Discharge Instructions|8540,8550|false|false|false|C0038895;C3244305;C3244306|ActInformationPrivacyReason - operations;HL7PublishingSubSection - operations;Surgical aspects|operations
Event|Event|Discharge Instructions|8552,8560|false|false|false|||diarrhea
Finding|Finding|Discharge Instructions|8552,8560|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|Discharge Instructions|8552,8560|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Event|Event|Discharge Instructions|8565,8570|false|false|false|||occur
Event|Event|Discharge Instructions|8584,8592|false|false|false|||diarrhea
Finding|Finding|Discharge Instructions|8584,8592|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|Discharge Instructions|8584,8592|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Drug|Organic Chemical|Discharge Instructions|8605,8618|false|false|false|C0718564|Anti-Diarrhea|anti-diarrhea
Drug|Pharmacologic Substance|Discharge Instructions|8605,8618|false|false|false|C0718564|Anti-Diarrhea|anti-diarrhea
Drug|Pharmacologic Substance|Discharge Instructions|8619,8628|false|false|false|C0013227|Pharmaceutical Preparations|medicines
Event|Event|Discharge Instructions|8619,8628|false|false|false|||medicines
Drug|Substance|Discharge Instructions|8647,8653|false|false|false|C0302908|Liquid substance|fluids
Event|Event|Discharge Instructions|8647,8653|false|false|false|||fluids
Finding|Body Substance|Discharge Instructions|8647,8653|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|8647,8653|false|false|false|C0016286|Fluid Therapy|fluids
Event|Event|Discharge Instructions|8658,8661|false|false|false|||see
Event|Event|Discharge Instructions|8668,8672|false|false|false|||goes
Event|Event|Discharge Instructions|8694,8696|false|false|false|||go
Event|Event|Discharge Instructions|8710,8716|false|false|false|||severe
Finding|Finding|Discharge Instructions|8710,8716|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Discharge Instructions|8710,8716|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Discharge Instructions|8725,8733|false|false|false|C0231218;C0557911;C2987492|Feel Ill Question;Feeling bad emotionally;Malaise|feel ill
Finding|Sign or Symptom|Discharge Instructions|8725,8733|false|false|false|C0231218;C0557911;C2987492|Feel Ill Question;Feeling bad emotionally;Malaise|feel ill
Finding|Sign or Symptom|Discharge Instructions|8730,8733|false|false|false|C0231218|Malaise|ill
Event|Event|Discharge Instructions|8742,8746|false|false|false|||call
Attribute|Clinical Attribute|Discharge Instructions|8752,8759|false|false|false|C5444295||surgeon
Attribute|Clinical Attribute|Discharge Instructions|8762,8766|false|false|false|C2598155||PAIN
Event|Event|Discharge Instructions|8762,8766|false|false|false|||PAIN
Finding|Functional Concept|Discharge Instructions|8762,8766|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|PAIN
Finding|Sign or Symptom|Discharge Instructions|8762,8766|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|PAIN
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|8762,8777|false|false|false|C0002766|Pain management (procedure)|PAIN MANAGEMENT
Event|Event|Discharge Instructions|8767,8777|false|false|false|||MANAGEMENT
Event|Occupational Activity|Discharge Instructions|8767,8777|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|MANAGEMENT
Procedure|Health Care Activity|Discharge Instructions|8767,8777|false|false|false|C0376636|Disease Management|MANAGEMENT
Event|Event|Discharge Instructions|8795,8805|false|false|false|||discharged
Attribute|Clinical Attribute|Discharge Instructions|8813,8825|false|false|false|C5886759|Prescription (attribute)|prescription
Event|Event|Discharge Instructions|8813,8825|false|false|false|||prescription
Finding|Intellectual Product|Discharge Instructions|8813,8825|false|false|false|C1521941|prescription document|prescription
Procedure|Health Care Activity|Discharge Instructions|8813,8825|false|false|false|C0033080|Prescription (procedure)|prescription
Drug|Organic Chemical|Discharge Instructions|8832,8841|false|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|Discharge Instructions|8832,8841|false|false|false|C0030049|oxycodone|oxycodone
Event|Event|Discharge Instructions|8832,8841|false|false|false|||oxycodone
Procedure|Laboratory Procedure|Discharge Instructions|8832,8841|false|false|false|C0524222|Oxycodone measurement|oxycodone
Attribute|Clinical Attribute|Discharge Instructions|8847,8851|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|8847,8851|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|8847,8851|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|8847,8851|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Discharge Instructions|8847,8859|false|false|false|C5548091|Demonstrates adequate pain control|pain control
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|8847,8859|false|false|false|C0002766;C1304888|Pain control;Pain management (procedure)|pain control
Drug|Organic Chemical|Discharge Instructions|8852,8859|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|Discharge Instructions|8852,8859|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|Discharge Instructions|8852,8859|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Event|Event|Discharge Instructions|8852,8859|false|false|false|||control
Finding|Conceptual Entity|Discharge Instructions|8852,8859|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|Discharge Instructions|8852,8859|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|Discharge Instructions|8852,8859|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Event|Event|Discharge Instructions|8869,8873|false|false|false|||take
Drug|Organic Chemical|Discharge Instructions|8874,8881|false|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|Discharge Instructions|8874,8881|false|false|false|C0699142|Tylenol|Tylenol
Event|Event|Discharge Instructions|8874,8881|false|false|false|||Tylenol
Event|Event|Discharge Instructions|8885,8893|false|false|false|||directed
Event|Event|Discharge Instructions|8910,8916|false|false|false|||3500mg
Event|Event|Discharge Instructions|8930,8934|false|false|false|||Take
Event|Event|Discharge Instructions|8967,8974|false|false|false|||surgery
Finding|Finding|Discharge Instructions|8967,8974|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Discharge Instructions|8967,8974|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Discharge Instructions|8967,8974|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|8967,8974|false|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Event|Discharge Instructions|8987,8991|false|false|false|||skip
Event|Event|Discharge Instructions|8994,8998|false|false|false|||dose
Event|Event|Discharge Instructions|9002,9010|false|false|false|||increase
Finding|Functional Concept|Discharge Instructions|9002,9010|false|true|false|C0442805|Increase|increase
Finding|Finding|Discharge Instructions|9011,9015|false|true|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Discharge Instructions|9011,9015|false|true|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Discharge Instructions|9011,9015|false|true|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|Discharge Instructions|9024,9029|false|false|false|||doses
Attribute|Clinical Attribute|Discharge Instructions|9053,9057|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|9053,9057|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|9053,9057|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|9053,9057|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Discharge Instructions|9078,9082|false|false|false|||need
Event|Event|Discharge Instructions|9096,9100|false|false|false|||take
Drug|Organic Chemical|Discharge Instructions|9105,9114|false|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|Discharge Instructions|9105,9114|false|false|false|C0030049|oxycodone|oxycodone
Event|Event|Discharge Instructions|9105,9114|false|false|false|||oxycodone
Procedure|Laboratory Procedure|Discharge Instructions|9105,9114|false|false|false|C0524222|Oxycodone measurement|oxycodone
Event|Event|Discharge Instructions|9119,9127|false|false|false|||moderate
Finding|Finding|Discharge Instructions|9119,9127|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|Discharge Instructions|9119,9127|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Finding|Discharge Instructions|9132,9138|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Discharge Instructions|9132,9138|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Finding|Discharge Instructions|9132,9143|false|false|false|C0278140;C4050465;C4521229|Neck Pain Score 6;Severe Extremity Pain;Severe pain|severe pain
Attribute|Clinical Attribute|Discharge Instructions|9139,9143|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|9139,9143|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|9139,9143|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|9139,9143|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Discharge Instructions|9148,9158|false|false|false|||controlled
Drug|Organic Chemical|Discharge Instructions|9167,9174|false|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|Discharge Instructions|9167,9174|false|false|false|C0699142|Tylenol|Tylenol
Event|Event|Discharge Instructions|9184,9188|false|false|false|||take
Finding|Body Substance|Discharge Instructions|9191,9196|false|false|false|C0015733|Feces|stool
Drug|Organic Chemical|Discharge Instructions|9191,9205|false|false|false|C0301470;C1154263|Stool Softener;Stool Softener brand of docusate sodium|stool softener
Drug|Pharmacologic Substance|Discharge Instructions|9191,9205|false|false|false|C0301470;C1154263|Stool Softener;Stool Softener brand of docusate sodium|stool softener
Event|Event|Discharge Instructions|9197,9205|false|false|false|||softener
Drug|Hazardous or Poisonous Substance|Discharge Instructions|9215,9224|false|false|false|C0027415|Narcotics|narcotics
Drug|Pharmacologic Substance|Discharge Instructions|9215,9224|false|false|false|C0027415|Narcotics|narcotics
Event|Event|Discharge Instructions|9215,9224|false|false|false|||narcotics
Event|Event|Discharge Instructions|9229,9233|false|false|false|||help
Event|Event|Discharge Instructions|9234,9241|false|false|false|||prevent
Event|Event|Discharge Instructions|9246,9258|false|false|false|||constipation
Finding|Sign or Symptom|Discharge Instructions|9246,9258|false|false|false|C0009806|Constipation|constipation
Event|Event|Discharge Instructions|9273,9278|false|false|false|||cause
Event|Event|Discharge Instructions|9288,9292|false|false|false|||wean
Attribute|Clinical Attribute|Discharge Instructions|9303,9314|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|9303,9314|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|9303,9314|false|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|9303,9314|false|false|false|C4284232|Medications|medications
Event|Event|Discharge Instructions|9318,9327|false|false|false|||tolerated
Attribute|Clinical Attribute|Discharge Instructions|9337,9341|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|9337,9341|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|9337,9341|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|9337,9341|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Discharge Instructions|9353,9359|false|false|false|||better
Finding|Idea or Concept|Discharge Instructions|9353,9359|false|false|false|C1550462|Observation Interpretation - better|better
Finding|Idea or Concept|Discharge Instructions|9360,9363|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Discharge Instructions|9360,9363|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Idea or Concept|Discharge Instructions|9367,9370|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Discharge Instructions|9367,9370|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Discharge Instructions|9379,9383|false|false|false|||find
Attribute|Clinical Attribute|Discharge Instructions|9388,9392|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|9388,9392|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|9388,9392|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|9388,9392|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Discharge Instructions|9405,9410|false|false|false|||worse
Finding|Finding|Discharge Instructions|9405,9410|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Idea or Concept|Discharge Instructions|9405,9410|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Idea or Concept|Discharge Instructions|9422,9428|false|false|false|C1550462|Observation Interpretation - better|better
Event|Event|Discharge Instructions|9437,9444|false|false|false|||contact
Attribute|Clinical Attribute|Discharge Instructions|9450,9457|false|false|false|C5444295||surgeon
Event|Event|Discharge Instructions|9467,9477|false|false|false|||experience
Event|Event|Discharge Instructions|9507,9514|false|false|false|||contact
Attribute|Clinical Attribute|Discharge Instructions|9521,9528|false|false|false|C5444295||surgeon
Finding|Finding|Discharge Instructions|9533,9538|false|false|false|C1444775;C1539835;C3890003|SPEN gene;SPEN wt Allele;Sharp sensation quality|sharp
Finding|Gene or Genome|Discharge Instructions|9533,9538|false|false|false|C1444775;C1539835;C3890003|SPEN gene;SPEN wt Allele;Sharp sensation quality|sharp
Finding|Sign or Symptom|Discharge Instructions|9533,9543|false|false|false|C0455270|Sharp pain|sharp pain
Attribute|Clinical Attribute|Discharge Instructions|9539,9543|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|9539,9543|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|9539,9543|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|9539,9543|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Discharge Instructions|9551,9557|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Discharge Instructions|9551,9557|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Finding|Discharge Instructions|9551,9562|false|false|false|C0278140;C4050465;C4521229|Neck Pain Score 6;Severe Extremity Pain;Severe pain|severe pain
Attribute|Clinical Attribute|Discharge Instructions|9558,9562|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|9558,9562|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|9558,9562|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|9558,9562|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Discharge Instructions|9568,9573|false|false|false|||lasts
Event|Event|Discharge Instructions|9582,9587|false|false|false|||hours
Anatomy|Body Location or Region|Discharge Instructions|9590,9595|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Discharge Instructions|9590,9595|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Discharge Instructions|9590,9600|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Discharge Instructions|9590,9600|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Discharge Instructions|9596,9600|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|9596,9600|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|9596,9600|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|9596,9600|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Discharge Instructions|9602,9610|false|false|false|||pressure
Finding|Finding|Discharge Instructions|9602,9610|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|Discharge Instructions|9602,9610|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|Discharge Instructions|9602,9610|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|Discharge Instructions|9602,9610|false|false|false|C0033095||pressure
Event|Event|Discharge Instructions|9612,9621|false|false|false|||squeezing
Event|Event|Discharge Instructions|9626,9635|false|false|false|||tightness
Drug|Organic Chemical|Discharge Instructions|9638,9643|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|Discharge Instructions|9638,9643|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|Discharge Instructions|9638,9643|false|false|false|||cough
Finding|Sign or Symptom|Discharge Instructions|9638,9643|false|false|false|C0010200|Coughing|cough
Event|Event|Discharge Instructions|9645,9654|false|false|false|||shortness
Attribute|Clinical Attribute|Discharge Instructions|9645,9664|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|Discharge Instructions|9645,9664|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|Discharge Instructions|9658,9664|false|false|false|C0225386|Breath|breath
Event|Event|Discharge Instructions|9666,9674|false|false|false|||wheezing
Finding|Sign or Symptom|Discharge Instructions|9666,9674|false|false|false|C0043144|Wheezing|wheezing
Attribute|Clinical Attribute|Discharge Instructions|9677,9681|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|9677,9681|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|9677,9681|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|9677,9681|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Discharge Instructions|9698,9703|false|false|false|||worse
Finding|Finding|Discharge Instructions|9698,9703|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Idea or Concept|Discharge Instructions|9698,9703|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Finding|Discharge Instructions|9709,9713|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Discharge Instructions|9709,9713|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Discharge Instructions|9709,9713|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Attribute|Clinical Attribute|Discharge Instructions|9717,9721|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|9717,9721|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|9717,9721|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|9717,9721|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Discharge Instructions|9727,9732|false|false|false|||fever
Finding|Finding|Discharge Instructions|9727,9732|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|Discharge Instructions|9727,9732|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|Discharge Instructions|9743,9749|false|false|false|||chills
Finding|Sign or Symptom|Discharge Instructions|9743,9749|false|false|false|C0085593|Chills|chills
Event|Event|Discharge Instructions|9751,9756|false|false|false|||fever
Finding|Finding|Discharge Instructions|9751,9756|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|Discharge Instructions|9751,9756|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|Discharge Instructions|9786,9792|false|false|false|||change
Finding|Functional Concept|Discharge Instructions|9786,9792|false|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|9786,9792|false|false|false|C4319952|Change - procedure|change
Finding|Functional Concept|Discharge Instructions|9786,9795|false|false|false|C0392747|Changing|change in
Event|Event|Discharge Instructions|9796,9802|false|false|false|||nature
Finding|Functional Concept|Discharge Instructions|9796,9802|false|false|false|C0349590;C1262865|Nature;Natures|nature
Finding|Idea or Concept|Discharge Instructions|9796,9802|false|false|false|C0349590;C1262865|Nature;Natures|nature
Event|Event|Discharge Instructions|9806,9813|false|false|false|||quality
Attribute|Clinical Attribute|Discharge Instructions|9822,9826|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|9822,9826|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|9822,9826|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|9822,9826|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|Discharge Instructions|9829,9835|false|false|false|C4255480||nausea
Event|Event|Discharge Instructions|9829,9835|false|false|false|||nausea
Finding|Sign or Symptom|Discharge Instructions|9829,9835|false|false|false|C0027497|Nausea|nausea
Finding|Sign or Symptom|Discharge Instructions|9829,9848|false|false|false|C0027498|Nausea and vomiting|nausea and vomiting
Event|Event|Discharge Instructions|9840,9848|false|false|false|||vomiting
Finding|Sign or Symptom|Discharge Instructions|9840,9848|false|false|false|C0042963|Vomiting|vomiting
Event|Event|Discharge Instructions|9850,9859|false|false|false|||inability
Drug|Substance|Discharge Instructions|9872,9878|false|false|false|C0302908|Liquid substance|fluids
Event|Event|Discharge Instructions|9872,9878|false|false|false|||fluids
Finding|Body Substance|Discharge Instructions|9872,9878|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|9872,9878|false|false|false|C0016286|Fluid Therapy|fluids
Drug|Food|Discharge Instructions|9880,9884|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Drug|Immunologic Factor|Discharge Instructions|9880,9884|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Drug|Pharmacologic Substance|Discharge Instructions|9880,9884|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Event|Event|Discharge Instructions|9880,9884|false|false|false|||food
Attribute|Clinical Attribute|Discharge Instructions|9895,9906|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|9895,9906|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|9895,9906|false|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|9895,9906|false|false|false|C4284232|Medications|medications
Disorder|Disease or Syndrome|Discharge Instructions|9928,9938|false|false|false|C0011175|Dehydration|dehydrated
Event|Event|Discharge Instructions|9928,9938|false|false|false|||dehydrated
Disorder|Disease or Syndrome|Discharge Instructions|9940,9949|false|false|false|C0043352|Xerostomia|dry mouth
Anatomy|Body Location or Region|Discharge Instructions|9944,9949|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Discharge Instructions|9944,9949|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Finding|Discharge Instructions|9951,9967|false|false|false|C0039231|Tachycardia|rapid heart beat
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|9957,9962|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|9957,9962|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Discharge Instructions|9957,9962|false|false|false|C0795691|HEART PROBLEM|heart
Finding|Organ or Tissue Function|Discharge Instructions|9957,9967|false|false|false|C0425583|Heart beat|heart beat
Event|Event|Discharge Instructions|9963,9967|false|false|false|||beat
Event|Event|Discharge Instructions|9970,9977|false|false|false|||feeling
Finding|Sign or Symptom|Discharge Instructions|9970,9983|false|false|false|C0849959|feeling dizzy|feeling dizzy
Finding|Sign or Symptom|Discharge Instructions|9978,9983|false|false|false|C0012833|Dizziness|dizzy
Event|Event|Discharge Instructions|9987,9992|false|false|false|||faint
Finding|Finding|Discharge Instructions|9987,9992|false|false|false|C0039070;C4554554|Faint - appearance;Syncope|faint
Finding|Sign or Symptom|Discharge Instructions|9987,9992|false|false|false|C0039070;C4554554|Faint - appearance;Syncope|faint
Event|Event|Discharge Instructions|10025,10031|false|false|false|||change
Finding|Functional Concept|Discharge Instructions|10025,10031|false|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10025,10031|false|false|false|C4319952|Change - procedure|change
Finding|Functional Concept|Discharge Instructions|10025,10034|false|false|false|C0392747|Changing|change in
Event|Event|Discharge Instructions|10040,10048|false|false|false|||symptoms
Finding|Functional Concept|Discharge Instructions|10040,10048|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Discharge Instructions|10040,10048|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|Discharge Instructions|10056,10064|false|false|false|||symptoms
Finding|Functional Concept|Discharge Instructions|10056,10064|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Discharge Instructions|10056,10064|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|Discharge Instructions|10070,10077|false|false|false|||concern
Finding|Functional Concept|Discharge Instructions|10083,10093|false|false|false|C1524062|Additional|Additional
Attribute|Clinical Attribute|Discharge Instructions|10099,10103|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|10099,10103|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|10099,10103|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|10099,10103|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Discharge Instructions|10120,10125|false|false|false|||worse
Finding|Finding|Discharge Instructions|10120,10125|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Idea or Concept|Discharge Instructions|10120,10125|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Finding|Discharge Instructions|10131,10135|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Discharge Instructions|10131,10135|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Discharge Instructions|10131,10135|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|Discharge Instructions|10140,10145|false|false|false|||going
Anatomy|Body Location or Region|Discharge Instructions|10154,10159|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Discharge Instructions|10154,10159|false|false|false|C0741025|Chest problem|chest
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|10172,10179|false|false|false|C0042027|Urinary tract|urinary
Event|Event|Discharge Instructions|10182,10189|false|false|false|||burning
Finding|Sign or Symptom|Discharge Instructions|10182,10189|false|false|false|C0085624|Burning sensation|burning
Disorder|Disease or Syndrome|Discharge Instructions|10193,10198|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Discharge Instructions|10193,10198|false|false|false|||blood
Finding|Body Substance|Discharge Instructions|10193,10198|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Event|Discharge Instructions|10207,10212|false|false|false|||urine
Finding|Body Substance|Discharge Instructions|10207,10212|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|Discharge Instructions|10207,10212|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|Discharge Instructions|10207,10212|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Event|Event|Medications|10258,10262|false|false|false|||Take
Drug|Pharmacologic Substance|Medications|10271,10280|false|false|false|C0013227|Pharmaceutical Preparations|medicines
Event|Event|Medications|10271,10280|false|false|false|||medicines
Event|Activity|Medications|10304,10313|false|false|false|C3241922|Operation Activity|operation
Event|Event|Medications|10304,10313|false|false|false|||operation
Procedure|Machine Activity|Medications|10304,10313|false|false|false|C0543467;C1880161|Computer Operation;Operative Surgical Procedures|operation
Procedure|Therapeutic or Preventive Procedure|Medications|10304,10313|false|false|false|C0543467;C1880161|Computer Operation;Operative Surgical Procedures|operation
Event|Event|Medications|10360,10364|false|false|false|||told
Event|Event|Medications|10396,10405|false|false|false|||questions
Drug|Pharmacologic Substance|Medications|10417,10425|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Event|Event|Medications|10417,10425|false|false|false|||medicine
Event|Event|Medications|10429,10433|false|false|false|||take
Procedure|Health Care Activity|Medications|10445,10449|false|false|false|C1515187|Take|take
Event|Event|Medications|10458,10462|false|false|false|||call
Attribute|Clinical Attribute|Medications|10468,10475|false|false|false|C5444295||surgeon
Disorder|Injury or Poisoning|Medications|10479,10484|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|WOUND
Event|Event|Medications|10479,10484|false|false|false|||WOUND
Finding|Body Substance|Medications|10479,10484|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|WOUND
Finding|Functional Concept|Medications|10479,10484|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|WOUND
Finding|Intellectual Product|Medications|10479,10484|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|WOUND
Procedure|Therapeutic or Preventive Procedure|Medications|10479,10489|false|false|false|C0886052;C1272654|Wound care management;wound care|WOUND CARE
Event|Activity|Medications|10485,10489|false|false|false|C1947933|care activity|CARE
Event|Event|Medications|10485,10489|false|false|false|||CARE
Finding|Finding|Medications|10485,10489|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|CARE
Finding|Intellectual Product|Medications|10485,10489|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|CARE
Drug|Biomedical or Dental Material|Medications|10494,10502|false|false|false|C1705365|Dressing Dosage Form|dressing
Event|Event|Medications|10494,10502|false|false|false|||dressing
Finding|Daily or Recreational Activity|Medications|10494,10502|false|false|false|C0518459;C1305428|Ability to dress|dressing
Finding|Finding|Medications|10494,10502|false|false|false|C0518459;C1305428|Ability to dress|dressing
Procedure|Health Care Activity|Medications|10494,10502|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Procedure|Therapeutic or Preventive Procedure|Medications|10494,10502|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Event|Activity|Medications|10503,10510|false|false|false|C1883720|Removing (action)|removal
Event|Event|Medications|10503,10510|false|false|false|||removal
Procedure|Therapeutic or Preventive Procedure|Medications|10503,10510|false|false|false|C0015252;C0185115;C0728940|Excision;Extraction;removal technique|removal
Event|Event|Medications|10522,10528|false|false|false|||remove
Event|Event|Medications|10534,10543|false|false|false|||dressings
Event|Event|Medications|10561,10567|false|false|false|||shower
Finding|Idea or Concept|Medications|10579,10582|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Medications|10579,10582|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biomedical or Dental Material|Medications|10592,10599|false|false|false|C2346961|Bandage Dosage Form|bandage
Event|Event|Medications|10600,10606|false|false|false|||strips
Event|Event|Medications|10619,10627|false|false|false|||covering
Event|Event|Medications|10648,10653|false|false|false|||scrub
Event|Event|Medications|10665,10669|false|false|false|||soak
Event|Event|Medications|10673,10677|false|false|false|||swim
Finding|Daily or Recreational Activity|Medications|10673,10677|false|false|false|C0039003|Swimming|swim
Disorder|Disease or Syndrome|Medications|10683,10686|false|false|false|C0030587|Paroxysmal atrial tachycardia|pat
Drug|Organic Chemical|Medications|10683,10686|false|false|false|C2825250|Fenamole|pat
Drug|Pharmacologic Substance|Medications|10683,10686|false|false|false|C2825250|Fenamole|pat
Event|Event|Medications|10683,10686|false|false|false|||pat
Finding|Molecular Function|Medications|10683,10686|false|false|false|C2247344;C2247346;C2248827|aspartate-prephenate aminotransferase activity;glutamate-prephenate aminotransferase activity;protein acetyltransferase activity|pat
Procedure|Diagnostic Procedure|Medications|10683,10686|false|false|false|C3897364|Thermoacoustic Computed Tomography|pat
Anatomy|Body Location or Region|Medications|10692,10700|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Medications|10692,10700|false|false|false|C0332803|Surgical wound|incision
Event|Event|Medications|10692,10700|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|Medications|10692,10700|false|false|false|C0184898|Surgical incisions|incision
Event|Event|Medications|10742,10746|false|false|false|||fall
Disorder|Disease or Syndrome|Medications|10791,10796|false|false|false|C1410088|Still|still
Event|Event|Medications|10791,10796|false|false|false|||still
Event|Event|Medications|10832,10839|false|false|false|||curling
Event|Event|Medications|10862,10866|false|false|false|||peel
Event|Event|Medications|10890,10895|false|false|false|||baths
Procedure|Health Care Activity|Medications|10890,10895|false|false|false|C0150141|Bathing|baths
Event|Event|Medications|10897,10901|false|false|false|||soak
Finding|Functional Concept|Medications|10897,10901|false|false|false|C1549544|Soak Administration|soak
Procedure|Therapeutic or Preventive Procedure|Medications|10897,10901|false|false|false|C0204774|Soak (procedure)|soak
Event|Event|Medications|10906,10910|false|false|false|||swim
Finding|Daily or Recreational Activity|Medications|10906,10910|false|false|false|C0039003|Swimming|swim
Finding|Finding|Medications|10923,10936|false|false|false|C0241311|post operative (finding)|after surgery
Event|Event|Medications|10929,10936|false|false|false|||surgery
Finding|Finding|Medications|10929,10936|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Medications|10929,10936|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Medications|10929,10936|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Medications|10929,10936|false|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Event|Medications|10945,10949|false|false|false|||told
Procedure|Health Care Activity|Medications|10968,10976|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|Medications|10968,10976|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Attribute|Clinical Attribute|Medications|10997,11004|false|false|false|C5444295||surgeon
Event|Event|Medications|11012,11018|false|false|false|||notice
Finding|Finding|Medications|11019,11027|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Finding|Idea or Concept|Medications|11019,11027|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Event|Event|Medications|11034,11042|false|false|false|||smelling
Finding|Organism Function|Medications|11034,11042|false|false|false|C0037361|Smell Perception|smelling
Event|Event|Medications|11045,11051|false|false|false|||bloody
Finding|Finding|Medications|11045,11051|false|false|false|C4554530|Bloody|bloody
Drug|Substance|Medications|11053,11056|false|false|false|C0444185|Pus specimen|pus
Event|Event|Medications|11053,11056|false|false|false|||pus
Finding|Body Substance|Medications|11053,11056|false|false|false|C0034161;C1546758|Pus;Pus Specimen Code|pus
Finding|Intellectual Product|Medications|11053,11056|false|false|false|C0034161;C1546758|Pus;Pus Specimen Code|pus
Finding|Idea or Concept|Medications|11058,11061|false|false|false|C1548556|Etc.|etc
Event|Event|Medications|11066,11075|false|false|false|||increased
Event|Event|Medications|11076,11084|false|false|false|||drainage
Finding|Body Substance|Medications|11076,11084|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|Medications|11076,11084|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|Medications|11076,11084|false|false|false|C0013103|Drainage procedure|drainage
Anatomy|Body Location or Region|Medications|11095,11103|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Medications|11095,11103|false|false|false|C0332803|Surgical wound|incision
Procedure|Therapeutic or Preventive Procedure|Medications|11095,11103|false|false|false|C0184898|Surgical incisions|incision
Anatomy|Body Location or Region|Medications|11104,11108|false|false|false|C1515974|Anatomic Site|site
Finding|Intellectual Product|Medications|11104,11108|false|false|false|C1546778||site
Event|Event|Medications|11111,11118|false|false|false|||opening
Anatomy|Body Location or Region|Medications|11127,11135|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Medications|11127,11135|false|false|false|C0332803|Surgical wound|incision
Event|Event|Medications|11127,11135|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|Medications|11127,11135|false|false|false|C0184898|Surgical incisions|incision
Finding|Finding|Medications|11140,11149|false|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Functional Concept|Medications|11140,11149|false|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Sign or Symptom|Medications|11140,11154|false|false|false|C5141269|Increased pain|increased pain
Attribute|Clinical Attribute|Medications|11150,11154|false|false|false|C2598155||pain
Event|Event|Medications|11150,11154|false|false|false|||pain
Finding|Functional Concept|Medications|11150,11154|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Medications|11150,11154|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Disorder|Injury or Poisoning|Medications|11158,11166|false|false|false|C0009938|Contusions|bruising
Event|Event|Medications|11158,11166|false|false|false|||bruising
Finding|Finding|Medications|11158,11166|false|false|false|C2136686|reported bruising (history)|bruising
Event|Event|Medications|11179,11184|false|false|false|||signs
Finding|Finding|Medications|11179,11184|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Medications|11179,11184|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Disorder|Disease or Syndrome|Medications|11188,11197|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|Medications|11188,11197|false|false|false|||infection
Finding|Pathologic Function|Medications|11188,11197|false|false|false|C3714514|Infection|infection
Disorder|Disease or Syndrome|Medications|11206,11213|false|false|false|C0041834|Erythema|redness
Event|Event|Medications|11206,11213|false|false|false|||redness
Finding|Finding|Medications|11206,11213|false|false|false|C0332575|Redness|redness
Event|Event|Medications|11215,11224|false|false|false|||streaking
Anatomy|Body System|Medications|11233,11237|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|Medications|11233,11237|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|Medications|11233,11237|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Finding|Body Substance|Medications|11233,11237|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|Medications|11233,11237|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Event|Event|Medications|11240,11248|false|false|false|||swelling
Finding|Finding|Medications|11240,11248|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|Medications|11240,11248|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Finding|Medications|11250,11259|false|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Functional Concept|Medications|11250,11259|false|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Sign or Symptom|Medications|11250,11264|false|false|false|C5141269|Increased pain|increased pain
Attribute|Clinical Attribute|Medications|11260,11264|false|false|false|C2598155||pain
Event|Event|Medications|11260,11264|false|false|false|||pain
Finding|Functional Concept|Medications|11260,11264|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Medications|11260,11264|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Medications|11279,11287|false|false|false|||drainage
Finding|Body Substance|Medications|11279,11287|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|Medications|11279,11287|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|Medications|11279,11287|false|false|false|C0013103|Drainage procedure|drainage
Event|Event|Medications|11298,11302|false|false|false|||call
Event|Event|Medications|11312,11321|false|false|false|||questions
Event|Event|Medications|11325,11333|false|false|false|||concerns
Event|Event|Medications|11350,11358|false|false|false|||allowing
Event|Event|Medications|11365,11376|false|false|false|||participate
Event|Activity|Medications|11385,11389|false|false|false|C1947933|care activity|care
Event|Event|Medications|11385,11389|false|false|false|||care
Finding|Finding|Medications|11385,11389|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Medications|11385,11389|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Event|Event|Medications|11417,11423|false|false|false|||return
Event|Event|Medications|11438,11442|false|false|false|||life
Finding|Idea or Concept|Medications|11438,11442|false|false|false|C0376558|Life|life
Procedure|Diagnostic Procedure|Medications|11438,11442|false|false|false|C1522684|Laser-Induced Fluorescence Endoscopy|life
Event|Activity|Medications|11447,11457|false|false|false|C0441655|Activities|activities
Event|Event|Medications|11447,11457|false|false|false|||activities
Finding|Finding|Medications|11447,11457|false|false|false|C2239122|activities (history)|activities
Event|Event|Medications|11460,11464|false|false|false|||Home
Finding|Idea or Concept|Medications|11460,11464|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Medications|11460,11464|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Medications|11460,11464|false|false|false|C1553498|home health encounter|Home
Event|Event|Medications|11491,11499|false|false|false|||catheter
Finding|Intellectual Product|Medications|11491,11499|false|false|false|C1546572||catheter
Anatomy|Body Part, Organ, or Organ Component|Medications|11508,11515|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|Medications|11508,11515|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Event|Event|Medications|11508,11515|false|false|false|||bladder
Procedure|Therapeutic or Preventive Procedure|Medications|11508,11515|false|false|false|C0872388|Procedures on bladder|bladder
Event|Event|Medications|11516,11522|false|false|false|||placed
Finding|Idea or Concept|Medications|11542,11545|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Medications|11542,11545|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Medications|11554,11561|false|false|false|||surgery
Finding|Finding|Medications|11554,11561|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Medications|11554,11561|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Medications|11554,11561|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Medications|11554,11561|false|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Event|Medications|11568,11578|false|false|false|||difficulty
Finding|Finding|Medications|11568,11578|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Event|Event|Medications|11579,11585|false|false|false|||trying
Event|Event|Medications|11589,11594|false|false|false|||place
Event|Event|Medications|11608,11612|false|false|false|||keep
Event|Event|Medications|11617,11625|false|false|false|||catheter
Finding|Intellectual Product|Medications|11617,11625|false|false|false|C1546572||catheter
Event|Activity|Medications|11637,11648|false|false|false|C0003629|Appointments|appointment
Event|Event|Medications|11637,11648|false|false|false|||appointment
Event|Event|Medications|11681,11685|false|false|false|||call
Event|Event|Medications|11690,11696|false|false|false|||number
Finding|Idea or Concept|Medications|11690,11696|false|false|false|C1554106|MDF AttributeType - Number|number
Event|Event|Medications|11706,11714|false|false|false|||schedule
Event|Activity|Medications|11721,11732|false|false|false|C0003629|Appointments|appointment
Event|Event|Medications|11721,11732|false|false|false|||appointment
Event|Event|Medications|11744,11750|false|false|false|||decide
Event|Event|Medications|11758,11762|false|false|false|||need
Event|Event|Medications|11776,11783|false|false|false|||attempt
Event|Event|Medications|11776,11783|false|false|false|C1516084|Attempt|attempt
Event|Event|Medications|11788,11794|false|false|false|||remove
Event|Event|Medications|11802,11805|false|false|false|||see
Event|Event|Medications|11817,11821|false|false|false|||able
Finding|Finding|Medications|11817,11821|false|false|false|C1299581|Able (qualifier value)|able
Event|Event|Medications|11825,11829|false|false|false|||void
Finding|Functional Concept|Medications|11832,11837|false|false|false|C5848602|Exhausted|Empty
Finding|Intellectual Product|Medications|11842,11845|false|false|false|C1552710|Bag Data Type|bag
Event|Event|Medications|11849,11855|false|false|false|||needed
Event|Event|Medications|11863,11868|false|false|false|||shown
Finding|Organism Function|Medications|11879,11886|false|false|false|C0006147|Breast Feeding|nursing
Procedure|Therapeutic or Preventive Procedure|Medications|11879,11886|false|false|false|C0028678|RNAx nursing therapy actions|nursing
Event|Event|Medications|11887,11892|false|false|false|||staff
Finding|Finding|Medications|11887,11892|false|false|false|C1551040|Encounter Special Courtesy - staff|staff
Anatomy|Body Part, Organ, or Organ Component|Medications|11915,11918|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Event|Event|Medications|11919,11922|false|false|false|||bag
Finding|Intellectual Product|Medications|11919,11922|false|false|false|C1552710|Bag Data Type|bag
Event|Event|Medications|11935,11944|false|false|false|||discharge
Finding|Body Substance|Medications|11935,11944|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Medications|11935,11944|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Medications|11935,11944|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Medications|11935,11944|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|Medications|11960,11963|false|false|false|||use
Finding|Functional Concept|Medications|11960,11963|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|Medications|11960,11963|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Phenomenon|Phenomenon or Process|Medications|11974,11979|false|false|false|C0221188|Tripping|trips
Event|Event|Medications|11999,12002|false|false|false|||bag
Finding|Intellectual Product|Medications|11999,12002|false|false|false|C1552710|Bag Data Type|bag
Anatomy|Body Part, Organ, or Organ Component|Medications|12024,12027|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Event|Event|Medications|12037,12041|false|false|false|||home
Finding|Idea or Concept|Medications|12037,12041|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Medications|12037,12041|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Medications|12037,12041|false|false|false|C1553498|home health encounter|home
Event|Event|Medications|12046,12050|false|false|false|||wear
Event|Event|Medications|12062,12071|false|false|false|||traveling
Event|Event|Medications|12086,12090|false|false|false|||home
Finding|Idea or Concept|Medications|12086,12090|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Medications|12086,12090|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Medications|12086,12090|false|false|false|C1553498|home health encounter|home
Event|Event|Medications|12097,12102|false|false|false|||holds
Finding|Intellectual Product|Medications|12113,12119|false|false|false|C1561574|Amount class - Amount|amount
Finding|Intellectual Product|Medications|12129,12132|false|false|false|C1552710|Bag Data Type|bag
Event|Event|Medications|12154,12159|false|false|false|||needs
Event|Event|Medications|12166,12173|false|false|false|||emptied
Finding|Intellectual Product|Medications|12179,12184|false|false|false|C4050225|Often - answer to question|often
Event|Event|Medications|12198,12202|false|false|false|||find
Event|Event|Medications|12217,12220|false|false|false|||use
Disorder|Disease or Syndrome|Medications|12232,12235|false|false|false|C4522181|Brachial Amyotrophic Diplegia|bad
Drug|Amino Acid, Peptide, or Protein|Medications|12232,12235|false|false|false|C1530798|BAD protein, human|bad
Drug|Biologically Active Substance|Medications|12232,12235|false|false|false|C1530798|BAD protein, human|bad
Event|Event|Medications|12232,12235|false|false|false|||bad
Finding|Gene or Genome|Medications|12232,12235|false|false|false|C1366450|BAD gene|bad
Finding|Finding|Medications|12250,12257|false|false|false|C4534363|At home|at home
Event|Event|Medications|12253,12257|false|false|false|||home
Finding|Idea or Concept|Medications|12253,12257|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Medications|12253,12257|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Medications|12253,12257|false|false|false|C1553498|home health encounter|home
Event|Event|Medications|12261,12266|false|false|false|||carry
Event|Activity|Medications|12295,12299|false|false|false|C1947933|care activity|Care
Finding|Finding|Medications|12295,12299|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Medications|12295,12299|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Attribute|Clinical Attribute|Medications|12295,12304|false|false|false|C4321316||Care Team
Finding|Finding|Medications|12295,12304|false|false|false|C4321315|Care team|Care Team
Procedure|Health Care Activity|Medications|12307,12315|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Medications|12316,12328|false|false|false|C3263700||Instructions
Event|Event|Medications|12316,12328|false|false|false|||Instructions
Finding|Intellectual Product|Medications|12316,12328|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

