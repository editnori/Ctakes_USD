 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|28,32
No|33,35
:|35,36
_|39,40
_|40,41
_|41,42
<EOL>|42,43
<EOL>|44,45
Admission|45,54
Date|55,59
:|59,60
_|62,63
_|63,64
_|64,65
Discharge|79,88
Date|89,93
:|93,94
_|97,98
_|98,99
_|99,100
<EOL>|100,101
<EOL>|102,103
Date|103,107
of|108,110
Birth|111,116
:|116,117
_|119,120
_|120,121
_|121,122
Sex|135,138
:|138,139
M|142,143
<EOL>|143,144
<EOL>|145,146
Service|146,153
:|153,154
PSYCHIATRY|155,165
<EOL>|165,166
<EOL>|167,168
Allergies|168,177
:|177,178
<EOL>|179,180
Patient|180,187
recorded|188,196
as|197,199
having|200,206
No|207,209
Known|210,215
Allergies|216,225
to|226,228
Drugs|229,234
<EOL>|234,235
<EOL>|236,237
Attending|237,246
:|246,247
_|248,249
_|249,250
_|250,251
<EOL>|251,252
<EOL>|253,254
Chief|254,259
Complaint|260,269
:|269,270
<EOL>|270,271
I|271,272
have|273,277
been|278,282
overwhelmed|283,294
and|295,298
I|299,300
felt|301,305
suicidal|306,314
.|314,315
"|315,316
<EOL>|316,317
<EOL>|317,318
<EOL>|319,320
Major|320,325
Surgical|326,334
or|335,337
Invasive|338,346
Procedure|347,356
:|356,357
<EOL>|357,358
none|358,362
<EOL>|362,363
<EOL>|363,364
<EOL>|365,366
History|366,373
of|374,376
Present|377,384
Illness|385,392
:|392,393
<EOL>|393,394
HPI|394,397
:|397,398
Mr.|400,403
_|404,405
_|405,406
_|406,407
is|408,410
a|411,412
_|413,414
_|414,415
_|415,416
yo|417,419
_|420,421
_|421,422
_|422,423
freshman|424,432
at|433,435
_|436,437
_|437,438
_|438,439
(|440,441
_|441,442
_|442,443
_|443,444
)|444,445
c|446,447
h|448,449
/|449,450
o|450,451
depressed|452,461
mood|462,466
and|467,470
anxiety|471,478
symptoms|479,487
<EOL>|487,488
(|488,489
panic|489,494
)|494,495
who|496,499
was|500,503
sent|504,508
to|509,511
_|512,513
_|513,514
_|514,515
at|516,518
recommendation|519,533
of|534,536
_|537,538
_|538,539
_|539,540
,|540,541
his|542,545
<EOL>|545,546
therapist|546,555
of|556,558
4|559,560
months|561,567
at|568,570
_|571,572
_|572,573
_|573,574
for|575,578
evaluation|579,589
of|590,592
3|593,594
weeks|595,600
of|601,603
<EOL>|603,604
worsening|604,613
depression|614,624
with|625,629
anhedonia|630,639
,|639,640
social|641,647
isolation|648,657
&|658,659
<EOL>|659,660
withdrawal|660,670
,|670,671
escalating|672,682
feelings|683,691
of|692,694
guilt|695,700
,|700,701
poor|702,706
sleep|707,712
secondary|713,722
<EOL>|723,724
to|724,726
<EOL>|726,727
ruminations|727,738
of|739,741
guilt|742,747
.|747,748
Patient|750,757
is|758,760
also|761,765
having|766,772
trouble|773,780
<EOL>|780,781
concentrating|781,794
and|795,798
going|799,804
to|805,807
his|808,811
other|812,817
classes|818,825
because|826,833
of|834,836
his|837,840
<EOL>|840,841
depression|841,851
and|852,855
anxiety|856,863
.|863,864
He|866,868
has|869,872
been|873,877
eating|878,884
fine|885,889
and|890,893
taking|894,900
care|901,905
<EOL>|905,906
of|906,908
himself|909,916
w|917,918
/|918,919
r|919,920
/|920,921
t|921,922
hygiene|923,930
.|930,931
Mr.|933,936
_|937,938
_|938,939
_|939,940
reported|941,949
that|950,954
what|955,959
seems|960,965
<EOL>|965,966
have|966,970
caused|971,977
his|978,981
recent|982,988
bout|989,993
of|994,996
anxiety|997,1004
is|1005,1007
the|1008,1011
culmination|1012,1023
of|1024,1026
<EOL>|1026,1027
stress|1027,1033
in|1034,1036
a|1037,1038
professional|1039,1051
relationship|1052,1064
with|1065,1069
one|1070,1073
of|1074,1076
his|1077,1080
teachers|1081,1089
<EOL>|1090,1091
at|1091,1093
<EOL>|1093,1094
his|1094,1097
program|1098,1105
.|1105,1106
For|1108,1111
reasons|1112,1119
that|1120,1124
are|1125,1128
not|1129,1132
completely|1133,1143
clear|1144,1149
,|1149,1150
patient|1151,1158
<EOL>|1158,1159
was|1159,1162
removed|1163,1170
from|1171,1175
a|1176,1177
studio|1178,1184
class|1185,1190
with|1191,1195
a|1196,1197
particular|1198,1208
instructor|1209,1219
.|1219,1220
<EOL>|1221,1222
Patient|1222,1229
referred|1230,1238
me|1239,1241
to|1242,1244
speak|1245,1250
with|1251,1255
_|1256,1257
_|1257,1258
_|1258,1259
to|1260,1262
explain|1263,1270
the|1271,1274
<EOL>|1275,1276
specifics|1276,1285
,|1285,1286
<EOL>|1286,1287
but|1287,1290
_|1291,1292
_|1292,1293
_|1293,1294
was|1295,1298
not|1299,1302
available|1303,1312
and|1313,1316
patient|1317,1324
felt|1325,1329
too|1330,1333
<EOL>|1333,1334
overwhelmed|1334,1345
to|1346,1348
give|1349,1353
me|1354,1356
the|1357,1360
story|1361,1366
in|1367,1369
detail|1370,1376
-|1376,1377
-|1377,1378
in|1378,1380
fact|1381,1385
had|1386,1389
a|1390,1391
panic|1392,1397
<EOL>|1397,1398
attack|1398,1404
during|1405,1411
our|1412,1415
talk|1416,1420
.|1420,1421
For|1423,1426
the|1427,1430
past|1431,1435
weeks|1436,1441
,|1441,1442
since|1443,1448
being|1449,1454
removed|1455,1462
<EOL>|1462,1463
from|1463,1467
the|1468,1471
class|1472,1477
,|1477,1478
Mr.|1479,1482
_|1483,1484
_|1484,1485
_|1485,1486
has|1487,1490
written|1491,1498
letters|1499,1506
,|1506,1507
called|1508,1514
(|1515,1516
did|1516,1519
<EOL>|1520,1521
not|1521,1524
<EOL>|1524,1525
leave|1525,1530
messages|1531,1539
)|1539,1540
and|1541,1544
emailed|1545,1552
this|1553,1557
instructor|1558,1568
w|1569,1570
/|1570,1571
o|1571,1572
getting|1573,1580
any|1581,1584
<EOL>|1584,1585
response|1585,1593
.|1593,1594
The|1596,1599
lack|1600,1604
of|1605,1607
response|1608,1616
has|1617,1620
caused|1621,1627
an|1628,1630
escalating|1631,1641
pattern|1642,1649
<EOL>|1649,1650
of|1650,1652
guilt|1653,1658
that|1659,1663
Mr.|1664,1667
_|1668,1669
_|1669,1670
_|1670,1671
has|1672,1675
been|1676,1680
dealing|1681,1688
with|1689,1693
by|1694,1696
cutting|1697,1704
<EOL>|1704,1705
himself|1705,1712
with|1713,1717
a|1718,1719
knife|1720,1725
(|1726,1727
cut|1727,1730
left|1731,1735
wrist|1736,1741
,|1741,1742
no|1743,1745
stitches|1746,1754
)|1754,1755
.|1755,1756
Last|1758,1762
night|1763,1768
,|1768,1769
<EOL>|1769,1770
in|1770,1772
the|1773,1776
context|1777,1784
of|1785,1787
this|1788,1792
guilt|1793,1798
,|1798,1799
not|1800,1803
sleeping|1804,1812
and|1813,1816
having|1817,1823
more|1824,1828
<EOL>|1828,1829
anxiety|1829,1836
,|1836,1837
Mr.|1838,1841
_|1842,1843
_|1843,1844
_|1844,1845
began|1846,1851
feeling|1852,1859
suicidal|1860,1868
and|1869,1872
developed|1873,1882
a|1883,1884
<EOL>|1885,1886
plan|1886,1890
<EOL>|1890,1891
to|1891,1893
kill|1894,1898
himself|1899,1906
by|1907,1909
cutting|1910,1917
himself|1918,1925
with|1926,1930
a|1931,1932
knife|1933,1938
.|1938,1939
He|1941,1943
decided|1944,1951
<EOL>|1952,1953
that|1953,1957
<EOL>|1957,1958
the|1958,1961
only|1962,1966
way|1967,1970
he|1971,1973
could|1974,1979
deal|1980,1984
with|1985,1989
his|1990,1993
overwhelming|1994,2006
feelings|2007,2015
would|2016,2021
<EOL>|2021,2022
be|2022,2024
suicide|2025,2032
.|2032,2033
Mr.|2035,2038
_|2039,2040
_|2040,2041
_|2041,2042
told|2043,2047
his|2048,2051
counselor|2052,2061
about|2062,2067
these|2068,2073
<EOL>|2074,2075
thoughts|2075,2083
<EOL>|2083,2084
and|2084,2087
his|2088,2091
counselor|2092,2101
recommended|2102,2113
that|2114,2118
he|2119,2121
come|2122,2126
to|2127,2129
the|2130,2133
ED|2134,2136
.|2136,2137
<EOL>|2139,2140
<EOL>|2140,2141
Mr.|2141,2144
_|2145,2146
_|2146,2147
_|2147,2148
reported|2149,2157
that|2158,2162
he|2163,2165
has|2166,2169
felt|2170,2174
"|2175,2176
highs|2176,2181
,|2181,2182
"|2182,2183
but|2184,2187
never|2188,2193
for|2194,2197
<EOL>|2197,2198
more|2198,2202
than|2203,2207
a|2208,2209
day|2210,2213
and|2214,2217
never|2218,2223
impacting|2224,2233
sleep|2234,2239
or|2240,2242
resulting|2243,2252
in|2253,2255
<EOL>|2255,2256
dramatically|2256,2268
impaired|2269,2277
decision|2278,2286
-|2286,2287
making|2287,2293
(|2294,2295
e.g|2295,2298
.|2298,2299
,|2299,2300
spending|2301,2309
too|2310,2313
much|2314,2318
,|2318,2319
<EOL>|2319,2320
indiscriminate|2320,2334
sexual|2335,2341
relationships|2342,2355
,|2355,2356
etc|2357,2360
)|2360,2361
.|2361,2362
Mr.|2364,2367
_|2368,2369
_|2369,2370
_|2370,2371
has|2372,2375
no|2376,2378
<EOL>|2378,2379
h|2379,2380
/|2380,2381
o|2381,2382
_|2383,2384
_|2384,2385
_|2385,2386
psychotic|2387,2396
symptoms|2397,2405
,|2405,2406
although|2407,2415
his|2416,2419
level|2420,2425
of|2426,2428
guilt|2429,2434
has|2435,2438
<EOL>|2438,2439
reached|2439,2446
a|2447,2448
near|2449,2453
psychotic|2454,2463
proportion|2464,2474
.|2474,2475
Mr.|2477,2480
_|2481,2482
_|2482,2483
_|2483,2484
denied|2485,2491
ever|2492,2496
<EOL>|2496,2497
being|2497,2502
asked|2503,2508
by|2509,2511
the|2512,2515
instructor|2516,2526
never|2527,2532
to|2533,2535
contact|2536,2543
him|2544,2547
,|2547,2548
but|2549,2552
he|2553,2555
feels|2556,2561
<EOL>|2561,2562
the|2562,2565
instructor|2566,2576
not|2577,2580
answering|2581,2590
his|2591,2594
calls|2595,2600
or|2601,2603
responding|2604,2614
to|2615,2617
emails|2618,2624
<EOL>|2624,2625
means|2625,2630
that|2631,2635
the|2636,2639
instructor|2640,2650
does|2651,2655
not|2656,2659
like|2660,2664
him|2665,2668
.|2668,2669
He|2671,2673
denied|2674,2680
any|2681,2684
<EOL>|2684,2685
thoughts|2685,2693
of|2694,2696
trying|2697,2703
to|2704,2706
harm|2707,2711
the|2712,2715
instructor|2716,2726
.|2726,2727
<EOL>|2729,2730
<EOL>|2730,2731
Mr.|2731,2734
_|2735,2736
_|2736,2737
_|2737,2738
reported|2739,2747
feeling|2748,2755
anxious|2756,2763
a|2764,2765
great|2766,2771
deal|2772,2776
,|2776,2777
having|2778,2784
a|2785,2786
<EOL>|2787,2788
rare|2788,2792
<EOL>|2792,2793
panic|2793,2798
attack|2799,2805
.|2805,2806
<EOL>|2807,2808
<EOL>|2808,2809
<EOL>|2810,2811
Past|2811,2815
Medical|2816,2823
History|2824,2831
:|2831,2832
<EOL>|2832,2833
PAST|2833,2837
PSYCH|2838,2843
HX|2844,2846
:|2846,2847
No|2849,2851
previous|2852,2860
medication|2861,2871
trials|2872,2878
or|2879,2881
psychiatric|2882,2893
<EOL>|2893,2894
hospitalizations|2894,2910
.|2910,2911
One|2913,2916
previous|2917,2925
episode|2926,2933
of|2934,2936
being|2937,2942
kept|2943,2947
in|2948,2950
a|2951,2952
<EOL>|2952,2953
psychiatric|2953,2964
ED|2965,2967
in|2968,2970
_|2971,2972
_|2972,2973
_|2973,2974
in|2975,2977
the|2978,2981
context|2982,2989
of|2990,2992
having|2993,2999
chest|3000,3005
<EOL>|3005,3006
pain|3006,3010
which|3011,3016
turned|3017,3023
out|3024,3027
to|3028,3030
be|3031,3033
a|3034,3035
panic|3036,3041
attack|3042,3048
.|3048,3049
Gets|3051,3055
occasional|3056,3066
<EOL>|3066,3067
panic|3067,3072
attacks|3073,3080
(|3081,3082
although|3082,3090
not|3091,3094
frequently|3095,3105
enough|3106,3112
to|3113,3115
make|3116,3120
a|3121,3122
<EOL>|3123,3124
diagnosis|3124,3133
<EOL>|3133,3134
of|3134,3136
panic|3137,3142
d|3143,3144
/|3144,3145
o|3145,3146
)|3146,3147
.|3147,3148
Has|3150,3153
been|3154,3158
seeing|3159,3165
a|3166,3167
counselor|3168,3177
_|3178,3179
_|3179,3180
_|3180,3181
at|3182,3184
_|3185,3186
_|3186,3187
_|3187,3188
x|3189,3190
4|3191,3192
<EOL>|3192,3193
months|3193,3199
.|3199,3200
Prior|3202,3207
to|3208,3210
3|3211,3212
weeks|3213,3218
ago|3219,3222
,|3222,3223
no|3224,3226
h|3227,3228
/|3228,3229
o|3229,3230
self|3231,3235
-|3235,3236
injurious|3236,3245
behaviors|3246,3255
,|3255,3256
<EOL>|3256,3257
although|3257,3265
has|3266,3269
had|3270,3273
suicidal|3274,3282
ideation|3283,3291
in|3292,3294
the|3295,3298
past|3299,3303
(|3304,3305
once|3305,3309
or|3310,3312
twice|3313,3318
<EOL>|3318,3319
prior|3319,3324
to|3325,3327
last|3328,3332
night|3333,3338
,|3338,3339
but|3340,3343
never|3344,3349
with|3350,3354
intent|3355,3361
like|3362,3366
now|3367,3370
)|3370,3371
.|3371,3372
Saw|3374,3377
a|3378,3379
<EOL>|3379,3380
counselor|3380,3389
in|3390,3392
high|3393,3397
school|3398,3404
to|3405,3407
help|3408,3412
with|3413,3417
"|3418,3419
coping|3419,3425
"|3425,3426
with|3427,3431
feeling|3432,3439
<EOL>|3439,3440
different|3440,3449
in|3450,3452
school|3453,3459
.|3459,3460
<EOL>|3460,3461
<EOL>|3461,3462
Mr.|3462,3465
_|3466,3467
_|3467,3468
_|3468,3469
reported|3470,3478
that|3479,3483
he|3484,3486
had|3487,3490
thoughts|3491,3499
of|3500,3502
fighting|3503,3511
with|3512,3516
a|3517,3518
<EOL>|3518,3519
fellow|3519,3525
student|3526,3533
a|3534,3535
few|3536,3539
months|3540,3546
ago|3547,3550
,|3550,3551
which|3552,3557
is|3558,3560
why|3561,3564
he|3565,3567
started|3568,3575
in|3576,3578
<EOL>|3578,3579
counseling|3579,3589
(|3590,3591
he|3591,3593
said|3594,3598
he|3599,3601
did|3602,3605
not|3606,3609
want|3610,3614
to|3615,3617
get|3618,3621
into|3622,3626
details|3627,3634
re|3635,3637
.|3637,3638
that|3639,3643
<EOL>|3643,3644
situation|3644,3653
)|3653,3654
.|3654,3655
He|3656,3658
said|3659,3663
that|3664,3668
ultimately|3669,3679
he|3680,3682
was|3683,3686
able|3687,3691
to|3692,3694
come|3695,3699
to|3700,3702
terms|3703,3708
<EOL>|3708,3709
with|3709,3713
this|3714,3718
person|3719,3725
w|3726,3727
/|3727,3728
o|3728,3729
fighting|3730,3738
.|3738,3739
He|3741,3743
denied|3744,3750
any|3751,3754
h|3755,3756
/|3756,3757
o|3757,3758
violent|3759,3766
<EOL>|3766,3767
behavior|3767,3775
.|3775,3776
<EOL>|3776,3777
<EOL>|3777,3778
PMH|3778,3781
:|3781,3782
Essentially|3784,3795
healthy|3796,3803
young|3804,3809
man|3810,3813
.|3813,3814
Had|3816,3819
repair|3820,3826
of|3827,3829
meniscus|3830,3838
of|3839,3841
<EOL>|3841,3842
left|3842,3846
knee|3847,3851
several|3852,3859
months|3860,3866
ago|3867,3870
secondary|3871,3880
to|3881,3883
injury|3884,3890
while|3891,3896
running|3897,3904
.|3904,3905
<EOL>|3906,3907
No|3907,3909
other|3910,3915
surgeries|3916,3925
.|3925,3926
<EOL>|3926,3927
<EOL>|3927,3928
<EOL>|3929,3930
Social|3930,3936
History|3937,3944
:|3944,3945
<EOL>|3945,3946
_|3946,3947
_|3947,3948
_|3948,3949
<EOL>|3949,3950
SOCIAL|3950,3956
/|3956,3957
FAMILY|3957,3963
HX|3964,3966
:|3966,3967
Only|3969,3973
child|3974,3979
born|3980,3984
to|3985,3987
now|3988,3991
divorced|3992,4000
parents|4001,4008
.|4008,4009
<EOL>|4010,4011
Parents|4011,4018
separated|4019,4028
when|4029,4033
patient|4034,4041
was|4042,4045
_|4046,4047
_|4047,4048
_|4048,4049
.|4049,4050
Raised|4052,4058
by|4059,4061
mother|4062,4068
in|4069,4071
<EOL>|4071,4072
_|4072,4073
_|4073,4074
_|4074,4075
,|4075,4076
but|4077,4080
also|4081,4085
has|4086,4089
a|4090,4091
relationship|4092,4104
with|4105,4109
father|4110,4116
.|4116,4117
Father|4119,4125
<EOL>|4125,4126
struggled|4126,4135
with|4136,4140
active|4141,4147
alcohol|4148,4155
dependence|4156,4166
for|4167,4170
many|4171,4175
years|4176,4181
,|4181,4182
but|4183,4186
is|4187,4189
<EOL>|4189,4190
now|4190,4193
sober|4194,4199
.|4199,4200
Patient|4202,4209
denied|4210,4216
any|4217,4220
h|4221,4222
/|4222,4223
o|4223,4224
physical|4225,4233
or|4234,4236
sexual|4237,4243
abuse|4244,4249
<EOL>|4250,4251
while|4251,4256
<EOL>|4256,4257
growing|4257,4264
up|4265,4267
.|4267,4268
Described|4270,4279
feeling|4280,4287
"|4288,4289
different|4289,4298
"|4298,4299
and|4300,4303
having|4304,4310
trouble|4311,4318
<EOL>|4318,4319
fitting|4319,4326
in|4327,4329
,|4329,4330
but|4331,4334
could|4335,4340
not|4341,4344
give|4345,4349
more|4350,4354
details|4355,4362
.|4362,4363
Had|4365,4368
some|4369,4373
<EOL>|4374,4375
behavioral|4375,4385
<EOL>|4385,4386
troubles|4386,4394
in|4395,4397
school|4398,4404
as|4405,4407
a|4408,4409
child|4410,4415
,|4415,4416
was|4417,4420
suspended|4421,4430
at|4431,4433
least|4434,4439
3|4440,4441
times|4442,4447
in|4448,4450
<EOL>|4450,4451
high|4451,4455
school|4456,4462
,|4462,4463
struggled|4464,4473
academically|4474,4486
,|4486,4487
but|4488,4491
did|4492,4495
graduate|4496,4504
.|4504,4505
<EOL>|4507,4508
Currently|4508,4517
<EOL>|4517,4518
a|4518,4519
freshman|4520,4528
at|4529,4531
_|4532,4533
_|4533,4534
_|4534,4535
with|4536,4540
an|4541,4543
area|4544,4548
of|4549,4551
concentration|4552,4565
in|4566,4568
the|4569,4572
clarinet|4573,4581
,|4581,4582
<EOL>|4582,4583
but|4583,4586
having|4587,4593
a|4594,4595
difficult|4596,4605
time|4606,4610
as|4611,4613
above|4614,4619
.|4619,4620
Mr.|4622,4625
_|4626,4627
_|4627,4628
_|4628,4629
lives|4630,4635
alone|4636,4641
<EOL>|4641,4642
in|4642,4644
student|4645,4652
housing|4653,4660
.|4660,4661
No|4663,4665
current|4666,4673
romantic|4674,4682
relationships|4683,4696
,|4696,4697
has|4698,4701
<EOL>|4702,4703
dated|4703,4708
<EOL>|4708,4709
a|4709,4710
girl|4711,4715
in|4716,4718
the|4719,4722
past|4723,4727
,|4727,4728
but|4729,4732
the|4733,4736
relationship|4737,4749
ended|4750,4755
because|4756,4763
the|4764,4767
girl|4768,4772
<EOL>|4772,4773
did|4773,4776
not|4777,4780
feel|4781,4785
ready|4786,4791
to|4792,4794
continue|4795,4803
.|4803,4804
Mr.|4806,4809
_|4810,4811
_|4811,4812
_|4812,4813
denied|4814,4820
any|4821,4824
legal|4825,4830
<EOL>|4830,4831
problems|4831,4839
and|4840,4843
denied|4844,4850
having|4851,4857
access|4858,4864
to|4865,4867
any|4868,4871
guns|4872,4876
.|4876,4877
<EOL>|4879,4880
<EOL>|4880,4881
<EOL>|4882,4883
Family|4883,4889
History|4890,4897
:|4897,4898
<EOL>|4898,4899
Family|4899,4905
history|4906,4913
remarkable|4914,4924
for|4925,4928
father|4929,4935
with|4936,4940
alcohol|4941,4948
problems|4949,4957
(|4958,4959
in|4959,4961
<EOL>|4961,4962
remission|4962,4971
)|4971,4972
and|4973,4976
mother|4977,4983
with|4984,4988
h|4989,4990
/|4990,4991
o|4991,4992
hypothyroidism|4993,5007
.|5007,5008
No|5010,5012
other|5013,5018
family|5019,5025
<EOL>|5025,5026
medical|5026,5033
or|5034,5036
psychiatric|5037,5048
problems|5049,5057
known|5058,5063
by|5064,5066
patient|5067,5074
.|5074,5075
<EOL>|5075,5076
<EOL>|5076,5077
<EOL>|5078,5079
Physical|5079,5087
Exam|5088,5092
:|5092,5093
<EOL>|5093,5094
MSE|5094,5097
-|5097,5098
Mr.|5099,5102
_|5103,5104
_|5104,5105
_|5105,5106
is|5107,5109
a|5110,5111
<EOL>|5111,5112
_|5112,5113
_|5113,5114
_|5114,5115
white|5116,5121
male|5122,5126
,|5126,5127
dressed|5128,5135
in|5136,5138
hospital|5139,5147
_|5148,5149
_|5149,5150
_|5150,5151
.|5151,5152
Appears|5154,5161
<EOL>|5161,5162
anxious|5162,5169
,|5169,5170
had|5171,5174
a|5175,5176
panic|5177,5182
attack|5183,5189
during|5190,5196
the|5197,5200
interview|5201,5210
.|5210,5211
Speech|5213,5219
normal|5220,5226
<EOL>|5226,5227
rate|5227,5231
,|5231,5232
tone|5233,5237
&|5238,5239
volume|5240,5246
.|5246,5247
Normal|5249,5255
language|5256,5264
.|5264,5265
Mood|5267,5271
is|5272,5274
"|5275,5276
depressed|5276,5285
"|5285,5286
with|5287,5291
<EOL>|5291,5292
a|5292,5293
constricted|5294,5305
affective|5306,5315
range|5316,5321
in|5322,5324
anxious|5325,5332
realm|5333,5338
.|5338,5339
Thoughts|5341,5349
<EOL>|5349,5350
organized|5350,5359
,|5359,5360
but|5361,5364
themes|5365,5371
of|5372,5374
guilt|5375,5380
.|5380,5381
Endorsed|5383,5391
suicidal|5392,5400
ideation|5401,5409
with|5410,5414
<EOL>|5414,5415
plan|5415,5419
to|5420,5422
commit|5423,5429
suicide|5430,5437
using|5438,5443
a|5444,5445
knife|5446,5451
to|5452,5454
cut|5455,5458
himself|5459,5466
,|5466,5467
vacillating|5468,5479
<EOL>|5479,5480
intent|5480,5486
.|5486,5487
Denied|5489,5495
thoughts|5496,5504
of|5505,5507
harming|5508,5515
others|5516,5522
.|5522,5523
Insight|5525,5532
into|5533,5537
need|5538,5542
<EOL>|5542,5543
for|5543,5546
help|5547,5551
is|5552,5554
good|5555,5559
,|5559,5560
judgment|5561,5569
fair|5570,5574
.|5574,5575
<EOL>|5575,5576
<EOL>|5576,5577
<EOL>|5578,5579
Pertinent|5579,5588
Results|5589,5596
:|5596,5597
<EOL>|5597,5598
_|5598,5599
_|5599,5600
_|5600,5601
03|5602,5604
:|5604,5605
58PM|5605,5609
GLUCOSE|5612,5619
-|5619,5620
96|5620,5622
UREA|5623,5627
N|5628,5629
-|5629,5630
17|5630,5632
CREAT|5633,5638
-|5638,5639
0.9|5639,5642
SODIUM|5643,5649
-|5649,5650
140|5650,5653
<EOL>|5654,5655
POTASSIUM|5655,5664
-|5664,5665
4.2|5665,5668
CHLORIDE|5669,5677
-|5677,5678
103|5678,5681
TOTAL|5682,5687
CO2|5688,5691
-|5691,5692
29|5692,5694
ANION|5695,5700
GAP|5701,5704
-|5704,5705
12|5705,5707
<EOL>|5707,5708
_|5708,5709
_|5709,5710
_|5710,5711
03|5712,5714
:|5714,5715
58PM|5715,5719
estGFR|5722,5728
-|5728,5729
Using|5729,5734
this|5735,5739
<EOL>|5739,5740
_|5740,5741
_|5741,5742
_|5742,5743
03|5744,5746
:|5746,5747
58PM|5747,5751
TSH|5754,5757
-|5757,5758
1.4|5758,5761
<EOL>|5761,5762
_|5762,5763
_|5763,5764
_|5764,5765
03|5766,5768
:|5768,5769
58PM|5769,5773
ASA|5776,5779
-|5779,5780
NEG|5780,5783
ETHANOL|5784,5791
-|5791,5792
NEG|5792,5795
ACETMNPHN|5796,5805
-|5805,5806
NEG|5806,5809
<EOL>|5810,5811
bnzodzpn|5811,5819
-|5819,5820
NEG|5820,5823
barbitrt|5824,5832
-|5832,5833
NEG|5833,5836
tricyclic|5837,5846
-|5846,5847
NEG|5847,5850
<EOL>|5850,5851
_|5851,5852
_|5852,5853
_|5853,5854
03|5855,5857
:|5857,5858
58PM|5858,5862
URINE|5863,5868
HOURS|5870,5875
-|5875,5876
RANDOM|5876,5882
<EOL>|5882,5883
_|5883,5884
_|5884,5885
_|5885,5886
03|5887,5889
:|5889,5890
58PM|5890,5894
URINE|5895,5900
HOURS|5902,5907
-|5907,5908
RANDOM|5908,5914
<EOL>|5914,5915
_|5915,5916
_|5916,5917
_|5917,5918
03|5919,5921
:|5921,5922
58PM|5922,5926
URINE|5927,5932
GR|5934,5936
HOLD|5937,5941
-|5941,5942
HOLD|5942,5946
<EOL>|5946,5947
_|5947,5948
_|5948,5949
_|5949,5950
03|5951,5953
:|5953,5954
58PM|5954,5958
URINE|5959,5964
bnzodzpn|5966,5974
-|5974,5975
NEG|5975,5978
barbitrt|5979,5987
-|5987,5988
NEG|5988,5991
opiates|5992,5999
-|5999,6000
NEG|6000,6003
<EOL>|6004,6005
cocaine|6005,6012
-|6012,6013
NEG|6013,6016
amphetmn|6017,6025
-|6025,6026
NEG|6026,6029
mthdone|6030,6037
-|6037,6038
NEG|6038,6041
<EOL>|6041,6042
_|6042,6043
_|6043,6044
_|6044,6045
03|6046,6048
:|6048,6049
58PM|6049,6053
WBC|6056,6059
-|6059,6060
7.6|6060,6063
RBC|6064,6067
-|6067,6068
5|6068,6069
.|6069,6070
09|6070,6072
HGB|6073,6076
-|6076,6077
14.5|6077,6081
HCT|6082,6085
-|6085,6086
42.6|6086,6090
MCV|6091,6094
-|6094,6095
84|6095,6097
<EOL>|6098,6099
MCH|6099,6102
-|6102,6103
28.5|6103,6107
MCHC|6108,6112
-|6112,6113
34.0|6113,6117
RDW|6118,6121
-|6121,6122
12.7|6122,6126
<EOL>|6126,6127
_|6127,6128
_|6128,6129
_|6129,6130
03|6131,6133
:|6133,6134
58PM|6134,6138
NEUTS|6141,6146
-|6146,6147
55.6|6147,6151
_|6152,6153
_|6153,6154
_|6154,6155
MONOS|6156,6161
-|6161,6162
3.7|6162,6165
EOS|6166,6169
-|6169,6170
1.4|6170,6173
<EOL>|6174,6175
BASOS|6175,6180
-|6180,6181
0.5|6181,6184
<EOL>|6184,6185
_|6185,6186
_|6186,6187
_|6187,6188
03|6189,6191
:|6191,6192
58PM|6192,6196
PLT|6199,6202
COUNT|6203,6208
-|6208,6209
287|6209,6212
<EOL>|6212,6213
_|6213,6214
_|6214,6215
_|6215,6216
03|6217,6219
:|6219,6220
58PM|6220,6224
URINE|6225,6230
COLOR|6232,6237
-|6237,6238
Yellow|6238,6244
APPEAR|6245,6251
-|6251,6252
Clear|6252,6257
SP|6258,6260
_|6261,6262
_|6262,6263
_|6263,6264
<EOL>|6264,6265
_|6265,6266
_|6266,6267
_|6267,6268
03|6269,6271
:|6271,6272
58PM|6272,6276
URINE|6277,6282
BLOOD|6284,6289
-|6289,6290
NEG|6290,6293
NITRITE|6294,6301
-|6301,6302
NEG|6302,6305
PROTEIN|6306,6313
-|6313,6314
NEG|6314,6317
<EOL>|6318,6319
GLUCOSE|6319,6326
-|6326,6327
NEG|6327,6330
KETONE|6331,6337
-|6337,6338
NEG|6338,6341
BILIRUBIN|6342,6351
-|6351,6352
NEG|6352,6355
UROBILNGN|6356,6365
-|6365,6366
NEG|6366,6369
PH|6370,6372
-|6372,6373
6.5|6373,6376
<EOL>|6377,6378
LEUK|6378,6382
-|6382,6383
NEG|6383,6386
<EOL>|6386,6387
<EOL>|6388,6389
Brief|6389,6394
Hospital|6395,6403
Course|6404,6410
:|6410,6411
<EOL>|6411,6412
1|6412,6413
)|6413,6414
Psychiatric|6415,6426
:|6426,6427
<EOL>|6427,6428
Pt|6428,6430
arrived|6431,6438
on|6439,6441
floor|6442,6447
denying|6448,6455
passive|6456,6463
abd|6464,6467
active|6468,6474
SI|6475,6477
,|6477,6478
intent|6479,6485
,|6485,6486
plan|6487,6491
<EOL>|6492,6493
but|6493,6496
admitted|6497,6505
to|6506,6508
still|6509,6514
feeling|6515,6522
depressed|6523,6532
,|6532,6533
anxious|6534,6541
.|6541,6542
he|6543,6545
was|6546,6549
eager|6550,6555
<EOL>|6556,6557
to|6557,6559
start|6560,6565
treatment|6566,6575
and|6576,6579
meds|6580,6584
.|6584,6585
Consequently|6586,6598
,|6598,6599
celexa|6600,6606
10|6607,6609
mg|6610,6612
and|6613,6616
<EOL>|6617,6618
klonopin|6618,6626
0.5|6627,6630
QHS|6631,6634
and|6635,6638
0.5|6639,6642
BID|6643,6646
prns|6647,6651
anxiety|6652,6659
were|6660,6664
started|6665,6672
.|6672,6673
No|6674,6676
side|6677,6681
<EOL>|6682,6683
effects|6683,6690
,|6690,6691
pt|6692,6694
reported|6695,6703
significant|6704,6715
anxiety|6716,6723
reduction|6724,6733
and|6734,6737
<EOL>|6738,6739
resolution|6739,6749
of|6750,6752
depressive|6753,6763
symptoms|6764,6772
(|6773,6774
slept|6774,6779
throughout|6780,6790
the|6791,6794
night|6795,6800
)|6800,6801
<EOL>|6802,6803
and|6803,6806
all|6807,6810
SI|6811,6813
/|6813,6814
SIB|6814,6817
urges|6818,6823
within|6824,6830
days|6831,6835
of|6836,6838
arrival|6839,6846
.|6846,6847
He|6848,6850
stated|6851,6857
he|6858,6860
<EOL>|6861,6862
realized|6862,6870
he|6871,6873
had|6874,6877
overreacted|6878,6889
in|6890,6892
his|6893,6896
dealings|6897,6905
with|6906,6910
the|6911,6914
teacher|6915,6922
and|6923,6926
<EOL>|6927,6928
wanted|6928,6934
to|6935,6937
be|6938,6940
discharged|6941,6951
so|6952,6954
that|6955,6959
he|6960,6962
could|6963,6968
return|6969,6975
to|6976,6978
school|6979,6985
.|6985,6986
<EOL>|6987,6988
However|6988,6995
,|6995,6996
in|6997,6999
speaking|7000,7008
with|7009,7013
_|7014,7015
_|7015,7016
_|7016,7017
(|7018,7019
counselor|7019,7028
at|7029,7031
_|7032,7033
_|7033,7034
_|7034,7035
)|7035,7036
<EOL>|7037,7038
_|7038,7039
_|7039,7040
_|7040,7041
and|7042,7045
the|7046,7049
Academic|7050,7058
_|7059,7060
_|7060,7061
_|7061,7062
@|7063,7064
_|7064,7065
_|7065,7066
_|7066,7067
,|7067,7068
_|7069,7070
_|7070,7071
_|7071,7072
<EOL>|7073,7074
_|7074,7075
_|7075,7076
_|7076,7077
,|7077,7078
both|7079,7083
expressed|7084,7093
concerns|7094,7102
over|7103,7107
pt|7108,7110
's|7110,7112
"|7113,7114
repeated|7114,7122
<EOL>|7122,7123
acts|7123,7127
of|7128,7130
impulsivity|7131,7142
(|7143,7144
apparently|7144,7154
in|7155,7157
_|7158,7159
_|7159,7160
_|7160,7161
he|7162,7164
got|7165,7168
in|7169,7171
a|7172,7173
fight|7174,7179
<EOL>|7180,7181
with|7181,7185
another|7186,7193
student|7194,7201
who|7202,7205
he|7206,7208
thought|7209,7216
was|7217,7220
talking|7221,7228
about|7229,7234
him|7235,7238
.|7238,7239
He|7240,7242
<EOL>|7243,7244
then|7244,7248
ran|7249,7252
back|7253,7257
to|7258,7260
his|7261,7264
roomatte|7265,7273
's|7273,7275
dorm|7276,7280
and|7281,7284
asked|7285,7290
the|7291,7294
roommate|7295,7303
to|7304,7306
<EOL>|7307,7308
kill|7308,7312
hm|7313,7315
by|7316,7318
cutting|7319,7326
his|7327,7330
throat|7331,7337
)|7337,7338
.|7338,7339
They|7340,7344
both|7345,7349
stated|7350,7356
the|7357,7360
pt|7361,7363
had|7364,7367
<EOL>|7368,7369
"|7369,7370
burned|7370,7376
a|7377,7378
lot|7379,7382
more|7383,7387
bridges|7388,7395
"|7395,7396
than|7397,7401
just|7402,7406
the|7407,7410
one|7411,7414
teacher|7415,7422
he|7423,7425
had|7426,7429
a|7430,7431
<EOL>|7432,7433
falling|7433,7440
out|7441,7444
<EOL>|7444,7445
with|7445,7449
,|7449,7450
that|7451,7455
other|7456,7461
teachers|7462,7470
at|7471,7473
_|7474,7475
_|7475,7476
_|7476,7477
are|7478,7481
still|7482,7487
"|7488,7489
unwilling|7489,7498
or|7499,7501
<EOL>|7502,7503
concerned|7503,7512
to|7513,7515
take|7516,7520
him|7521,7524
on|7525,7527
as|7528,7530
a|7531,7532
student|7533,7540
given|7541,7546
his|7547,7550
growing|7551,7558
<EOL>|7559,7560
reputation|7560,7570
as|7571,7573
impulsive|7574,7583
"|7583,7584
.|7584,7585
They|7586,7590
stated|7591,7597
the|7598,7601
NEC|7602,7605
may|7606,7609
<EOL>|7609,7610
recommend|7610,7619
pt|7620,7622
take|7623,7627
the|7628,7631
rest|7632,7636
of|7637,7639
the|7640,7643
semester|7644,7652
off|7653,7656
on|7657,7659
medical|7660,7667
leave|7668,7673
.|7673,7674
<EOL>|7675,7676
<EOL>|7676,7677
<EOL>|7677,7678
We|7678,7680
had|7681,7684
a|7685,7686
meeting|7687,7694
with|7695,7699
team|7700,7704
,|7704,7705
the|7706,7709
academic|7710,7718
_|7719,7720
_|7720,7721
_|7721,7722
of|7723,7725
_|7726,7727
_|7727,7728
_|7728,7729
,|7729,7730
and|7731,7734
the|7735,7738
<EOL>|7739,7740
patient|7740,7747
where|7748,7753
all|7754,7757
parties|7758,7765
agreed|7766,7772
that|7773,7777
the|7778,7781
pt|7782,7784
should|7785,7791
take|7792,7796
the|7797,7800
<EOL>|7801,7802
rest|7802,7806
of|7807,7809
the|7810,7813
semester|7814,7822
off|7823,7826
on|7827,7829
medical|7830,7837
leave|7838,7843
of|7844,7846
absence|7847,7854
with|7855,7859
the|7860,7863
<EOL>|7864,7865
possibility|7865,7876
of|7877,7879
returning|7880,7889
next|7890,7894
year|7895,7899
.|7899,7900
The|7901,7904
patient|7905,7912
stated|7913,7919
,|7919,7920
after|7921,7926
<EOL>|7927,7928
speaking|7928,7936
with|7937,7941
his|7942,7945
family|7946,7952
,|7952,7953
that|7954,7958
he|7959,7961
would|7962,7967
return|7968,7974
to|7975,7977
_|7978,7979
_|7979,7980
_|7980,7981
<EOL>|7982,7983
_|7983,7984
_|7984,7985
_|7985,7986
immediately|7987,7998
to|7999,8001
be|8002,8004
close|8005,8010
to|8011,8013
his|8014,8017
family|8018,8024
,|8024,8025
"|8026,8027
for|8027,8030
extra|8031,8036
support|8037,8044
"|8044,8045
<EOL>|8046,8047
during|8047,8053
his|8054,8057
time|8058,8062
of|8063,8065
medical|8066,8073
leave.|8074,8080
he|8081,8083
strongly|8084,8092
agreed|8093,8099
that|8100,8104
he|8105,8107
<EOL>|8108,8109
needed|8109,8115
to|8116,8118
continue|8119,8127
taking|8128,8134
his|8135,8138
medications|8139,8150
and|8151,8154
would|8155,8160
followup|8161,8169
<EOL>|8170,8171
with|8171,8175
psychiatric|8176,8187
care|8188,8192
arranged|8193,8201
in|8202,8204
_|8205,8206
_|8206,8207
_|8207,8208
for|8209,8212
him|8213,8216
.|8216,8217
The|8218,8221
school|8222,8228
<EOL>|8229,8230
was|8230,8233
satisfied|8234,8243
with|8244,8248
his|8249,8252
mental|8253,8259
status|8260,8266
at|8267,8269
this|8270,8274
joint|8275,8280
meeting|8281,8288
and|8289,8292
<EOL>|8293,8294
felt|8294,8298
he|8299,8301
was|8302,8305
safe|8306,8310
to|8311,8313
be|8314,8316
discharged.|8317,8328
Pt|8329,8331
continued|8332,8341
to|8342,8344
deny|8345,8349
<EOL>|8350,8351
depression|8351,8361
,|8361,8362
SI|8363,8365
,|8365,8366
SIB|8367,8370
,|8370,8371
was|8372,8375
future|8376,8382
oriented|8383,8391
and|8392,8395
goal|8396,8400
oriented|8401,8409
and|8410,8413
<EOL>|8414,8415
was|8415,8418
deemed|8419,8425
safe|8426,8430
for|8431,8434
discharge|8435,8444
on|8445,8447
_|8448,8449
_|8449,8450
_|8450,8451
.|8451,8452
<EOL>|8452,8453
<EOL>|8453,8454
2|8454,8455
)|8455,8456
Medical|8457,8464
:|8464,8465
<EOL>|8465,8466
No|8466,8468
active|8469,8475
issues|8476,8482
during|8483,8489
hospital|8490,8498
stay|8499,8503
.|8503,8504
<EOL>|8504,8505
<EOL>|8505,8506
3|8506,8507
)|8507,8508
Groups|8509,8515
/|8515,8516
Behavioral|8516,8526
:|8526,8527
<EOL>|8527,8528
Pt|8528,8530
attended|8531,8539
groups|8540,8546
,|8546,8547
remained|8548,8556
visible|8557,8564
and|8565,8568
calm|8570,8574
in|8575,8577
unit|8578,8582
milieu|8583,8589
.|8589,8590
<EOL>|8592,8593
no|8593,8595
disruptive|8596,8606
or|8607,8609
threatening|8610,8621
behavior|8622,8630
.|8630,8631
no|8633,8635
quiet|8636,8641
room|8642,8646
,|8646,8647
1|8648,8649
:|8649,8650
1|8650,8651
<EOL>|8652,8653
sitter|8653,8659
,|8659,8660
physical|8661,8669
or|8670,8672
chemical|8673,8681
restraints|8682,8692
needed|8693,8699
at|8700,8702
any|8703,8706
time|8707,8711
.|8711,8712
<EOL>|8712,8713
<EOL>|8713,8714
4|8714,8715
)|8715,8716
Legal|8717,8722
:|8722,8723
<EOL>|8723,8724
_|8724,8725
_|8725,8726
_|8726,8727
<EOL>|8727,8728
Medications|8728,8739
on|8740,8742
Admission|8743,8752
:|8752,8753
<EOL>|8753,8754
none|8754,8758
<EOL>|8758,8759
<EOL>|8760,8761
Discharge|8761,8770
Medications|8771,8782
:|8782,8783
<EOL>|8783,8784
1.|8784,8786
Citalopram|8787,8797
20|8798,8800
mg|8801,8803
Tablet|8804,8810
Sig|8811,8814
:|8814,8815
One|8816,8819
(|8820,8821
1|8821,8822
)|8822,8823
Tablet|8824,8830
PO|8831,8833
DAILY|8834,8839
(|8840,8841
Daily|8841,8846
)|8846,8847
.|8847,8848
<EOL>|8848,8849
Disp|8849,8853
:|8853,8854
*|8854,8855
30|8855,8857
Tablet|8858,8864
(|8864,8865
s|8865,8866
)|8866,8867
*|8867,8868
Refills|8869,8876
:|8876,8877
*|8877,8878
0|8878,8879
*|8879,8880
<EOL>|8880,8881
2.|8881,8883
Clonazepam|8884,8894
0.5|8895,8898
mg|8899,8901
Tablet|8902,8908
Sig|8909,8912
:|8912,8913
One|8914,8917
(|8918,8919
1|8919,8920
)|8920,8921
Tablet|8922,8928
PO|8929,8931
QAM|8932,8935
and|8936,8939
QHS|8940,8943
.|8943,8944
<EOL>|8944,8945
Disp|8945,8949
:|8949,8950
*|8950,8951
12|8951,8953
Tablet|8954,8960
(|8960,8961
s|8961,8962
)|8962,8963
*|8963,8964
Refills|8965,8972
:|8972,8973
*|8973,8974
0|8974,8975
*|8975,8976
<EOL>|8976,8977
<EOL>|8977,8978
<EOL>|8979,8980
Discharge|8980,8989
Disposition|8990,9001
:|9001,9002
<EOL>|9002,9003
Home|9003,9007
<EOL>|9007,9008
<EOL>|9009,9010
Discharge|9010,9019
Diagnosis|9020,9029
:|9029,9030
<EOL>|9030,9031
Axis|9031,9035
I|9036,9037
:|9037,9038
<EOL>|9038,9039
Major|9039,9044
depressive|9045,9055
disorder|9056,9064
,|9064,9065
severe|9066,9072
,|9072,9073
without|9074,9081
psychotic|9082,9091
features|9092,9100
<EOL>|9100,9101
Anxiety|9101,9108
disorder|9109,9117
not|9118,9121
otherwise|9122,9131
specified|9132,9141
<EOL>|9141,9142
II|9142,9144
-|9144,9145
deferred|9146,9154
<EOL>|9154,9155
III|9155,9158
-|9158,9159
status|9160,9166
post|9167,9171
meniscus|9172,9180
repair|9181,9187
(|9188,9189
knee|9189,9193
)|9193,9194
<EOL>|9194,9195
IV|9195,9197
-|9197,9198
moderately|9199,9209
severe|9210,9216
psychosocial|9217,9229
stressors|9230,9239
identified|9240,9250
<EOL>|9250,9251
V|9251,9252
-|9252,9253
GAF|9254,9257
upon|9258,9262
discharge|9263,9272
:|9272,9273
45|9274,9276
<EOL>|9276,9277
<EOL>|9277,9278
<EOL>|9279,9280
Discharge|9280,9289
Condition|9290,9299
:|9299,9300
<EOL>|9300,9301
MSE|9301,9304
:|9304,9305
general|9305,9312
-|9312,9313
thin|9314,9318
caucasian|9319,9328
man|9329,9332
,|9332,9333
seated|9333,9339
,|9339,9340
NAD|9341,9344
<EOL>|9344,9345
behavior|9345,9353
=|9353,9354
calm|9355,9359
,|9359,9360
no|9361,9363
tremors|9364,9371
,|9371,9372
no|9373,9375
PMA|9376,9379
<EOL>|9379,9380
speech|9380,9386
-|9386,9387
normal|9388,9394
,|9394,9395
not|9396,9399
pressured|9400,9409
<EOL>|9410,9411
affect|9411,9417
:|9417,9418
more|9420,9424
emotionally|9425,9436
reactive|9437,9445
than|9446,9450
<EOL>|9450,9451
prior|9451,9456
,|9456,9457
smiles|9458,9464
appropriately|9465,9478
,|9478,9479
even|9480,9484
and|9485,9488
euthymic|9489,9497
<EOL>|9497,9498
TC|9498,9500
:|9500,9501
no|9502,9504
delusions|9505,9514
,|9514,9515
no|9516,9518
AVH|9519,9522
<EOL>|9522,9523
TP|9523,9525
:|9525,9526
linear|9527,9533
and|9534,9537
goal|9538,9542
-|9542,9543
directed|9543,9551
;|9551,9552
<EOL>|9552,9553
safety|9553,9559
-|9559,9560
denies|9561,9567
SI|9568,9570
,|9570,9571
SIB|9572,9575
,|9575,9576
intent|9577,9583
,|9583,9584
plan|9585,9589
<EOL>|9590,9591
cog|9591,9594
:|9594,9595
AOx3|9596,9600
<EOL>|9600,9601
I|9601,9602
/|9602,9603
J|9603,9604
;|9604,9605
fair|9606,9610
/|9610,9611
fair|9611,9615
<EOL>|9615,9616
<EOL>|9616,9617
<EOL>|9618,9619
Discharge|9619,9628
Instructions|9629,9641
:|9641,9642
<EOL>|9642,9643
Please|9643,9649
take|9650,9654
medications|9655,9666
as|9667,9669
prescribed|9670,9680
.|9680,9681
<EOL>|9681,9682
Please|9682,9688
attend|9689,9695
outpatient|9696,9706
appointments|9707,9719
as|9720,9722
scheduled|9723,9732
.|9732,9733
<EOL>|9733,9734
If|9734,9736
you|9737,9740
are|9741,9744
feeling|9745,9752
unsafe|9753,9759
or|9760,9762
that|9763,9767
your|9768,9772
condition|9773,9782
is|9783,9785
worsening|9786,9795
,|9795,9796
<EOL>|9797,9798
call|9798,9802
_|9803,9804
_|9804,9805
_|9805,9806
or|9807,9809
go|9810,9812
to|9813,9815
your|9816,9820
nearest|9821,9828
ED|9829,9831
<EOL>|9831,9832
<EOL>|9832,9833
<EOL>|9834,9835
Followup|9835,9843
Instructions|9844,9856
:|9856,9857
<EOL>|9857,9858
_|9858,9859
_|9859,9860
_|9860,9861
<EOL>|9861,9862

