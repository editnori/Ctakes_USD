 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|25,29
No|30,32
:|32,33
_|36,37
_|37,38
_|38,39
<EOL>|39,40
<EOL>|41,42
Admission|42,51
Date|52,56
:|56,57
_|59,60
_|60,61
_|61,62
Discharge|76,85
Date|86,90
:|90,91
_|94,95
_|95,96
_|96,97
<EOL>|97,98
<EOL>|99,100
Date|100,104
of|105,107
Birth|108,113
:|113,114
_|116,117
_|117,118
_|118,119
Sex|132,135
:|135,136
F|139,140
<EOL>|140,141
<EOL>|142,143
Service|143,150
:|150,151
MEDICINE|152,160
<EOL>|160,161
<EOL>|162,163
No|175,177
Known|178,183
Allergies|184,193
/|194,195
Adverse|196,203
Drug|204,208
Reactions|209,218
<EOL>|218,219
<EOL>|220,221
Attending|221,230
:|230,231
_|232,233
_|233,234
_|234,235
.|235,236
<EOL>|236,237
<EOL>|238,239
Fever|256,261
,|261,262
non-productive|263,277
cough|278,283
<EOL>|283,284
<EOL>|285,286
Major|286,291
Surgical|292,300
or|301,303
Invasive|304,312
Procedure|313,322
:|322,323
<EOL>|323,324
None|324,328
<EOL>|328,329
<EOL>|329,330
<EOL>|331,332
_|360,361
_|361,362
_|362,363
yo|364,366
F|367,368
w|369,370
/|370,371
HTN|372,375
,|375,376
CAD|377,380
,|380,381
COPD|382,386
p|387,388
/|388,389
w|389,390
fevers|391,397
,|397,398
non-productive|399,413
cough|414,419
,|419,420
<EOL>|421,422
since|422,427
_|428,429
_|429,430
_|430,431
.|431,432
Pt|433,435
said|436,440
she|441,444
was|445,448
in|449,451
her|452,455
usual|456,461
state|462,467
of|468,470
health|471,477
until|478,483
<EOL>|484,485
_|485,486
_|486,487
_|487,488
evening|489,496
when|497,501
she|502,505
developed|506,515
a|516,517
cough|518,523
producing|524,533
_|534,535
_|535,536
_|536,537
<EOL>|538,539
sputum|539,545
.|545,546
She|548,551
took|552,556
some|557,561
robitussin|562,572
and|573,576
went|577,581
to|582,584
bed|585,588
.|588,589
She|591,594
woke|595,599
up|600,602
<EOL>|603,604
the|604,607
next|608,612
morning|613,620
and|621,624
had|625,628
general|629,636
malaise|637,644
,|644,645
nasal|646,651
congestion|652,662
,|662,663
<EOL>|664,665
intermittently|665,679
productive|680,690
cough|691,696
.|696,697
She|699,702
did|703,706
not|707,710
want|711,715
to|716,718
eat|719,722
and|723,726
<EOL>|727,728
had|728,731
4|732,733
episodes|734,742
of|743,745
water|746,751
diarrhea|752,760
and|761,764
one|765,768
episode|769,776
of|777,779
vomiting|780,788
<EOL>|789,790
without|790,797
nausea|798,804
.|804,805
She|807,810
denied|811,817
fevers|818,824
,|824,825
chills|826,832
or|833,835
sweats|836,842
at|843,845
that|846,850
<EOL>|851,852
time|852,856
.|856,857
She|859,862
called|863,869
her|870,873
PCP|874,877
who|878,881
prescribed|882,892
_|893,894
_|894,895
_|895,896
Z|897,898
-|898,899
pack|899,903
.|903,904
Her|906,909
symptoms|910,918
<EOL>|919,920
persisted|920,929
and|930,933
she|934,937
developed|938,947
pain|948,952
with|953,957
coughing|958,966
around|967,973
her|974,977
upper|978,983
<EOL>|984,985
abdomen|985,992
and|993,996
lower|997,1002
chest|1003,1008
.|1008,1009
Denies|1011,1017
other|1018,1023
joint|1024,1029
or|1030,1032
muscle|1033,1039
pain|1040,1044
.|1044,1045
<EOL>|1047,1048
She|1048,1051
went|1052,1056
to|1057,1059
see|1060,1063
her|1064,1067
PCP|1068,1071
on|1072,1074
the|1075,1078
day|1079,1082
of|1083,1085
admission|1086,1095
.|1095,1096
In|1098,1100
her|1101,1104
PCP|1105,1108
's|1108,1110
<EOL>|1111,1112
office|1112,1118
was|1119,1122
hypoxic|1123,1130
on|1131,1133
RA|1134,1136
,|1136,1137
here|1138,1142
is|1143,1145
89|1146,1148
%|1148,1149
on|1150,1152
RA|1153,1155
.|1155,1156
Has|1157,1160
had|1161,1164
flu|1165,1168
vaccine|1169,1176
<EOL>|1177,1178
this|1178,1182
year|1183,1187
and|1188,1191
pneumovax|1192,1201
last|1202,1206
year|1207,1211
.|1211,1212
wheezy|1213,1219
on|1220,1222
exam|1223,1227
,|1227,1228
on|1229,1231
2L|1232,1234
with|1235,1239
o2|1240,1242
<EOL>|1243,1244
sat|1244,1247
mid-90s|1248,1255
.|1255,1256
<EOL>|1258,1259
.|1259,1260
<EOL>|1260,1261
In|1261,1263
ED|1264,1266
VS|1267,1269
were|1270,1274
afebrile|1275,1283
70|1284,1286
113|1287,1290
/|1290,1291
66|1291,1293
94|1294,1296
%|1296,1297
2L|1297,1299
,|1299,1300
On|1301,1303
exam|1304,1308
had|1309,1312
wheezes|1313,1320
with|1321,1325
<EOL>|1326,1327
peak|1327,1331
flow|1332,1336
of|1337,1339
150|1340,1343
(|1344,1345
no|1345,1347
baseline|1348,1356
)|1356,1357
,|1357,1358
speaking|1359,1367
in|1368,1370
full|1371,1375
sentences|1376,1385
and|1386,1389
<EOL>|1390,1391
no|1391,1393
accessory|1394,1403
muscle|1404,1410
use|1411,1414
,|1414,1415
euvolemic|1416,1425
and|1426,1429
no|1430,1432
_|1433,1434
_|1434,1435
_|1435,1436
edema|1437,1442
.|1442,1443
Flu|1445,1448
screen|1449,1455
<EOL>|1456,1457
not|1457,1460
performed|1461,1470
,|1470,1471
CXR|1472,1475
unremarkable|1476,1488
compared|1489,1497
to|1498,1500
prior|1501,1506
.|1506,1507
Given|1509,1514
<EOL>|1515,1516
levoflox|1516,1524
,|1524,1525
nebs|1526,1530
,|1530,1531
pred|1532,1536
50|1537,1539
mg|1540,1542
.|1542,1543
<EOL>|1543,1544
<EOL>|1544,1545
<EOL>|1546,1547
ASTHMA|1569,1575
<EOL>|1578,1579
HYPERTENSION|1579,1591
<EOL>|1594,1595
HYPERLIPIDEMIA|1595,1609
<EOL>|1612,1613
HEADACHE|1613,1621
<EOL>|1624,1625
OSTEOARTHRITIS|1625,1639
<EOL>|1642,1643
ATYPICAL|1643,1651
CHEST|1652,1657
PAIN|1658,1662
<EOL>|1665,1666
TOBACCO|1666,1673
ABUSE|1674,1679
<EOL>|1682,1683
ABNORMAL|1683,1691
CHEST|1692,1697
XRAY|1698,1702
<EOL>|1705,1706
COPD|1706,1710
<EOL>|1712,1713
<EOL>|1714,1715
:|1729,1730
<EOL>|1730,1731
_|1731,1732
_|1732,1733
_|1733,1734
<EOL>|1734,1735
:|1749,1750
<EOL>|1750,1751
Mother|1751,1757
:|1757,1758
_|1759,1760
_|1760,1761
_|1761,1762
,|1762,1763
HTN|1764,1767
<EOL>|1769,1770
Father|1770,1776
:|1776,1777
_|1778,1779
_|1779,1780
_|1780,1781
CA|1782,1784
<EOL>|1786,1787
Brother|1787,1794
:|1794,1795
CA|1796,1798
?|1798,1799
<EOL>|1801,1802
Brother|1802,1809
:|1809,1810
_|1811,1812
_|1812,1813
_|1813,1814
<EOL>|1816,1817
<EOL>|1817,1818
<EOL>|1819,1820
Physical|1820,1828
_|1829,1830
_|1830,1831
_|1831,1832
:|1832,1833
<EOL>|1833,1834
On|1834,1836
Admission|1837,1846
:|1846,1847
<EOL>|1847,1848
VS|1848,1850
:|1850,1851
T|1852,1853
:|1853,1854
,|1856,1857
BP|1858,1860
:|1860,1861
142|1862,1865
/|1865,1866
70|1866,1868
,|1868,1869
HR|1870,1872
:|1872,1873
70|1874,1876
,|1876,1877
RR|1878,1880
20|1881,1883
,|1883,1884
O2|1885,1887
93|1888,1890
%|1890,1891
on|1892,1894
RA|1895,1897
(|1898,1899
96|1899,1901
%|1901,1902
2L|1903,1905
)|1905,1906
<EOL>|1906,1907
GA|1907,1909
:|1909,1910
AOx3|1911,1915
,|1915,1916
pt|1917,1919
with|1920,1924
nasal|1925,1930
cannula|1931,1938
on|1939,1941
in|1942,1944
no|1945,1947
respiratory|1948,1959
distress|1960,1968
<EOL>|1968,1969
HEENT|1969,1974
:|1974,1975
MMM|1977,1980
.|1980,1981
no|1982,1984
LAD|1985,1988
.|1988,1989
no|1990,1992
JVD|1993,1996
.|1996,1997
neck|1998,2002
supple|2003,2009
.|2009,2010
<EOL>|2011,2012
Cards|2012,2017
:|2017,2018
RRR|2019,2022
S1|2023,2025
/|2025,2026
S2|2026,2028
heard|2029,2034
.|2034,2035
no|2036,2038
murmurs|2039,2046
/|2046,2047
gallops|2047,2054
/|2054,2055
rubs|2055,2059
.|2059,2060
<EOL>|2060,2061
Pulm|2061,2065
:|2065,2066
CTAB|2067,2071
no|2072,2074
crackles|2075,2083
or|2084,2086
wheezes|2087,2094
,|2094,2095
good|2096,2100
inspiratory|2101,2112
effort|2113,2119
,|2119,2120
but|2121,2124
<EOL>|2125,2126
not|2126,2129
great|2130,2135
air|2136,2139
movement|2140,2148
,|2148,2149
slightly|2150,2158
prolonged|2159,2168
expiratory|2169,2179
phase|2180,2185
.|2185,2186
<EOL>|2186,2187
Abd|2187,2190
:|2190,2191
soft|2192,2196
,|2196,2197
NT|2198,2200
,|2200,2201
+|2202,2203
BS|2203,2205
.|2205,2206
no|2207,2209
g|2210,2211
/|2211,2212
rt|2212,2214
.|2214,2215
neg|2216,2219
HSM|2220,2223
.|2223,2224
<EOL>|2224,2225
Extremities|2225,2236
:|2236,2237
wwp|2238,2241
,|2241,2242
no|2243,2245
edema|2246,2251
.|2251,2252
DPs|2253,2256
,|2256,2257
PTs|2258,2261
2|2262,2263
+|2263,2264
.|2264,2265
<EOL>|2265,2266
Skin|2266,2270
:|2270,2271
no|2272,2274
noticeable|2275,2285
rashes|2286,2292
<EOL>|2292,2293
Neuro|2293,2298
/|2298,2299
Psych|2299,2304
:|2304,2305
CNs|2306,2309
II|2310,2312
-|2312,2313
XII|2313,2316
intact|2317,2323
<EOL>|2323,2324
.|2324,2325
<EOL>|2325,2326
ON|2326,2328
DISCHARGE|2329,2338
:|2338,2339
<EOL>|2339,2340
VS|2340,2342
:|2342,2343
T|2344,2345
:|2345,2346
,|2348,2349
BP|2350,2352
:|2352,2353
142|2354,2357
/|2357,2358
70|2358,2360
,|2360,2361
HR|2362,2364
:|2364,2365
70|2366,2368
,|2368,2369
RR|2370,2372
20|2373,2375
,|2375,2376
O2|2377,2379
93|2380,2382
%|2382,2383
on|2384,2386
RA|2387,2389
(|2390,2391
96|2391,2393
%|2393,2394
2L|2395,2397
)|2397,2398
<EOL>|2398,2399
GA|2399,2401
:|2401,2402
AOx3|2403,2407
,|2407,2408
pt|2409,2411
with|2412,2416
nasal|2417,2422
cannula|2423,2430
on|2431,2433
in|2434,2436
no|2437,2439
respiratory|2440,2451
distress|2452,2460
<EOL>|2460,2461
HEENT|2461,2466
:|2466,2467
MMM|2469,2472
.|2472,2473
no|2474,2476
LAD|2477,2480
.|2480,2481
no|2482,2484
JVD|2485,2488
.|2488,2489
neck|2490,2494
supple|2495,2501
.|2501,2502
<EOL>|2503,2504
Cards|2504,2509
:|2509,2510
RRR|2511,2514
S1|2515,2517
/|2517,2518
S2|2518,2520
heard|2521,2526
.|2526,2527
no|2528,2530
murmurs|2531,2538
/|2538,2539
gallops|2539,2546
/|2546,2547
rubs|2547,2551
.|2551,2552
<EOL>|2552,2553
Pulm|2553,2557
:|2557,2558
CTAB|2559,2563
no|2564,2566
crackles|2567,2575
or|2576,2578
wheezes|2579,2586
,|2586,2587
good|2588,2592
inspiratory|2593,2604
effort|2605,2611
,|2611,2612
but|2613,2616
<EOL>|2617,2618
not|2618,2621
great|2622,2627
air|2628,2631
movement|2632,2640
,|2640,2641
slightly|2642,2650
prolonged|2651,2660
expiratory|2661,2671
phase|2672,2677
.|2677,2678
<EOL>|2678,2679
Abd|2679,2682
:|2682,2683
soft|2684,2688
,|2688,2689
NT|2690,2692
,|2692,2693
+|2694,2695
BS|2695,2697
.|2697,2698
no|2699,2701
g|2702,2703
/|2703,2704
rt|2704,2706
.|2706,2707
neg|2708,2711
HSM|2712,2715
.|2715,2716
<EOL>|2716,2717
Extremities|2717,2728
:|2728,2729
wwp|2730,2733
,|2733,2734
no|2735,2737
edema|2738,2743
.|2743,2744
DPs|2745,2748
,|2748,2749
PTs|2750,2753
2|2754,2755
+|2755,2756
.|2756,2757
<EOL>|2757,2758
Skin|2758,2762
:|2762,2763
no|2764,2766
noticeable|2767,2777
rashes|2778,2784
<EOL>|2784,2785
Neuro|2785,2790
/|2790,2791
Psych|2791,2796
:|2796,2797
CNs|2798,2801
II|2802,2804
-|2804,2805
XII|2805,2808
intact|2809,2815
<EOL>|2815,2816
<EOL>|2817,2818
Pertinent|2818,2827
Results|2828,2835
:|2835,2836
<EOL>|2836,2837
LABS|2837,2841
:|2841,2842
<EOL>|2842,2843
_|2843,2844
_|2844,2845
_|2845,2846
03|2847,2849
:|2849,2850
26PM|2850,2854
BLOOD|2855,2860
WBC|2861,2864
-|2864,2865
4.9|2865,2868
RBC|2869,2872
-|2872,2873
4.25|2873,2877
Hgb|2878,2881
-|2881,2882
12.7|2882,2886
Hct|2887,2890
-|2890,2891
36.5|2891,2895
MCV|2896,2899
-|2899,2900
86|2900,2902
<EOL>|2903,2904
MCH|2904,2907
-|2907,2908
30.0|2908,2912
MCHC|2913,2917
-|2917,2918
34.9|2918,2922
RDW|2923,2926
-|2926,2927
15.3|2927,2931
Plt|2932,2935
_|2936,2937
_|2937,2938
_|2938,2939
<EOL>|2939,2940
_|2940,2941
_|2941,2942
_|2942,2943
06|2944,2946
:|2946,2947
50AM|2947,2951
BLOOD|2952,2957
WBC|2958,2961
-|2961,2962
8|2962,2963
.|2963,2964
2|2964,2965
#|2965,2966
RBC|2967,2970
-|2970,2971
4|2971,2972
.|2972,2973
03|2973,2975
*|2975,2976
Hgb|2977,2980
-|2980,2981
12.2|2981,2985
Hct|2986,2989
-|2989,2990
34|2990,2992
.|2992,2993
8|2993,2994
*|2994,2995
<EOL>|2996,2997
MCV|2997,3000
-|3000,3001
87|3001,3003
MCH|3004,3007
-|3007,3008
30.4|3008,3012
MCHC|3013,3017
-|3017,3018
35|3018,3020
.|3020,3021
1|3021,3022
*|3022,3023
RDW|3024,3027
-|3027,3028
15.3|3028,3032
Plt|3033,3036
_|3037,3038
_|3038,3039
_|3039,3040
<EOL>|3040,3041
_|3041,3042
_|3042,3043
_|3043,3044
03|3045,3047
:|3047,3048
26PM|3048,3052
BLOOD|3053,3058
Glucose|3059,3066
-|3066,3067
123|3067,3070
*|3070,3071
UreaN|3072,3077
-|3077,3078
14|3078,3080
Creat|3081,3086
-|3086,3087
0.9|3087,3090
Na|3091,3093
-|3093,3094
136|3094,3097
<EOL>|3098,3099
K|3099,3100
-|3100,3101
3.3|3101,3104
Cl|3105,3107
-|3107,3108
97|3108,3110
HCO3|3111,3115
-|3115,3116
31|3116,3118
AnGap|3119,3124
-|3124,3125
_|3125,3126
_|3126,3127
_|3127,3128
06|3129,3131
:|3131,3132
50AM|3132,3136
BLOOD|3137,3142
Glucose|3143,3150
-|3150,3151
95|3151,3153
UreaN|3154,3159
-|3159,3160
17|3160,3162
Creat|3163,3168
-|3168,3169
0.8|3169,3172
Na|3173,3175
-|3175,3176
139|3176,3179
<EOL>|3180,3181
K|3181,3182
-|3182,3183
3.5|3183,3186
Cl|3187,3189
-|3189,3190
98|3190,3192
HCO3|3193,3197
-|3197,3198
30|3198,3200
AnGap|3201,3206
-|3206,3207
15|3207,3209
<EOL>|3209,3210
.|3210,3211
<EOL>|3211,3212
MICRO|3212,3217
:|3217,3218
<EOL>|3218,3219
*|3223,3224
*|3224,3225
FINAL|3225,3230
REPORT|3231,3237
_|3238,3239
_|3239,3240
_|3240,3241
<EOL>|3241,3242
<EOL>|3242,3243
DIRECT|3246,3252
INFLUENZA|3253,3262
A|3263,3264
ANTIGEN|3265,3272
TEST|3273,3277
(|3278,3279
Final|3279,3284
_|3285,3286
_|3286,3287
_|3287,3288
:|3288,3289
<EOL>|3290,3291
POSITIVE|3297,3305
FOR|3306,3309
INFLUENZA|3310,3319
A|3320,3321
VIRAL|3322,3327
ANTIGEN|3328,3335
.|3335,3336
<EOL>|3337,3338
REPORTED|3347,3355
BY|3356,3358
PHONE|3359,3364
TO|3365,3367
_|3368,3369
_|3369,3370
_|3370,3371
AT|3372,3374
1153|3375,3379
_|3381,3382
_|3382,3383
_|3383,3384
.|3384,3385
<EOL>|3385,3386
.|3386,3387
<EOL>|3387,3388
IMAGING|3388,3395
:|3395,3396
<EOL>|3396,3397
CXR|3397,3400
_|3401,3402
_|3402,3403
_|3403,3404
:|3404,3405
<EOL>|3405,3406
1|3419,3420
.|3420,3421
No|3422,3424
acute|3425,3430
chest|3431,3436
pathology|3437,3446
with|3447,3451
stable|3452,3458
pleural|3459,3466
parenchymal|3467,3478
<EOL>|3479,3480
scar|3480,3484
.|3484,3485
<EOL>|3486,3487
2.|3487,3489
Flattening|3490,3500
of|3501,3503
the|3504,3507
hemidiaphragms|3508,3522
consistent|3523,3533
with|3534,3538
COPD|3539,3543
.|3543,3544
<EOL>|3545,3546
<EOL>|3546,3547
<EOL>|3548,3549
A|3572,3573
/|3573,3574
P|3574,3575
:|3575,3576
_|3577,3578
_|3578,3579
_|3579,3580
year|3581,3585
old|3586,3589
woman|3590,3595
with|3596,3600
recent|3601,3607
onset|3608,3613
of|3614,3616
fevers|3617,3623
,|3623,3624
productive|3625,3635
<EOL>|3636,3637
cough|3637,3642
and|3643,3646
costochondral|3647,3660
vs|3661,3663
.|3663,3664
pleuritic|3665,3674
pain|3675,3679
who|3680,3683
tested|3684,3690
positive|3691,3699
<EOL>|3700,3701
for|3701,3704
influenza|3705,3714
A|3715,3716
.|3716,3717
<EOL>|3717,3718
.|3718,3719
<EOL>|3719,3720
#|3720,3721
Fevers|3722,3728
,|3728,3729
malaise|3730,3737
,|3737,3738
cough|3739,3744
:|3744,3745
Pt|3746,3748
seemed|3749,3755
to|3756,3758
have|3759,3763
onset|3764,3769
of|3770,3772
symptoms|3773,3781
<EOL>|3782,3783
consistent|3783,3793
with|3794,3798
viral|3799,3804
infection|3805,3814
.|3814,3815
She|3817,3820
was|3821,3824
admitted|3825,3833
to|3834,3836
the|3837,3840
<EOL>|3841,3842
hospital|3842,3850
and|3851,3854
placed|3855,3861
on|3862,3864
droplet|3865,3872
precautions|3873,3884
because|3885,3892
there|3893,3898
was|3899,3902
<EOL>|3903,3904
concern|3904,3911
that|3912,3916
she|3917,3920
had|3921,3924
the|3925,3928
flu|3929,3932
.|3932,3933
She|3935,3938
was|3939,3942
empirically|3943,3954
started|3955,3962
on|3963,3965
<EOL>|3966,3967
Oseltamivir|3967,3978
75mg|3979,3983
PO|3984,3986
BID|3987,3990
.|3990,3991
nasopharyngeal|3993,4007
swab|4008,4012
was|4013,4016
positive|4017,4025
for|4026,4029
<EOL>|4030,4031
influenza|4031,4040
A.|4041,4043
She|4045,4048
was|4049,4052
continued|4053,4062
on|4063,4065
a|4066,4067
five|4068,4072
day|4073,4076
regiment|4077,4085
of|4086,4088
<EOL>|4089,4090
oseltamivir|4090,4101
for|4102,4105
her|4106,4109
flu|4110,4113
and|4114,4117
will|4118,4122
follow|4123,4129
up|4130,4132
with|4133,4137
Dr.|4138,4141
_|4142,4143
_|4143,4144
_|4144,4145
in|4146,4148
the|4149,4152
<EOL>|4153,4154
outpatient|4154,4164
setting|4165,4172
.|4172,4173
<EOL>|4173,4174
.|4174,4175
<EOL>|4175,4176
#|4176,4177
COPD|4178,4182
exacerbation|4183,4195
:|4195,4196
Pt|4198,4200
tested|4201,4207
positive|4208,4216
for|4217,4220
the|4221,4224
flu|4225,4228
,|4228,4229
but|4230,4233
seemed|4234,4240
<EOL>|4241,4242
to|4242,4244
also|4245,4249
be|4250,4252
having|4253,4259
a|4260,4261
COPD|4262,4266
exacerbation|4267,4279
with|4280,4284
worsening|4285,4294
dyspnea|4295,4302
and|4303,4306
<EOL>|4307,4308
sputum|4308,4314
production|4315,4325
.|4325,4326
She|4328,4331
was|4332,4335
started|4336,4343
on|4344,4346
prednisone|4347,4357
50mg|4358,4362
PO|4363,4365
Daily|4366,4371
,|4371,4372
<EOL>|4373,4374
Azithromycin|4374,4386
and|4387,4390
O2|4391,4393
via|4394,4397
nasal|4398,4403
cannula|4404,4411
.|4411,4412
Her|4414,4417
resting|4418,4425
O2|4426,4428
sat|4429,4432
was|4433,4436
<EOL>|4437,4438
initially|4438,4447
85|4448,4450
%|4450,4451
,|4451,4452
but|4453,4456
at|4457,4459
the|4460,4463
time|4464,4468
of|4469,4471
discharge|4472,4481
she|4482,4485
was|4486,4489
satting|4490,4497
96|4498,4500
%|4500,4501
<EOL>|4502,4503
on|4503,4505
RA|4506,4508
,|4508,4509
but|4510,4513
would|4514,4519
desaturate|4520,4530
to|4531,4533
84|4534,4536
%|4536,4537
after|4538,4543
walking|4544,4551
75|4552,4554
-|4554,4555
100feet|4555,4562
.|4562,4563
<EOL>|4565,4566
She|4566,4569
Was|4570,4573
given|4574,4579
a|4580,4581
5|4582,4583
day|4584,4587
course|4588,4594
of|4595,4597
azithromycin|4598,4610
,|4610,4611
5|4612,4613
days|4614,4618
of|4619,4621
<EOL>|4622,4623
prednisone|4623,4633
at|4634,4636
50mg|4637,4641
PO|4642,4644
Daily|4645,4650
and|4651,4654
then|4655,4659
a|4660,4661
week|4662,4666
long|4667,4671
taper|4672,4677
and|4678,4681
<EOL>|4682,4683
discharged|4683,4693
on|4694,4696
home|4697,4701
O2|4702,4704
while|4705,4710
her|4711,4714
symptoms|4715,4723
improved|4724,4732
.|4732,4733
The|4735,4738
patient|4739,4746
<EOL>|4747,4748
was|4748,4751
breathing|4752,4761
more|4762,4766
comfortably|4767,4778
and|4779,4782
ambulating|4783,4793
well|4794,4798
at|4799,4801
the|4802,4805
time|4806,4810
<EOL>|4811,4812
of|4812,4814
discharge|4815,4824
.|4824,4825
She|4827,4830
will|4831,4835
follow|4836,4842
up|4843,4845
with|4846,4850
Dr.|4851,4854
_|4855,4856
_|4856,4857
_|4857,4858
as|4859,4861
well|4862,4866
as|4867,4869
Dr|4870,4872
.|4872,4873
<EOL>|4874,4875
_|4875,4876
_|4876,4877
_|4877,4878
in|4879,4881
the|4882,4885
outpatient|4886,4896
setting|4897,4904
.|4904,4905
<EOL>|4905,4906
.|4906,4907
<EOL>|4907,4908
#|4908,4909
ASTHMA|4910,4916
:|4916,4917
pt|4918,4920
with|4921,4925
wheezing|4926,4934
in|4935,4937
the|4938,4941
ED|4942,4944
and|4945,4948
at|4949,4951
PCP|4952,4955
office|4956,4962
,|4962,4963
but|4964,4967
not|4968,4971
<EOL>|4972,4973
present|4973,4980
on|4981,4983
my|4984,4986
exams|4987,4992
,|4992,4993
however|4994,5001
,|5001,5002
she|5003,5006
had|5007,5010
received|5011,5019
duonebs|5020,5027
prior|5028,5033
to|5034,5036
<EOL>|5037,5038
my|5038,5040
exam|5041,5045
.|5045,5046
Likely|5048,5054
having|5055,5061
asthma|5062,5068
symptoms|5069,5077
in|5078,5080
setting|5081,5088
of|5089,5091
COPD|5092,5096
<EOL>|5097,5098
exacerbations|5098,5111
.|5111,5112
She|5114,5117
was|5118,5121
continued|5122,5131
on|5132,5134
her|5135,5138
home|5139,5143
regiment|5144,5152
and|5153,5156
also|5157,5161
<EOL>|5162,5163
on|5163,5165
standing|5166,5174
nebulizers|5175,5185
.|5185,5186
She|5188,5191
was|5192,5195
discharged|5196,5206
with|5207,5211
nebulizer|5212,5221
<EOL>|5222,5223
treamtents|5223,5233
as|5234,5236
well|5237,5241
as|5242,5244
her|5245,5248
home|5249,5253
medications|5254,5265
.|5265,5266
Respiratory|5268,5279
status|5280,5286
<EOL>|5287,5288
was|5288,5291
described|5292,5301
above|5302,5307
.|5307,5308
<EOL>|5308,5309
.|5309,5310
<EOL>|5310,5311
HYPERTENSION|5311,5323
:|5323,5324
Pt|5325,5327
slightly|5328,5336
hypertensive|5337,5349
in|5350,5352
the|5353,5356
ED|5357,5359
,|5359,5360
but|5361,5364
will|5365,5369
<EOL>|5370,5371
continue|5371,5379
meds|5380,5384
at|5385,5387
current|5388,5395
regiment|5396,5404
and|5405,5408
reassess|5409,5417
in|5418,5420
the|5421,5424
morning|5425,5432
.|5432,5433
<EOL>|5435,5436
Her|5436,5439
BP|5440,5442
meds|5443,5447
are|5448,5451
actively|5452,5460
being|5461,5466
uptitrated|5467,5477
in|5478,5480
the|5481,5484
outpatient|5485,5495
<EOL>|5496,5497
setting|5497,5504
.|5504,5505
She|5507,5510
remained|5511,5519
normotensive|5520,5532
during|5533,5539
her|5540,5543
hospital|5544,5552
stay|5553,5557
on|5558,5560
<EOL>|5561,5562
the|5562,5565
floor|5566,5571
.|5571,5572
We|5574,5576
continued|5577,5586
Diltiazem|5587,5596
ER|5597,5599
360mg|5600,5605
PO|5606,5608
Q24H|5609,5613
,|5613,5614
HCTZ|5615,5619
12.5|5620,5624
mg|5624,5626
<EOL>|5627,5628
PO|5628,5630
DAILY|5631,5636
,|5636,5637
IMDUR|5638,5643
ER|5644,5646
60|5647,5649
mg|5650,5652
PO|5653,5655
DAILY|5656,5661
.|5661,5662
<EOL>|5662,5663
.|5663,5664
<EOL>|5666,5667
GERD|5667,5671
:|5671,5672
Currently|5673,5682
asymptomatic|5683,5695
.|5695,5696
We|5698,5700
continued|5701,5710
omeprazole|5711,5721
20mg|5722,5726
PO|5727,5729
<EOL>|5730,5731
Daily|5731,5736
<EOL>|5736,5737
.|5737,5738
<EOL>|5739,5740
CAD|5740,5743
:|5743,5744
Pt|5745,5747
was|5748,5751
recently|5752,5760
diagnosed|5761,5770
with|5771,5775
single|5776,5782
vessel|5783,5789
disease|5790,5797
.|5797,5798
She|5800,5803
<EOL>|5804,5805
is|5805,5807
asymptomatic|5808,5820
at|5821,5823
this|5824,5828
time|5829,5833
,|5833,5834
but|5835,5838
we|5839,5841
will|5842,5846
continue|5847,5855
to|5856,5858
monitor|5859,5866
<EOL>|5867,5868
her|5868,5871
for|5872,5875
symptoms|5876,5884
during|5885,5891
this|5892,5896
admission|5897,5906
.|5906,5907
<EOL>|5908,5909
We|5909,5911
continued|5912,5921
aspirin|5922,5929
81mg|5930,5934
PO|5935,5937
DAILY|5938,5943
<EOL>|5943,5944
.|5944,5945
<EOL>|5945,5946
TOBACCO|5946,5953
ABUSE|5954,5959
:|5959,5960
Pt|5961,5963
had|5964,5967
been|5968,5972
smoking|5973,5980
for|5981,5984
many|5985,5989
years|5990,5995
,|5995,5996
but|5997,6000
said|6001,6005
that|6006,6010
<EOL>|6011,6012
she|6012,6015
quit|6016,6020
yesterday|6021,6030
and|6031,6034
has|6035,6038
no|6039,6041
need|6042,6046
for|6047,6050
a|6051,6052
nicotine|6053,6061
patch|6062,6067
or|6068,6070
gum|6071,6074
<EOL>|6075,6076
at|6076,6078
this|6079,6083
time|6084,6088
.|6088,6089
<EOL>|6091,6092
.|6092,6093
<EOL>|6093,6094
<EOL>|6094,6095
<EOL>|6096,6097
Medications|6097,6108
on|6109,6111
Admission|6112,6121
:|6121,6122
<EOL>|6122,6123
1.|6123,6125
Lisinopril|6126,6136
5mg|6137,6140
PO|6141,6143
Daily|6144,6149
<EOL>|6149,6150
2|6150,6151
.|6151,6152
B|6153,6154
complex|6155,6162
-|6162,6163
vitamin|6163,6170
C|6171,6172
-|6172,6173
folic|6173,6178
acid|6179,6183
1|6184,6185
mg|6186,6188
Capsule|6189,6196
Sig|6197,6200
:|6200,6201
One|6202,6205
(|6206,6207
1|6207,6208
)|6208,6209
Cap|6210,6213
<EOL>|6215,6216
<EOL>|6216,6217
PO|6217,6219
DAILY|6220,6225
(|6226,6227
Daily|6227,6232
)|6232,6233
.|6233,6234
<EOL>|6236,6237
3.|6237,6239
cinacalcet|6240,6250
30|6251,6253
mg|6254,6256
Tablet|6257,6263
Sig|6264,6267
:|6267,6268
Two|6269,6272
(|6273,6274
2|6274,6275
)|6275,6276
Tablet|6277,6283
PO|6284,6286
DAILY|6287,6292
(|6293,6294
Daily|6294,6299
)|6299,6300
.|6300,6301
<EOL>|6302,6303
<EOL>|6304,6305
4.|6305,6307
simvastatin|6308,6319
10|6320,6322
mg|6323,6325
Tablet|6326,6332
Sig|6333,6336
:|6336,6337
Two|6338,6341
(|6342,6343
2|6343,6344
)|6344,6345
Tablet|6346,6352
PO|6353,6355
DAILY|6356,6361
<EOL>|6363,6364
(|6364,6365
Daily|6365,6370
)|6370,6371
.|6371,6372
<EOL>|6374,6375
5.|6375,6377
metoprolol|6378,6388
succinate|6389,6398
100|6399,6402
mg|6403,6405
Tablet|6406,6412
Sustained|6413,6422
Release|6423,6430
24|6431,6433
hr|6434,6436
<EOL>|6438,6439
Sig|6439,6442
:|6442,6443
One|6444,6447
(|6448,6449
1|6449,6450
)|6450,6451
Tablet|6452,6458
Sustained|6459,6468
Release|6469,6476
24|6477,6479
hr|6480,6482
PO|6483,6485
once|6486,6490
a|6491,6492
day|6493,6496
.|6496,6497
<EOL>|6499,6500
6.|6500,6502
doxazosin|6503,6512
4|6513,6514
mg|6515,6517
Tablet|6518,6524
Sig|6525,6528
:|6528,6529
Two|6530,6533
(|6534,6535
2|6535,6536
)|6536,6537
Tablet|6538,6544
PO|6545,6547
HS|6548,6550
(|6551,6552
at|6552,6554
bedtime|6555,6562
)|6562,6563
.|6563,6564
<EOL>|6565,6566
<EOL>|6567,6568
7.|6568,6570
aspirin|6571,6578
81|6579,6581
mg|6582,6584
Tablet|6585,6591
,|6591,6592
Chewable|6593,6601
Sig|6602,6605
:|6605,6606
One|6607,6610
(|6611,6612
1|6612,6613
)|6613,6614
Tablet|6615,6621
,|6621,6622
Chewable|6623,6631
<EOL>|6633,6634
<EOL>|6634,6635
PO|6635,6637
DAILY|6638,6643
(|6644,6645
Daily|6645,6650
)|6650,6651
.|6651,6652
<EOL>|6654,6655
8.|6655,6657
venlafaxine|6658,6669
75|6670,6672
mg|6673,6675
Capsule|6676,6683
,|6683,6684
Sust|6685,6689
.|6689,6690
Release|6691,6698
24|6699,6701
hr|6702,6704
Sig|6705,6708
:|6708,6709
Two|6710,6713
(|6714,6715
2|6715,6716
)|6716,6717
<EOL>|6719,6720
Capsule|6720,6727
,|6727,6728
Sust|6729,6733
.|6733,6734
Release|6735,6742
24|6743,6745
hr|6746,6748
PO|6749,6751
DAILY|6752,6757
(|6758,6759
Daily|6759,6764
)|6764,6765
.|6765,6766
<EOL>|6768,6769
9.|6769,6771
venlafaxine|6772,6783
37.5|6784,6788
mg|6789,6791
Capsule|6792,6799
,|6799,6800
Sust|6801,6805
.|6805,6806
Release|6807,6814
24|6815,6817
hr|6818,6820
Sig|6821,6824
:|6824,6825
One|6826,6829
(|6830,6831
1|6831,6832
)|6832,6833
<EOL>|6834,6835
<EOL>|6836,6837
Capsule|6837,6844
,|6844,6845
Sust|6846,6850
.|6850,6851
Release|6852,6859
24|6860,6862
hr|6863,6865
PO|6866,6868
DAILY|6869,6874
(|6875,6876
Daily|6876,6881
)|6881,6882
.|6882,6883
<EOL>|6885,6886
10.|6886,6889
sevelamer|6890,6899
HCl|6900,6903
400|6904,6907
mg|6908,6910
Tablet|6911,6917
Sig|6918,6921
:|6921,6922
Six|6923,6926
(|6927,6928
6|6928,6929
)|6929,6930
Tablet|6931,6937
PO|6938,6940
TID|6941,6944
<EOL>|6946,6947
W|6947,6948
/|6948,6949
MEALS|6949,6954
(|6955,6956
3|6956,6957
TIMES|6958,6963
A|6964,6965
DAY|6966,6969
WITH|6970,6974
MEALS|6975,6980
)|6980,6981
.|6981,6982
<EOL>|6984,6985
Disp|6985,6989
:|6989,6990
*|6990,6991
540|6991,6994
Tablet|6995,7001
(|7001,7002
s|7002,7003
)|7003,7004
*|7004,7005
Refills|7006,7013
:|7013,7014
*|7014,7015
2|7015,7016
*|7016,7017
<EOL>|7019,7020
11.|7020,7023
clonazepam|7024,7034
1|7035,7036
mg|7037,7039
Tablet|7040,7046
Sig|7047,7050
:|7050,7051
One|7052,7055
(|7056,7057
1|7057,7058
)|7058,7059
Tablet|7060,7066
PO|7067,7069
at|7070,7072
bedtime|7073,7080
.|7080,7081
<EOL>|7083,7084
<EOL>|7084,7085
<EOL>|7086,7087
Discharge|7087,7096
Medications|7097,7108
:|7108,7109
<EOL>|7109,7110
1.|7110,7112
acetaminophen|7113,7126
325|7127,7130
mg|7131,7133
Tablet|7134,7140
Sig|7141,7144
:|7144,7145
One|7146,7149
(|7150,7151
1|7151,7152
)|7152,7153
Tablet|7154,7160
PO|7161,7163
every|7164,7169
four|7170,7174
<EOL>|7175,7176
(|7176,7177
4|7177,7178
)|7178,7179
hours|7180,7185
as|7186,7188
needed|7189,7195
for|7196,7199
pain|7200,7204
.|7204,7205
<EOL>|7207,7208
2.|7208,7210
albuterol|7211,7220
sulfate|7221,7228
90|7229,7231
mcg|7232,7235
/|7235,7236
Actuation|7236,7245
HFA|7246,7249
Aerosol|7250,7257
Inhaler|7258,7265
Sig|7266,7269
:|7269,7270
<EOL>|7271,7272
Two|7272,7275
(|7276,7277
2|7277,7278
)|7278,7279
Inhalation|7281,7291
every|7292,7297
_|7298,7299
_|7299,7300
_|7300,7301
hours|7302,7307
.|7307,7308
<EOL>|7310,7311
3.|7311,7313
azithromycin|7314,7326
250|7327,7330
mg|7331,7333
Tablet|7334,7340
Sig|7341,7344
:|7344,7345
One|7346,7349
(|7350,7351
1|7351,7352
)|7352,7353
Tablet|7354,7360
PO|7361,7363
Q24H|7364,7368
(|7369,7370
every|7370,7375
<EOL>|7376,7377
24|7377,7379
hours|7380,7385
)|7385,7386
for|7387,7390
2|7391,7392
days|7393,7397
.|7397,7398
<EOL>|7398,7399
Disp|7399,7403
:|7403,7404
*|7404,7405
2|7405,7406
Tablet|7407,7413
(|7413,7414
s|7414,7415
)|7415,7416
*|7416,7417
Refills|7418,7425
:|7425,7426
*|7426,7427
0|7427,7428
*|7428,7429
<EOL>|7429,7430
4.|7430,7432
oseltamivir|7433,7444
75|7445,7447
mg|7448,7450
Capsule|7451,7458
Sig|7459,7462
:|7462,7463
One|7464,7467
(|7468,7469
1|7469,7470
)|7470,7471
Capsule|7472,7479
PO|7480,7482
BID|7483,7486
(|7487,7488
2|7488,7489
<EOL>|7490,7491
times|7491,7496
a|7497,7498
day|7499,7502
)|7502,7503
for|7504,7507
3|7508,7509
days|7510,7514
.|7514,7515
<EOL>|7515,7516
Disp|7516,7520
:|7520,7521
*|7521,7522
5|7522,7523
Capsule|7524,7531
(|7531,7532
s|7532,7533
)|7533,7534
*|7534,7535
Refills|7536,7543
:|7543,7544
*|7544,7545
0|7545,7546
*|7546,7547
<EOL>|7547,7548
5.|7548,7550
prednisone|7551,7561
10|7562,7564
mg|7565,7567
Tablet|7568,7574
Sig|7575,7578
:|7578,7579
Five|7580,7584
(|7585,7586
5|7586,7587
)|7587,7588
Tablet|7589,7595
PO|7596,7598
once|7599,7603
a|7604,7605
day|7606,7609
<EOL>|7610,7611
for|7611,7614
7|7615,7616
days|7617,7621
:|7621,7622
Take|7623,7627
5|7628,7629
tabs|7630,7634
for|7635,7638
2|7639,7640
days|7641,7645
,|7645,7646
then|7647,7651
4|7652,7653
tabs|7654,7658
for|7659,7662
2|7663,7664
days|7665,7669
,|7669,7670
then|7671,7675
<EOL>|7676,7677
2|7677,7678
tabs|7679,7683
for|7684,7687
2|7688,7689
days|7690,7694
,|7694,7695
then|7696,7700
1|7701,7702
tab|7703,7706
for|7707,7710
2|7711,7712
days|7713,7717
.|7717,7718
<EOL>|7718,7719
Disp|7719,7723
:|7723,7724
*|7724,7725
19|7725,7727
Tablet|7728,7734
(|7734,7735
s|7735,7736
)|7736,7737
*|7737,7738
Refills|7739,7746
:|7746,7747
*|7747,7748
0|7748,7749
*|7749,7750
<EOL>|7750,7751
6.|7751,7753
diltiazem|7754,7763
HCl|7764,7767
180|7768,7771
mg|7772,7774
Capsule|7775,7782
,|7782,7783
Extended|7784,7792
Release|7793,7800
Sig|7801,7804
:|7804,7805
Two|7806,7809
(|7810,7811
2|7811,7812
)|7812,7813
<EOL>|7814,7815
Capsule|7815,7822
,|7822,7823
Extended|7824,7832
Release|7833,7840
PO|7841,7843
DAILY|7844,7849
(|7850,7851
Daily|7851,7856
)|7856,7857
.|7857,7858
<EOL>|7860,7861
7.|7861,7863
fluticasone|7864,7875
50|7876,7878
mcg|7879,7882
/|7882,7883
Actuation|7883,7892
Spray|7893,7898
,|7898,7899
Suspension|7900,7910
Sig|7911,7914
:|7914,7915
One|7916,7919
(|7920,7921
1|7921,7922
)|7922,7923
<EOL>|7924,7925
Spray|7925,7930
Nasal|7931,7936
DAILY|7937,7942
(|7943,7944
Daily|7944,7949
)|7949,7950
.|7950,7951
<EOL>|7953,7954
8.|7954,7956
fluticasone|7957,7968
-|7968,7969
salmeterol|7969,7979
500|7980,7983
-|7983,7984
50|7984,7986
mcg|7987,7990
/|7990,7991
dose|7991,7995
Disk|7996,8000
with|8001,8005
Device|8006,8012
Sig|8013,8016
:|8016,8017
<EOL>|8018,8019
One|8019,8022
(|8023,8024
1|8024,8025
)|8025,8026
Disk|8027,8031
with|8032,8036
Device|8037,8043
Inhalation|8044,8054
BID|8055,8058
(|8059,8060
2|8060,8061
times|8062,8067
a|8068,8069
day|8070,8073
)|8073,8074
.|8074,8075
<EOL>|8077,8078
9.|8078,8080
hydrochlorothiazide|8081,8100
12.5|8101,8105
mg|8106,8108
Capsule|8109,8116
Sig|8117,8120
:|8120,8121
One|8122,8125
(|8126,8127
1|8127,8128
)|8128,8129
Capsule|8130,8137
PO|8138,8140
<EOL>|8141,8142
DAILY|8142,8147
(|8148,8149
Daily|8149,8154
)|8154,8155
.|8155,8156
<EOL>|8158,8159
10.|8159,8162
isosorbide|8163,8173
mononitrate|8174,8185
60|8186,8188
mg|8189,8191
Tablet|8192,8198
Extended|8199,8207
Release|8208,8215
24|8216,8218
hr|8219,8221
<EOL>|8222,8223
Sig|8223,8226
:|8226,8227
One|8228,8231
(|8232,8233
1|8233,8234
)|8234,8235
Tablet|8236,8242
Extended|8243,8251
Release|8252,8259
24|8260,8262
hr|8263,8265
PO|8266,8268
DAILY|8269,8274
(|8275,8276
Daily|8276,8281
)|8281,8282
.|8282,8283
<EOL>|8285,8286
11.|8286,8289
montelukast|8290,8301
10|8302,8304
mg|8305,8307
Tablet|8308,8314
Sig|8315,8318
:|8318,8319
One|8320,8323
(|8324,8325
1|8325,8326
)|8326,8327
Tablet|8328,8334
PO|8335,8337
DAILY|8338,8343
<EOL>|8344,8345
(|8345,8346
Daily|8346,8351
)|8351,8352
.|8352,8353
<EOL>|8355,8356
12.|8356,8359
omeprazole|8360,8370
20|8371,8373
mg|8374,8376
Capsule|8377,8384
,|8384,8385
Delayed|8386,8393
Release|8394,8401
(|8401,8402
E.C|8402,8405
.|8405,8406
)|8406,8407
Sig|8408,8411
:|8411,8412
One|8413,8416
(|8417,8418
1|8418,8419
)|8419,8420
<EOL>|8421,8422
Capsule|8422,8429
,|8429,8430
Delayed|8431,8438
Release|8439,8446
(|8446,8447
E.C|8447,8450
.|8450,8451
)|8451,8452
PO|8453,8455
DAILY|8456,8461
(|8462,8463
Daily|8463,8468
)|8468,8469
.|8469,8470
<EOL>|8472,8473
13.|8473,8476
tiotropium|8477,8487
bromide|8488,8495
18|8496,8498
mcg|8499,8502
Capsule|8503,8510
,|8510,8511
w|8512,8513
/|8513,8514
Inhalation|8514,8524
Device|8525,8531
Sig|8532,8535
:|8535,8536
<EOL>|8537,8538
One|8538,8541
(|8542,8543
1|8543,8544
)|8544,8545
Cap|8546,8549
Inhalation|8550,8560
DAILY|8561,8566
(|8567,8568
Daily|8568,8573
)|8573,8574
.|8574,8575
<EOL>|8577,8578
14.|8578,8581
calcium|8582,8589
carbonate|8590,8599
200|8600,8603
mg|8604,8606
(|8607,8608
500|8608,8611
mg|8612,8614
)|8614,8615
Tablet|8616,8622
,|8622,8623
Chewable|8624,8632
Sig|8633,8636
:|8636,8637
One|8638,8641
<EOL>|8642,8643
(|8643,8644
1|8644,8645
)|8645,8646
Tablet|8647,8653
,|8653,8654
Chewable|8655,8663
PO|8664,8666
DAILY|8667,8672
(|8673,8674
Daily|8674,8679
)|8679,8680
.|8680,8681
<EOL>|8683,8684
15.|8684,8687
multivitamin|8688,8700
Tablet|8705,8711
Sig|8712,8715
:|8715,8716
One|8717,8720
(|8721,8722
1|8722,8723
)|8723,8724
Tablet|8725,8731
PO|8732,8734
DAILY|8735,8740
<EOL>|8741,8742
(|8742,8743
Daily|8743,8748
)|8748,8749
.|8749,8750
<EOL>|8752,8753
16.|8753,8756
aspirin|8757,8764
81|8765,8767
mg|8768,8770
Tablet|8771,8777
Sig|8778,8781
:|8781,8782
One|8783,8786
(|8787,8788
1|8788,8789
)|8789,8790
Tablet|8791,8797
PO|8798,8800
once|8801,8805
a|8806,8807
day|8808,8811
.|8811,8812
<EOL>|8814,8815
17.|8815,8818
Oxygen|8819,8825
<EOL>|8825,8826
Home|8826,8830
Oxygen|8831,8837
@|8838,8839
2LPM|8840,8844
Continuous|8845,8855
via|8856,8859
nasal|8860,8865
cannula|8866,8873
,|8873,8874
conserving|8875,8885
<EOL>|8886,8887
device|8887,8893
for|8894,8897
portability|8898,8909
.|8909,8910
Pulse|8912,8917
dose|8918,8922
for|8923,8926
portability|8927,8938
.|8938,8939
<EOL>|8939,8940
<EOL>|8940,8941
<EOL>|8942,8943
Discharge|8943,8952
Disposition|8953,8964
:|8964,8965
<EOL>|8965,8966
Home|8966,8970
With|8971,8975
Service|8976,8983
<EOL>|8983,8984
<EOL>|8985,8986
Facility|8986,8994
:|8994,8995
<EOL>|8995,8996
_|8996,8997
_|8997,8998
_|8998,8999
<EOL>|8999,9000
<EOL>|9001,9002
Discharge|9002,9011
Diagnosis|9012,9021
:|9021,9022
<EOL>|9022,9023
Influenza|9042,9051
<EOL>|9051,9052
COPD|9052,9056
exacerbation|9057,9069
<EOL>|9069,9070
.|9070,9071
<EOL>|9071,9072
Secondary|9072,9081
Diagnosis|9082,9091
:|9091,9092
<EOL>|9092,9093
ASTHMA|9093,9099
<EOL>|9102,9103
HYPERTENSION|9103,9115
<EOL>|9118,9119
HYPERLIPIDEMIA|9119,9133
<EOL>|9136,9137
HEADACHE|9137,9145
<EOL>|9148,9149
OSTEOARTHRITIS|9149,9163
<EOL>|9166,9167
ATYPICAL|9167,9175
CHEST|9176,9181
PAIN|9182,9186
<EOL>|9189,9190
TOBACCO|9190,9197
ABUSE|9198,9203
<EOL>|9206,9207
ABNORMAL|9207,9215
CHEST|9216,9221
XRAY|9222,9226
<EOL>|9229,9230
COPD|9230,9234
<EOL>|9235,9236
<EOL>|9236,9237
<EOL>|9238,9239
Mental|9260,9266
Status|9267,9273
:|9273,9274
Clear|9275,9280
and|9281,9284
coherent|9285,9293
.|9293,9294
<EOL>|9294,9295
Level|9295,9300
of|9301,9303
Consciousness|9304,9317
:|9317,9318
Alert|9319,9324
and|9325,9328
interactive|9329,9340
.|9340,9341
<EOL>|9341,9342
Activity|9342,9350
Status|9351,9357
:|9357,9358
Ambulatory|9359,9369
-|9370,9371
Independent|9372,9383
.|9383,9384
<EOL>|9384,9385
<EOL>|9385,9386
<EOL>|9387,9388
You|9412,9415
are|9416,9419
being|9420,9425
discharged|9426,9436
from|9437,9441
_|9442,9443
_|9443,9444
_|9444,9445
.|9445,9446
It|9448,9450
<EOL>|9451,9452
was|9452,9455
a|9456,9457
pleasure|9458,9466
taking|9467,9473
care|9474,9478
of|9479,9481
you|9482,9485
.|9485,9486
You|9488,9491
were|9492,9496
admitted|9497,9505
to|9506,9508
the|9509,9512
<EOL>|9513,9514
hospital|9514,9522
for|9523,9526
symptoms|9527,9535
that|9536,9540
were|9541,9545
similar|9546,9553
to|9554,9556
a|9557,9558
common|9559,9565
cold|9566,9570
as|9571,9573
well|9574,9578
<EOL>|9579,9580
as|9580,9582
worsening|9583,9592
respiratory|9593,9604
status|9605,9611
.|9611,9612
You|9614,9617
tested|9618,9624
positive|9625,9633
for|9634,9637
the|9638,9641
<EOL>|9642,9643
flu|9643,9646
and|9647,9650
we|9651,9653
also|9654,9658
believe|9659,9666
that|9667,9671
you|9672,9675
are|9676,9679
having|9680,9686
a|9687,9688
COPD|9689,9693
exacerbation|9694,9706
.|9706,9707
<EOL>|9708,9709
You|9710,9713
were|9714,9718
started|9719,9726
on|9727,9729
high|9730,9734
dose|9735,9739
steroids|9740,9748
,|9748,9749
azithromycin|9750,9762
,|9762,9763
tamiflu|9764,9771
<EOL>|9772,9773
and|9773,9776
nebulizers|9777,9787
.|9787,9788
You|9790,9793
were|9794,9798
also|9799,9803
placed|9804,9810
on|9811,9813
oxygen|9814,9820
.|9820,9821
You|9823,9826
are|9827,9830
now|9831,9834
<EOL>|9835,9836
doing|9836,9841
better|9842,9848
,|9848,9849
but|9850,9853
may|9854,9857
require|9858,9865
O2|9866,9868
at|9869,9871
home|9872,9876
for|9877,9880
some|9881,9885
time|9886,9890
as|9891,9893
your|9894,9898
<EOL>|9899,9900
infection|9900,9909
resolves|9910,9918
and|9919,9922
your|9923,9927
inflammation|9928,9940
improves|9941,9949
.|9949,9950
<EOL>|9950,9951
.|9951,9952
<EOL>|9952,9953
The|9953,9956
Following|9957,9966
medications|9967,9978
were|9979,9983
STARTED|9984,9991
:|9991,9992
<EOL>|9992,9993
Prednisone|9993,10003
50mg|10004,10008
1|10009,10010
day|10011,10014
,|10014,10015
on|10016,10018
_|10019,10020
_|10020,10021
_|10021,10022
decrease|10023,10031
to|10032,10034
40mg|10035,10039
Daily|10040,10045
for|10046,10049
2|10050,10051
<EOL>|10052,10053
days|10053,10057
,|10057,10058
on|10059,10061
_|10062,10063
_|10063,10064
_|10064,10065
decrease|10066,10074
to|10075,10077
20mg|10078,10082
Daily|10083,10088
for|10089,10092
2|10093,10094
days|10095,10099
,|10099,10100
on|10101,10103
_|10104,10105
_|10105,10106
_|10106,10107
<EOL>|10108,10109
take|10109,10113
10mg|10114,10118
Daily|10119,10124
for|10125,10128
2|10129,10130
days|10131,10135
then|10136,10140
stop|10141,10145
<EOL>|10147,10148
Azithromycin|10148,10160
250mg|10161,10166
by|10167,10169
mouth|10170,10175
Daily|10176,10181
1|10182,10183
day|10184,10187
(|10188,10189
last|10189,10193
dose|10194,10198
on|10199,10201
_|10202,10203
_|10203,10204
_|10204,10205
<EOL>|10205,10206
Tamiflu|10206,10213
75mg|10214,10218
two|10219,10222
times|10223,10228
a|10229,10230
day|10231,10234
for|10235,10238
2.5|10239,10242
days|10243,10247
(|10248,10249
last|10249,10253
dose|10254,10258
on|10259,10261
_|10262,10263
_|10263,10264
_|10264,10265
<EOL>|10265,10266
You|10266,10269
will|10270,10274
also|10275,10279
be|10280,10282
sent|10283,10287
on|10288,10290
home|10291,10295
O2|10296,10298
<EOL>|10298,10299
.|10299,10300
<EOL>|10300,10301
Please|10301,10307
take|10308,10312
your|10313,10317
other|10318,10323
medications|10324,10335
as|10336,10338
prescribed|10339,10349
.|10349,10350
<EOL>|10350,10351
<EOL>|10352,10353
Followup|10353,10361
Instructions|10362,10374
:|10374,10375
<EOL>|10375,10376
_|10376,10377
_|10377,10378
_|10378,10379
<EOL>|10379,10380

