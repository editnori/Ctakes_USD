 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|46,55|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|46,55|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|46,60|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|80,89|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|80,89|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|80,94|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|136,139|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|147,154|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|147,154|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|156,164|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Drug|Organic Chemical|Allergies|179,186|false|false|false|C0009214|codeine|Codeine
Drug|Pharmacologic Substance|Allergies|179,186|false|false|false|C0009214|codeine|Codeine
Event|Event|Allergies|189,198|false|false|false|||Attending
Finding|Functional Concept|Allergies|189,198|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|Chief Complaint|224,229|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Finding|Sign or Symptom|Chief Complaint|224,229|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Finding|Classification|Chief Complaint|232,237|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|238,246|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|238,246|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|250,268|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|259,268|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|259,268|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|259,268|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|259,268|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|259,268|false|false|false|C0184661|Interventional procedure|Procedure
Attribute|Clinical Attribute|History of Present Illness|320,325|false|false|false|C1300072|Tumor stage|stage
Disorder|Neoplastic Process|History of Present Illness|320,348|false|false|false|C0854988|Adenocarcinoma of lung, stage IV|stage IV lung adenocarcinoma
Anatomy|Body Location or Region|History of Present Illness|329,333|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|329,333|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|History of Present Illness|329,333|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|History of Present Illness|329,333|false|false|false|C0740941|Lung Problem|lung
Disorder|Neoplastic Process|History of Present Illness|329,348|false|false|false|C0152013|Adenocarcinoma of lung (disorder)|lung adenocarcinoma
Disorder|Neoplastic Process|History of Present Illness|334,348|false|false|false|C0001418;C5551397|Adenocarcinoma;Malignant adenomatous neoplasm|adenocarcinoma
Event|Event|History of Present Illness|334,348|false|false|false|||adenocarcinoma
Drug|Organic Chemical|History of Present Illness|353,363|false|false|false|C0210657|pemetrexed|pemetrexed
Drug|Pharmacologic Substance|History of Present Illness|353,363|false|false|false|C0210657|pemetrexed|pemetrexed
Event|Event|History of Present Illness|353,363|false|false|false|||pemetrexed
Disorder|Disease or Syndrome|History of Present Illness|365,368|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|365,368|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|History of Present Illness|365,368|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|History of Present Illness|365,368|false|false|false|||CAD
Finding|Gene or Genome|History of Present Illness|365,368|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|History of Present Illness|365,368|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|History of Present Illness|365,368|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|365,368|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|History of Present Illness|370,373|false|false|false|C0001365;C0038454|Acute ill-defined cerebrovascular disease;Cerebrovascular accident|CVA
Drug|Pharmacologic Substance|History of Present Illness|370,373|false|false|false|C5779650|Cyclophosphamide/Doxorubicin/Vincristine|CVA
Event|Event|History of Present Illness|370,373|false|false|false|||CVA
Event|Event|History of Present Illness|374,383|false|false|false|||presented
Event|Event|History of Present Illness|389,394|false|false|false|||fever
Finding|Finding|History of Present Illness|389,394|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|History of Present Illness|389,394|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|History of Present Illness|400,404|false|false|false|||home
Finding|Idea or Concept|History of Present Illness|400,404|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|History of Present Illness|400,404|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|History of Present Illness|400,404|false|false|false|C1553498|home health encounter|home
Finding|Body Substance|History of Present Illness|406,413|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|406,413|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|406,413|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|History of Present Illness|419,424|false|false|false|||found
Event|Event|History of Present Illness|433,437|false|false|false|||temp
Finding|Gene or Genome|History of Present Illness|433,437|false|false|false|C1823816|C1orf210 gene|temp
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|433,437|false|false|false|C0279848|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|temp
Phenomenon|Natural Phenomenon or Process|History of Present Illness|486,490|false|false|false|C0678568||cool
Event|Event|History of Present Illness|491,501|false|false|false|||compresses
Drug|Organic Chemical|History of Present Illness|506,519|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Drug|Pharmacologic Substance|History of Present Illness|506,519|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Event|Event|History of Present Illness|506,519|false|false|false|||acetaminophen
Procedure|Laboratory Procedure|History of Present Illness|506,519|false|false|false|C0373527|Acetaminophen measurement|acetaminophen
Finding|Body Substance|History of Present Illness|521,528|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|521,528|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|521,528|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|History of Present Illness|529,536|false|false|false|||reports
Event|Event|History of Present Illness|576,582|false|false|false|||coughs
Finding|Finding|History of Present Illness|576,582|false|false|false|C0010200;C0687152|Coughing;Does cough|coughs
Finding|Sign or Symptom|History of Present Illness|576,582|false|false|false|C0010200;C0687152|Coughing;Does cough|coughs
Finding|Intellectual Product|History of Present Illness|584,588|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Sign or Symptom|History of Present Illness|589,593|false|false|false|C0234233;C1442877|Sore skin;Sore to touch|sore
Disorder|Disease or Syndrome|History of Present Illness|589,600|false|false|false|C0031350|Pharyngitis|sore throat
Drug|Organic Chemical|History of Present Illness|589,600|false|false|false|C0723402;C3244654|Sore Throat brand of Phenol;Sore Throat brand of benzocaine & menthol|sore throat
Drug|Pharmacologic Substance|History of Present Illness|589,600|false|false|false|C0723402;C3244654|Sore Throat brand of Phenol;Sore Throat brand of benzocaine & menthol|sore throat
Finding|Sign or Symptom|History of Present Illness|589,600|false|false|false|C0242429|Sore Throat|sore throat
Anatomy|Body Location or Region|History of Present Illness|594,600|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|594,600|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Drug|Pharmacologic Substance|History of Present Illness|594,600|false|false|false|C1950455|Throat Homeopathic Medication|throat
Event|Event|History of Present Illness|594,600|false|false|false|||throat
Finding|Body Substance|History of Present Illness|594,600|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Finding|Intellectual Product|History of Present Illness|594,600|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|607,612|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|History of Present Illness|607,612|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|History of Present Illness|607,612|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|History of Present Illness|607,612|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|History of Present Illness|607,612|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|History of Present Illness|607,612|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Sign or Symptom|History of Present Illness|607,623|false|false|false|C0027424|Nasal congestion (finding)|nasal congestion
Event|Event|History of Present Illness|613,623|false|false|false|||congestion
Finding|Pathologic Function|History of Present Illness|613,623|false|false|false|C0700148|Congestion|congestion
Event|Event|History of Present Illness|650,656|false|false|false|||states
Finding|Intellectual Product|History of Present Illness|680,701|false|false|false|C4526595|More Tired Than Usual|more tired than usual
Event|Event|History of Present Illness|685,690|false|false|false|||tired
Finding|Finding|History of Present Illness|685,690|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Finding|Intellectual Product|History of Present Illness|685,690|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Finding|Sign or Symptom|History of Present Illness|685,690|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Event|Event|History of Present Illness|696,701|false|false|false|||usual
Finding|Body Substance|History of Present Illness|703,710|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|703,710|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|703,710|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|History of Present Illness|715,723|false|false|false|||referred
Event|Event|History of Present Illness|751,753|false|false|false|||HR
Event|Event|History of Present Illness|783,787|false|false|false|||Exam
Finding|Functional Concept|History of Present Illness|783,787|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|History of Present Illness|783,787|false|false|false|C0582103|Medical Examination|Exam
Event|Event|History of Present Illness|789,801|false|false|false|||unremarkable
Event|Event|History of Present Illness|803,807|false|false|false|||Labs
Lab|Laboratory or Test Result|History of Present Illness|803,807|false|false|false|C0587081|Laboratory test finding|Labs
Event|Event|History of Present Illness|820,823|false|false|false|||ANC
Procedure|Laboratory Procedure|History of Present Illness|820,823|false|false|false|C0948762|Absolute neutrophil count|ANC
Drug|Biomedical or Dental Material|History of Present Illness|854,862|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|History of Present Illness|854,862|false|false|false|||baseline
Finding|Idea or Concept|History of Present Illness|854,862|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|History of Present Illness|873,876|false|false|false|||CXR
Procedure|Diagnostic Procedure|History of Present Illness|873,876|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|History of Present Illness|877,883|false|false|false|||showed
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|888,891|false|false|false|C1261077|Structure of left lower lobe of lung|LLL
Disorder|Disease or Syndrome|History of Present Illness|892,905|false|false|false|C0521530|Lung consolidation|consolidation
Event|Event|History of Present Illness|892,905|false|false|false|||consolidation
Finding|Finding|History of Present Illness|913,916|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|History of Present Illness|913,916|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|918,925|false|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|History of Present Illness|918,925|false|false|false|C1951340|Process Pharmacologic Substance|process
Event|Event|History of Present Illness|918,925|false|false|false|||process
Finding|Functional Concept|History of Present Illness|918,925|false|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|History of Present Illness|918,925|false|false|false|C1522240|Process|process
Event|Event|History of Present Illness|927,935|false|false|false|||Admitted
Event|Event|History of Present Illness|939,943|false|false|false|||OMED
Event|Event|History of Present Illness|956,966|false|false|false|||management
Event|Occupational Activity|History of Present Illness|956,966|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|History of Present Illness|956,966|false|false|false|C0376636|Disease Management|management
Attribute|Clinical Attribute|Patient History|1013,1018|false|false|false|C1300072|Tumor stage|Stage
Disorder|Neoplastic Process|Patient History|1013,1041|false|false|false|C0854988|Adenocarcinoma of lung, stage IV|Stage IV lung adenocarcinoma
Anatomy|Body Location or Region|Patient History|1022,1026|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Patient History|1022,1026|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Patient History|1022,1026|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Patient History|1022,1026|false|false|false|C0740941|Lung Problem|lung
Disorder|Neoplastic Process|Patient History|1022,1041|false|false|false|C0152013|Adenocarcinoma of lung (disorder)|lung adenocarcinoma
Disorder|Neoplastic Process|Patient History|1027,1041|false|false|false|C0001418;C5551397|Adenocarcinoma;Malignant adenomatous neoplasm|adenocarcinoma
Event|Event|Patient History|1027,1041|false|false|false|||adenocarcinoma
Event|Event|Patient History|1053,1062|false|false|false|||diagnosed
Attribute|Clinical Attribute|Patient History|1068,1073|false|false|false|C1300072|Tumor stage|stage
Anatomy|Body Location or Region|Patient History|1077,1081|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Patient History|1077,1081|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Patient History|1077,1081|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Patient History|1077,1081|false|false|false|C0740941|Lung Problem|lung
Event|Event|Patient History|1097,1106|false|false|false|||admission
Procedure|Health Care Activity|Patient History|1097,1106|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Disorder|Disease or Syndrome|Patient History|1111,1116|false|false|false|C1536220|ST segment elevation myocardial infarction|STEMI
Event|Event|Patient History|1111,1116|false|false|false|||STEMI
Finding|Finding|Patient History|1111,1116|false|false|false|C3538872|ST Elevation Myocardial Infarction by ECG Finding|STEMI
Event|Event|Patient History|1118,1126|false|false|false|||Received
Event|Event|Patient History|1137,1142|false|false|false|||cycle
Drug|Organic Chemical|Patient History|1146,1156|false|false|false|C0210657|pemetrexed|pemetrexed
Drug|Pharmacologic Substance|Patient History|1146,1156|false|false|false|C0210657|pemetrexed|pemetrexed
Event|Event|Patient History|1178,1183|false|false|false|||chemo
Procedure|Therapeutic or Preventive Procedure|Patient History|1178,1183|false|false|false|C0392920;C3665472|Chemotherapy;Chemotherapy Regimen|chemo
Drug|Organic Chemical|Patient History|1194,1204|false|false|false|C0210657|pemetrexed|pemetrexed
Drug|Pharmacologic Substance|Patient History|1194,1204|false|false|false|C0210657|pemetrexed|pemetrexed
Event|Event|Patient History|1227,1234|false|false|false|||treated
Event|Event|Patient History|1244,1250|false|false|false|||course
Finding|Idea or Concept|Patient History|1263,1267|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|Patient History|1263,1267|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|Patient History|1283,1290|false|false|false|||courses
Drug|Antibiotic|Patient History|1294,1305|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|Patient History|1294,1305|false|false|false|||antibiotics
Anatomy|Body Part, Organ, or Organ Component|Patient History|1310,1313|false|false|false|C1261075|Structure of right lower lobe of lung|RLL
Finding|Finding|Patient History|1310,1313|false|false|false|C5703311|Radiolucent Lines|RLL
Disorder|Disease or Syndrome|Patient History|1314,1323|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|Patient History|1314,1323|false|false|false|||pneumonia
Event|Event|Patient History|1331,1337|false|false|false|||failed
Event|Event|Patient History|1342,1349|false|false|false|||resolve
Finding|Conceptual Entity|Patient History|1342,1349|false|false|false|C2699488|Resolution|resolve
Procedure|Diagnostic Procedure|Patient History|1342,1349|false|false|false|C5401470|RESOLVE Multishot Diffusion Weighted Echoplanar Imaging|resolve
Finding|Intellectual Product|Patient History|1353,1359|false|false|false|C0031082|Periodicals|serial
Anatomy|Body Location or Region|Patient History|1360,1365|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Patient History|1360,1365|false|false|false|C0741025|Chest problem|chest
Procedure|Diagnostic Procedure|Patient History|1360,1373|false|false|false|C1531652|Chest imaging|chest imaging
Event|Event|Patient History|1366,1373|false|false|false|||imaging
Finding|Finding|Patient History|1366,1373|false|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|Patient History|1366,1373|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Disorder|Disease or Syndrome|Patient History|1402,1414|false|false|false|C0242339|Dyslipidemias|Dyslipidemia
Event|Event|Patient History|1402,1414|false|false|false|||Dyslipidemia
Disorder|Disease or Syndrome|Patient History|1417,1429|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|Patient History|1417,1429|false|false|false|||Hypertension
Disorder|Disease or Syndrome|Patient History|1434,1437|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Patient History|1434,1437|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Patient History|1434,1437|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Patient History|1434,1437|false|false|false|||CAD
Finding|Gene or Genome|Patient History|1434,1437|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Patient History|1434,1437|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Patient History|1434,1437|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Patient History|1434,1437|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Anatomy|Body Location or Region|Patient History|1466,1472|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|Patient History|1466,1472|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Event|Event|Patient History|1473,1477|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|Patient History|1473,1477|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Anatomy|Body Part, Organ, or Organ Component|Patient History|1484,1487|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|Patient History|1484,1487|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|Patient History|1484,1487|false|false|false|||LAD
Finding|Gene or Genome|Patient History|1484,1487|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Disorder|Disease or Syndrome|Patient History|1494,1497|false|false|false|C0006430|Burning Mouth Syndrome|BMS
Event|Event|Patient History|1494,1497|false|false|false|||BMS
Anatomy|Body Part, Organ, or Organ Component|Patient History|1501,1504|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|Patient History|1501,1504|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|Patient History|1501,1504|false|false|false|||LAD
Finding|Gene or Genome|Patient History|1501,1504|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Disorder|Disease or Syndrome|Patient History|1518,1526|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Disorder|Disease or Syndrome|Patient History|1527,1532|false|false|false|C1536220|ST segment elevation myocardial infarction|STEMI
Event|Event|Patient History|1527,1532|false|false|false|||STEMI
Finding|Finding|Patient History|1527,1532|false|false|false|C3538872|ST Elevation Myocardial Infarction by ECG Finding|STEMI
Disorder|Disease or Syndrome|Patient History|1535,1538|false|false|false|C0001365;C0038454|Acute ill-defined cerebrovascular disease;Cerebrovascular accident|CVA
Drug|Pharmacologic Substance|Patient History|1535,1538|false|false|false|C5779650|Cyclophosphamide/Doxorubicin/Vincristine|CVA
Event|Event|Patient History|1535,1538|false|false|false|||CVA
Finding|Functional Concept|Patient History|1547,1551|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Disorder|Disease or Syndrome|Patient History|1552,1561|false|false|false|C0751438|Posterior pituitary disease|posterior
Event|Event|Patient History|1570,1577|false|false|false|||infarct
Finding|Pathologic Function|Patient History|1570,1577|false|false|false|C0021308|Infarction|infarct
Event|Event|Patient History|1591,1594|false|false|false|||PFO
Event|Event|Patient History|1605,1617|false|false|false|||Degereration
Finding|Conceptual Entity|Family Medical History|1660,1666|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Finding|Idea or Concept|Family Medical History|1660,1666|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Event|Event|Family Medical History|1667,1671|false|false|false|||died
Disorder|Disease or Syndrome|Family Medical History|1679,1682|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Family Medical History|1679,1682|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Family Medical History|1679,1682|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Family Medical History|1679,1682|false|false|false|||CAD
Finding|Gene or Genome|Family Medical History|1679,1682|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Family Medical History|1679,1682|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Family Medical History|1679,1682|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Family Medical History|1679,1682|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Attribute|Clinical Attribute|Family Medical History|1686,1689|false|false|false|C1114365||age
Drug|Biologically Active Substance|Family Medical History|1686,1689|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|Family Medical History|1686,1689|false|false|false|C0162574|Glycation End Products, Advanced|age
Event|Event|Family Medical History|1686,1689|false|false|false|||age
Finding|Idea or Concept|Family Medical History|1699,1705|false|false|false|C1546508|Relationship - Mother|mother
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1710,1717|false|false|false|C0038351;C3714551;C4266636|Abdomen>Stomach;Stomach;Stomach structure|stomach
Disorder|Disease or Syndrome|Family Medical History|1710,1717|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Disorder|Neoplastic Process|Family Medical History|1710,1717|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Event|Event|Family Medical History|1710,1717|false|false|false|||stomach
Finding|Finding|Family Medical History|1710,1717|false|false|false|C0577027|Stomach problem|stomach
Procedure|Therapeutic or Preventive Procedure|Family Medical History|1710,1717|false|false|false|C0872393|Procedure on stomach|stomach
Disorder|Neoplastic Process|Family Medical History|1719,1725|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Family Medical History|1719,1725|false|false|false|||cancer
Disorder|Neoplastic Process|Family Medical History|1730,1742|false|false|false|C0029463;C0585442|Osteosarcoma;Osteosarcoma of bone|osteosarcoma
Event|Event|Family Medical History|1730,1742|false|false|false|||osteosarcoma
Finding|Gene or Genome|Family Medical History|1730,1742|false|false|false|C0694889|RB1 gene|osteosarcoma
Event|Event|Family Medical History|1747,1754|false|false|false|||history
Finding|Conceptual Entity|Family Medical History|1747,1754|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|1747,1754|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Family Medical History|1747,1754|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|1747,1757|false|false|false|C0262926|Medical History|history of
Anatomy|Body Location or Region|Family Medical History|1758,1762|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1758,1762|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Family Medical History|1758,1762|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Family Medical History|1758,1762|false|false|false|C0740941|Lung Problem|lung
Disorder|Neoplastic Process|Family Medical History|1758,1769|true|false|false|C0242379;C0684249|Carcinoma of lung;Malignant neoplasm of lung|lung cancer
Disorder|Neoplastic Process|Family Medical History|1763,1769|true|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Family Medical History|1763,1769|false|false|false|||cancer
Disorder|Neoplastic Process|Family Medical History|1763,1776|true|false|false|C0007102|Malignant tumor of colon|cancer, colon
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1771,1776|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|Family Medical History|1771,1776|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|Family Medical History|1771,1776|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Finding|Finding|Family Medical History|1771,1776|false|false|false|C0750873|COLON PROBLEM|colon
Disorder|Neoplastic Process|Family Medical History|1771,1783|true|false|false|C0007102;C0346629;C0699790|Colon Carcinoma;Malignant neoplasm of large intestine;Malignant tumor of colon|colon cancer
Disorder|Neoplastic Process|Family Medical History|1777,1783|true|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Family Medical History|1777,1783|false|false|false|||cancer
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1788,1794|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|Family Medical History|1788,1794|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Event|Event|Family Medical History|1788,1794|false|false|false|||breast
Finding|Finding|Family Medical History|1788,1794|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|Family Medical History|1788,1794|false|false|false|C0191838|Procedures on breast|breast
Disorder|Neoplastic Process|Family Medical History|1788,1801|false|false|false|C0006142;C0678222|Breast Carcinoma;Malignant neoplasm of breast|breast cancer
Disorder|Neoplastic Process|Family Medical History|1795,1801|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Family Medical History|1795,1801|false|false|false|||cancer
Finding|Classification|General Exam|1820,1823|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Finding|Gene or Genome|General Exam|1820,1823|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Event|Event|General Exam|1833,1838|false|false|false|||woman
Disorder|Disease or Syndrome|General Exam|1842,1845|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|1842,1845|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|1842,1845|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|1842,1845|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|1842,1845|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|General Exam|1842,1845|false|false|false|||NAD
Finding|Finding|General Exam|1842,1845|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|General Exam|1846,1851|false|false|false|C1512338|HEENT|HEENT
Event|Event|General Exam|1853,1857|false|false|false|||EOMI
Event|Event|General Exam|1876,1882|false|false|false|||lesion
Finding|Finding|General Exam|1876,1882|true|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|General Exam|1876,1882|true|false|false|C0221198;C1546698|Lesion|lesion
Anatomy|Body Location or Region|General Exam|1883,1887|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|General Exam|1883,1887|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|General Exam|1883,1887|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|General Exam|1889,1895|false|false|false|||supple
Finding|Functional Concept|General Exam|1889,1895|false|false|false|C0332254|Supple|supple
Anatomy|Body Part, Organ, or Organ Component|General Exam|1900,1903|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|General Exam|1900,1903|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|General Exam|1900,1903|false|false|false|||LAD
Finding|Gene or Genome|General Exam|1900,1903|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Event|General Exam|1908,1911|false|false|false|||RRR
Anatomy|Body Part, Organ, or Organ Component|General Exam|1936,1941|false|false|false|C0024109|Lung|Lungs
Finding|Intellectual Product|General Exam|1943,1947|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|Poor
Event|Event|General Exam|1948,1956|false|false|false|||aeration
Procedure|Therapeutic or Preventive Procedure|General Exam|1948,1956|false|false|false|C2215609|aeration|aeration
Anatomy|Body Location or Region|General Exam|1962,1966|false|false|false|C2987514|Anatomical base|base
Drug|Biomedical or Dental Material|General Exam|1962,1966|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Chemical Viewed Functionally|General Exam|1962,1966|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|1962,1966|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Finding|Gene or Genome|General Exam|1962,1966|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Finding|Idea or Concept|General Exam|1962,1966|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Anatomy|Body Location or Region|General Exam|1967,1970|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|Abd
Disorder|Cell or Molecular Dysfunction|General Exam|1967,1970|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|Abd
Disorder|Disease or Syndrome|General Exam|1972,1976|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|General Exam|1972,1976|false|false|false|||soft
Event|Event|General Exam|1989,1996|false|false|false|||present
Finding|Finding|General Exam|1989,1996|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|General Exam|1989,1996|false|false|false|C0150312;C0449450|Present;Presentation|present
Disorder|Congenital Abnormality|General Exam|1997,2000|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|General Exam|1997,2000|false|false|false|||Ext
Finding|Gene or Genome|General Exam|1997,2000|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Anatomy|Cell|General Exam|2032,2035|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|2042,2045|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|2042,2045|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|2042,2045|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|2052,2055|false|false|false|C0019046|Hemoglobin|HGB
Drug|Biologically Active Substance|General Exam|2052,2055|false|false|false|C0019046|Hemoglobin|HGB
Event|Event|General Exam|2052,2055|false|false|false|||HGB
Finding|Gene or Genome|General Exam|2052,2055|false|false|false|C1424337|CYGB gene|HGB
Lab|Laboratory or Test Result|General Exam|2052,2055|false|false|false|C0019029|Hemoglobin concentration|HGB
Procedure|Laboratory Procedure|General Exam|2061,2064|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|General Exam|2061,2064|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Disorder|Virus|General Exam|2071,2074|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|2071,2074|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|2071,2074|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|2071,2074|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|2071,2074|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Event|Event|General Exam|2095,2101|false|false|false|||LYMPHS
Finding|Body Substance|General Exam|2095,2101|false|false|false|C0024202|Lymph|LYMPHS
Drug|Antibiotic|General Exam|2106,2111|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Biomedical or Dental Material|General Exam|2106,2111|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Organic Chemical|General Exam|2106,2111|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Disorder|Disease or Syndrome|General Exam|2116,2119|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|EOS
Event|Event|General Exam|2116,2119|false|false|false|||EOS
Finding|Gene or Genome|General Exam|2116,2119|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|EOS
Event|Event|General Exam|2153,2156|false|false|false|||PLT
Procedure|Laboratory Procedure|General Exam|2153,2156|false|false|false|C0201617|Primed lymphocyte test|PLT
Drug|Biologically Active Substance|General Exam|2169,2176|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|General Exam|2169,2176|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|General Exam|2169,2176|false|false|false|C0017725|glucose|GLUCOSE
Event|Event|General Exam|2169,2176|false|false|false|||GLUCOSE
Lab|Laboratory or Test Result|General Exam|2169,2176|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|General Exam|2169,2176|false|false|false|C0337438|Glucose measurement|GLUCOSE
Drug|Biologically Active Substance|General Exam|2182,2186|false|false|false|C0041942|urea|UREA
Drug|Organic Chemical|General Exam|2182,2186|false|false|false|C0041942|urea|UREA
Drug|Pharmacologic Substance|General Exam|2182,2186|false|false|false|C0041942|urea|UREA
Event|Event|General Exam|2182,2186|false|false|false|||UREA
Procedure|Laboratory Procedure|General Exam|2182,2186|false|false|false|C0523961|Urea measurement|UREA
Drug|Biologically Active Substance|General Exam|2204,2210|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Element, Ion, or Isotope|General Exam|2204,2210|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Pharmacologic Substance|General Exam|2204,2210|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Event|Event|General Exam|2204,2210|false|false|false|||SODIUM
Finding|Physiologic Function|General Exam|2204,2210|false|false|false|C4553025|Sodium metabolic function|SODIUM
Procedure|Laboratory Procedure|General Exam|2204,2210|false|false|false|C0337443|Sodium measurement|SODIUM
Drug|Biologically Active Substance|General Exam|2216,2225|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Element, Ion, or Isotope|General Exam|2216,2225|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Food|General Exam|2216,2225|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Inorganic Chemical|General Exam|2216,2225|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Pharmacologic Substance|General Exam|2216,2225|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Finding|Physiologic Function|General Exam|2216,2225|false|false|false|C4553027|Potassium metabolic function|POTASSIUM
Procedure|Laboratory Procedure|General Exam|2216,2225|false|false|false|C0202194|Potassium measurement|POTASSIUM
Drug|Element, Ion, or Isotope|General Exam|2231,2239|false|false|false|C0008203;C0596019|Chlorides;chloride ion|CHLORIDE
Event|Event|General Exam|2231,2239|false|false|false|||CHLORIDE
Finding|Physiologic Function|General Exam|2231,2239|false|false|false|C4553021|Chloride metabolic function|CHLORIDE
Procedure|Laboratory Procedure|General Exam|2231,2239|false|false|false|C0201952|Chloride measurement|CHLORIDE
Drug|Biologically Active Substance|General Exam|2249,2252|false|false|false|C0007012|carbon dioxide|CO2
Drug|Inorganic Chemical|General Exam|2249,2252|false|false|false|C0007012|carbon dioxide|CO2
Event|Event|General Exam|2249,2252|false|false|false|||CO2
Finding|Finding|General Exam|2249,2252|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Finding|Gene or Genome|General Exam|2249,2252|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Drug|Organic Chemical|General Exam|2256,2263|false|false|false|C0022924;C0376261|Lactates;lactate|LACTATE
Drug|Pharmacologic Substance|General Exam|2256,2263|false|false|false|C0022924;C0376261|Lactates;lactate|LACTATE
Event|Event|General Exam|2256,2263|false|false|false|||LACTATE
Procedure|Laboratory Procedure|General Exam|2256,2263|false|false|false|C0202115|Lactic acid measurement|LACTATE
Finding|Body Substance|General Exam|2269,2274|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|2269,2274|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|2269,2274|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Finding|General Exam|2269,2281|false|false|false|C0278030|Color of urine|URINE  COLOR
Drug|Biomedical or Dental Material|General Exam|2276,2281|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|COLOR
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|2276,2281|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|COLOR
Event|Event|General Exam|2276,2281|false|false|false|||COLOR
Finding|Idea or Concept|General Exam|2296,2301|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Body Substance|General Exam|2309,2314|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|2309,2314|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|2309,2314|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Disorder|Disease or Syndrome|General Exam|2309,2321|false|false|false|C0018965|Hematuria|URINE  BLOOD
Disorder|Disease or Syndrome|General Exam|2316,2321|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2316,2321|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2316,2321|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Biologically Active Substance|General Exam|2325,2332|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Drug|Inorganic Chemical|General Exam|2325,2332|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Drug|Pharmacologic Substance|General Exam|2325,2332|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Finding|Finding|General Exam|2333,2336|false|false|false|C5848551|Neg - answer|NEG
Drug|Amino Acid, Peptide, or Protein|General Exam|2337,2344|false|false|false|C0033684|Proteins|PROTEIN
Drug|Biologically Active Substance|General Exam|2337,2344|false|false|false|C0033684|Proteins|PROTEIN
Event|Event|General Exam|2337,2344|false|false|false|||PROTEIN
Finding|Conceptual Entity|General Exam|2337,2344|false|false|false|C1521746|Protein Info|PROTEIN
Procedure|Laboratory Procedure|General Exam|2337,2344|false|false|false|C0202202|Protein measurement|PROTEIN
Drug|Biologically Active Substance|General Exam|2348,2355|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|General Exam|2348,2355|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|General Exam|2348,2355|false|false|false|C0017725|glucose|GLUCOSE
Event|Event|General Exam|2348,2355|false|false|false|||GLUCOSE
Lab|Laboratory or Test Result|General Exam|2348,2355|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|General Exam|2348,2355|false|false|false|C0337438|Glucose measurement|GLUCOSE
Event|Event|General Exam|2356,2359|false|false|false|||NEG
Finding|Finding|General Exam|2356,2359|false|false|false|C5848551|Neg - answer|NEG
Drug|Organic Chemical|General Exam|2360,2366|false|false|false|C0022634|Ketones|KETONE
Event|Event|General Exam|2360,2366|false|false|false|||KETONE
Event|Event|General Exam|2367,2370|false|false|false|||NEG
Finding|Finding|General Exam|2367,2370|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|General Exam|2372,2381|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Drug|Organic Chemical|General Exam|2372,2381|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Drug|Pharmacologic Substance|General Exam|2372,2381|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Procedure|Laboratory Procedure|General Exam|2372,2381|false|false|false|C0201913;C0863174|Bilirubin, total measurement;blood bilirubin level test|BILIRUBIN
Event|Event|General Exam|2382,2385|false|false|false|||NEG
Finding|Finding|General Exam|2382,2385|false|false|false|C5848551|Neg - answer|NEG
Event|Event|General Exam|2396,2399|false|false|false|||NEG
Finding|Finding|General Exam|2396,2399|false|false|false|C5848551|Neg - answer|NEG
Event|Event|General Exam|2412,2415|false|false|false|||NEG
Finding|Finding|General Exam|2412,2415|false|false|false|C5848551|Neg - answer|NEG
Finding|Body Substance|General Exam|2416,2421|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|2416,2421|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|2416,2421|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|2427,2435|false|false|false|C1510439|bacteria aspects|BACTERIA
Drug|Food|General Exam|2440,2445|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Immunologic Factor|General Exam|2440,2445|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|2440,2445|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Pharmacologic Substance|General Exam|2440,2445|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Event|Event|General Exam|2440,2445|false|false|false|||YEAST
Event|Event|General Exam|2446,2450|false|false|false|||NONE
Event|Event|General Exam|2455,2460|false|false|false|||TRANS
Finding|Finding|General Exam|2455,2460|false|false|false|C0558141|Transsexual (finding)|TRANS
Event|Event|General Exam|2467,2474|false|false|false|||STUDIES
Procedure|Research Activity|General Exam|2467,2474|false|false|false|C0947630|Scientific Study|STUDIES
Anatomy|Body Location or Region|General Exam|2477,2482|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|General Exam|2477,2482|false|false|false|C0741025|Chest problem|Chest
Procedure|Diagnostic Procedure|General Exam|2477,2487|false|false|false|C0039985|Plain chest X-ray|Chest Xray
Phenomenon|Natural Phenomenon or Process|General Exam|2483,2487|false|false|false|C0043309|Roentgen Rays|Xray
Procedure|Diagnostic Procedure|General Exam|2483,2487|false|false|false|C0043299|Diagnostic radiologic examination|Xray
Finding|Mental Process|General Exam|2500,2507|false|false|false|C0542559|contextual factors|setting
Disorder|Neoplastic Process|General Exam|2521,2546|false|false|false|C0007120|Bronchioloalveolar Adenocarcinoma|bronchoalveolar carcinoma
Disorder|Neoplastic Process|General Exam|2537,2546|false|false|false|C0007097|Carcinoma|carcinoma
Event|Event|General Exam|2537,2546|false|false|false|||carcinoma
Disorder|Anatomical Abnormality|General Exam|2557,2564|false|false|false|C1689985|Absence (morphologic abnormality)|absence
Event|Event|General Exam|2557,2564|false|false|false|||absence
Finding|Functional Concept|General Exam|2557,2564|false|false|false|C0332197|Absent|absence
Finding|Functional Concept|General Exam|2557,2567|false|false|false|C0332197|Absent|absence of
Event|Event|General Exam|2587,2594|false|false|false|||studies
Procedure|Research Activity|General Exam|2587,2594|false|false|false|C0947630|Scientific Study|studies
Finding|Finding|General Exam|2596,2599|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|General Exam|2596,2599|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Disorder|Disease or Syndrome|General Exam|2600,2609|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|General Exam|2600,2609|false|false|false|||pneumonia
Event|Event|General Exam|2619,2628|false|false|false|||difficult
Finding|Finding|General Exam|2619,2628|false|false|false|C0332218|Difficult (qualifier value)|difficult
Event|Event|General Exam|2633,2642|false|false|false|||recognize
Finding|Functional Concept|General Exam|2650,2655|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|General Exam|2656,2661|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|2656,2661|false|false|false|C2003888|Lower (action)|lower
Finding|Intellectual Product|General Exam|2666,2672|false|false|false|C1552826|Table Cell Vertical Align - middle|middle
Anatomy|Body Part, Organ, or Organ Component|General Exam|2673,2678|false|false|false|C0796494|lobe|lobes
Attribute|Clinical Attribute|General Exam|2682,2690|false|false|false|C0881858||CT Chest
Procedure|Diagnostic Procedure|General Exam|2682,2690|false|false|false|C0202823|Chest CT|CT Chest
Anatomy|Body Location or Region|General Exam|2685,2690|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|General Exam|2685,2690|false|false|false|C0741025|Chest problem|Chest
Event|Event|General Exam|2700,2709|false|false|false|||Increased
Anatomy|Body Part, Organ, or Organ Component|General Exam|2710,2719|false|false|false|C0205039;C1442216|Bronchial;Bronchial system|bronchial
Drug|Organic Chemical|General Exam|2710,2719|false|false|false|C0719022|Bronchial brand of guaifenesin-theophylline|bronchial
Drug|Pharmacologic Substance|General Exam|2710,2719|false|false|false|C0719022|Bronchial brand of guaifenesin-theophylline|bronchial
Event|Event|General Exam|2710,2719|false|false|false|||bronchial
Finding|Body Substance|General Exam|2710,2719|false|false|false|C1546565;C1550618|Bronchial Specimen;Bronchial Specimen Source Codes|bronchial
Finding|Intellectual Product|General Exam|2710,2719|false|false|false|C1546565;C1550618|Bronchial Specimen;Bronchial Specimen Source Codes|bronchial
Event|Event|General Exam|2738,2745|false|false|false|||nodules
Disorder|Disease or Syndrome|General Exam|2759,2764|false|false|false|C2676739|Chromosome 2q32-Q33 Deletion Syndrome|glass
Drug|Hazardous or Poisonous Substance|General Exam|2759,2764|false|false|false|C0025611|methamphetamine|glass
Drug|Organic Chemical|General Exam|2759,2764|false|false|false|C0025611|methamphetamine|glass
Drug|Pharmacologic Substance|General Exam|2759,2764|false|false|false|C0025611|methamphetamine|glass
Event|Event|General Exam|2759,2764|false|false|false|||glass
Event|Event|General Exam|2783,2796|false|false|false|||predominating
Finding|Intellectual Product|General Exam|2807,2813|false|false|false|C1552826|Table Cell Vertical Align - middle|middle
Anatomy|Body Part, Organ, or Organ Component|General Exam|2814,2819|false|false|false|C0796494|lobe|lobes
Event|Event|General Exam|2827,2837|false|false|false|||consistent
Finding|Idea or Concept|General Exam|2827,2837|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|General Exam|2827,2842|false|false|false|C0332290|Consistent with|consistent with
Disorder|Disease or Syndrome|General Exam|2843,2852|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|General Exam|2843,2852|false|false|false|||infection
Finding|Pathologic Function|General Exam|2843,2852|false|false|false|C3714514|Infection|infection
Finding|Intellectual Product|General Exam|2858,2864|false|false|false|C1547311|Patient Condition Code - Stable|Stable
Finding|Functional Concept|General Exam|2865,2870|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|General Exam|2865,2881|false|false|false|C1261075|Structure of right lower lobe of lung|right lower lobe
Anatomy|Body Location or Region|General Exam|2871,2876|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|2871,2876|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|General Exam|2871,2881|false|false|false|C0225758|Structure of lower lobe of lung|lower lobe
Anatomy|Body Part, Organ, or Organ Component|General Exam|2877,2881|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|General Exam|2877,2881|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Event|Event|General Exam|2892,2901|false|false|false|||opacities
Finding|Finding|General Exam|2892,2901|false|true|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacities
Finding|Pathologic Function|General Exam|2892,2901|false|true|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacities
Event|Event|General Exam|2907,2912|false|false|false|||areas
Disorder|Disease or Syndrome|General Exam|2917,2930|false|false|false|C0521530|Lung consolidation|consolidation
Event|Event|General Exam|2917,2930|false|false|false|||consolidation
Event|Event|General Exam|2947,2954|false|false|false|||nodules
Event|Event|General Exam|2969,2978|false|false|false|||involving
Finding|Functional Concept|General Exam|2983,2988|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Finding|Intellectual Product|General Exam|3000,3006|false|false|false|C1552826|Table Cell Vertical Align - middle|middle
Anatomy|Body Part, Organ, or Organ Component|General Exam|3008,3013|false|false|false|C0796494|lobe|lobes
Event|Event|General Exam|3015,3025|false|false|false|||consistent
Finding|Idea or Concept|General Exam|3015,3025|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|General Exam|3015,3030|false|false|false|C0332290|Consistent with|consistent with
Anatomy|Cell|General Exam|3054,3058|false|false|false|C0007634|Cells|cell
Finding|Gene or Genome|General Exam|3054,3058|false|false|false|C1413336;C1413337|CEL gene;CELP gene|cell
Disorder|Neoplastic Process|General Exam|3059,3068|false|false|false|C0007097|Carcinoma|carcinoma
Event|Event|General Exam|3059,3068|false|false|false|||carcinoma
Finding|Intellectual Product|General Exam|3074,3080|false|false|false|C1547311|Patient Condition Code - Stable|Stable
Finding|Gene or Genome|General Exam|3081,3086|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Finding|Functional Concept|General Exam|3087,3091|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|General Exam|3092,3099|false|false|false|C0040132|Thyroid Gland|thyroid
Disorder|Disease or Syndrome|General Exam|3092,3099|false|false|false|C0040128|Thyroid Diseases|thyroid
Drug|Amino Acid, Peptide, or Protein|General Exam|3092,3099|false|false|false|C0040134;C3540038;C5781115|THYROID;THYROID DIAGNOSTIC RADIOPHARMACEUTICALS;thyroid (USP)|thyroid
Drug|Hormone|General Exam|3092,3099|false|false|false|C0040134;C3540038;C5781115|THYROID;THYROID DIAGNOSTIC RADIOPHARMACEUTICALS;thyroid (USP)|thyroid
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|3092,3099|false|false|false|C0040134;C3540038;C5781115|THYROID;THYROID DIAGNOSTIC RADIOPHARMACEUTICALS;thyroid (USP)|thyroid
Drug|Organic Chemical|General Exam|3092,3099|false|false|false|C0040134;C3540038;C5781115|THYROID;THYROID DIAGNOSTIC RADIOPHARMACEUTICALS;thyroid (USP)|thyroid
Drug|Pharmacologic Substance|General Exam|3092,3099|false|false|false|C0040134;C3540038;C5781115|THYROID;THYROID DIAGNOSTIC RADIOPHARMACEUTICALS;thyroid (USP)|thyroid
Procedure|Health Care Activity|General Exam|3092,3099|false|false|false|C2228489|examination of thyroid|thyroid
Finding|Finding|General Exam|3092,3104|false|false|false|C0349453|Mass of thyroid gland|thyroid mass
Event|Event|General Exam|3100,3104|false|false|false|||mass
Finding|Finding|General Exam|3100,3104|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|General Exam|3100,3104|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|General Exam|3100,3104|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|General Exam|3110,3116|false|false|false|C1547311|Patient Condition Code - Stable|Stable
Anatomy|Body Location or Region|General Exam|3117,3126|false|false|false|C0000726|Abdomen|abdominal
Anatomy|Body Part, Organ, or Organ Component|General Exam|3127,3133|false|false|false|C0003483|Aorta|aortic
Event|Event|General Exam|3142,3155|false|false|false|||calcification
Finding|Organ or Tissue Function|General Exam|3142,3155|false|false|false|C0006660;C0006663;C1533591|Calcification;Calcinosis;Physiologic calcification|calcification
Finding|Pathologic Function|General Exam|3142,3155|false|false|false|C0006660;C0006663;C1533591|Calcification;Calcinosis;Physiologic calcification|calcification
Event|Event|General Exam|3156,3168|false|false|false|||displacement
Finding|Mental Process|General Exam|3156,3168|false|false|false|C0012725|Psychologic Displacement|displacement
Phenomenon|Phenomenon or Process|General Exam|3156,3168|false|false|false|C2347509|Physical Shift|displacement
Finding|Intellectual Product|General Exam|3174,3180|false|false|false|C1547311|Patient Condition Code - Stable|Stable
Anatomy|Body Part, Organ, or Organ Component|General Exam|3181,3186|false|false|false|C0022646|Kidney|renal
Disorder|Disease or Syndrome|General Exam|3181,3186|false|false|false|C0042075|Urologic Diseases|renal
Disorder|Disease or Syndrome|General Exam|3181,3192|false|false|false|C3887499|Renal cyst|renal cysts
Disorder|Anatomical Abnormality|General Exam|3187,3192|false|false|false|C0010709|Cyst|cysts
Event|Event|General Exam|3187,3192|false|false|false|||cysts
Finding|Functional Concept|General Exam|3219,3224|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|General Exam|3219,3230|false|false|false|C0227613|Right kidney|right renal
Anatomy|Body Part, Organ, or Organ Component|General Exam|3225,3230|false|false|false|C0022646|Kidney|renal
Disorder|Disease or Syndrome|General Exam|3225,3230|false|false|false|C0042075|Urologic Diseases|renal
Event|Event|General Exam|3232,3240|false|false|false|||calculus
Finding|Body Substance|General Exam|3232,3240|false|false|false|C0006736|Calculi|calculus
Procedure|Laboratory Procedure|General Exam|3232,3240|false|false|false|C3668917|Calculus (lab procedure)|calculus
Finding|Finding|General Exam|3246,3254|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|General Exam|3246,3254|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Disorder|Disease or Syndrome|General Exam|3255,3264|false|false|false|C0034067|Pulmonary Emphysema|emphysema
Event|Event|General Exam|3255,3264|false|false|false|||emphysema
Finding|Pathologic Function|General Exam|3255,3264|false|false|false|C0013990|Pathological accumulation of air in tissues|emphysema
Finding|Idea or Concept|Hospital Course|3295,3299|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|Hospital Course|3295,3299|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|Hospital Course|3300,3303|false|false|false|||old
Attribute|Clinical Attribute|Hospital Course|3315,3320|false|false|false|C1300072|Tumor stage|stage
Anatomy|Body Location or Region|Hospital Course|3324,3328|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|3324,3328|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Hospital Course|3324,3328|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Hospital Course|3324,3328|false|false|false|C0740941|Lung Problem|lung
Event|Event|Hospital Course|3329,3336|false|false|false|||adenoca
Disorder|Disease or Syndrome|Hospital Course|3338,3341|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|3338,3341|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|3338,3341|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Hospital Course|3338,3341|false|false|false|||CAD
Finding|Gene or Genome|Hospital Course|3338,3341|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|3338,3341|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|3338,3341|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3338,3341|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|Hospital Course|3346,3355|false|false|false|||presented
Event|Event|Hospital Course|3362,3367|false|false|false|||fever
Finding|Finding|Hospital Course|3362,3367|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|Hospital Course|3362,3367|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Finding|Hospital Course|3368,3375|false|false|false|C4534363|At home|at home
Event|Event|Hospital Course|3371,3375|false|false|false|||home
Finding|Idea or Concept|Hospital Course|3371,3375|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|3371,3375|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|3371,3375|false|false|false|C1553498|home health encounter|home
Finding|Finding|Hospital Course|3381,3386|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Finding|Sign or Symptom|Hospital Course|3381,3386|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Event|Event|Hospital Course|3392,3401|false|false|false|||presented
Event|Event|Hospital Course|3420,3427|false|false|false|||fatigue
Finding|Sign or Symptom|Hospital Course|3420,3427|false|false|false|C0015672|Fatigue|fatigue
Event|Event|Hospital Course|3429,3442|false|false|false|||nonproductive
Drug|Organic Chemical|Hospital Course|3444,3449|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|Hospital Course|3444,3449|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|Hospital Course|3444,3449|false|false|false|||cough
Finding|Sign or Symptom|Hospital Course|3444,3449|false|false|false|C0010200|Coughing|cough
Event|Event|Hospital Course|3458,3465|false|false|false|||chronic
Finding|Intellectual Product|Hospital Course|3458,3465|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Hospital Course|3458,3465|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Finding|Idea or Concept|Hospital Course|3473,3476|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|3473,3476|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|3480,3486|false|false|false|||fevers
Finding|Sign or Symptom|Hospital Course|3480,3486|false|false|false|C0015967|Fever|fevers
Anatomy|Body Location or Region|Hospital Course|3489,3494|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|Hospital Course|3489,3494|false|false|false|C0741025|Chest problem|Chest
Procedure|Diagnostic Procedure|Hospital Course|3489,3499|false|false|false|C0039985|Plain chest X-ray|Chest xray
Event|Event|Hospital Course|3495,3499|false|false|false|||xray
Phenomenon|Natural Phenomenon or Process|Hospital Course|3495,3499|false|false|false|C0043309|Roentgen Rays|xray
Procedure|Diagnostic Procedure|Hospital Course|3495,3499|false|false|false|C0043299|Diagnostic radiologic examination|xray
Event|Event|Hospital Course|3505,3517|false|false|false|||unremarkable
Event|Event|Hospital Course|3532,3536|false|false|false|||rule
Disorder|Disease or Syndrome|Hospital Course|3541,3550|false|true|true|C0009450|Communicable Diseases|infection
Event|Event|Hospital Course|3541,3550|false|false|false|||infection
Finding|Pathologic Function|Hospital Course|3541,3550|false|true|true|C3714514|Infection|infection
Anatomy|Body Location or Region|Hospital Course|3561,3569|false|false|false|C1515974|Anatomic Site|location
Finding|Intellectual Product|Hospital Course|3561,3569|false|true|false|C1555588|Transaction counts and value totals - location|location
Anatomy|Body Location or Region|Hospital Course|3578,3582|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|3578,3582|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Hospital Course|3578,3582|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Hospital Course|3578,3582|false|false|false|C0740941|Lung Problem|lung
Disorder|Neoplastic Process|Hospital Course|3578,3589|false|false|false|C0242379;C0684249|Carcinoma of lung;Malignant neoplasm of lung|lung cancer
Disorder|Neoplastic Process|Hospital Course|3583,3589|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Hospital Course|3583,3589|false|false|false|||cancer
Event|Event|Hospital Course|3600,3608|false|false|false|||negative
Finding|Classification|Hospital Course|3600,3608|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|3600,3608|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|3600,3608|false|false|false|C5237010|Expression Negative|negative
Disorder|Disease or Syndrome|Hospital Course|3609,3614|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Hospital Course|3609,3614|false|false|false|||blood
Finding|Body Substance|Hospital Course|3609,3614|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Body Substance|Hospital Course|3619,3624|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|Hospital Course|3619,3624|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|Hospital Course|3619,3624|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Event|Event|Hospital Course|3625,3633|false|false|false|||cultures
Finding|Idea or Concept|Hospital Course|3625,3633|false|false|false|C0010453|Culture (Anthropological)|cultures
Attribute|Clinical Attribute|Hospital Course|3651,3659|false|false|false|C0881858||CT chest
Procedure|Diagnostic Procedure|Hospital Course|3651,3659|false|false|false|C0202823|Chest CT|CT chest
Anatomy|Body Location or Region|Hospital Course|3654,3659|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|3654,3659|false|false|false|C0741025|Chest problem|chest
Event|Event|Hospital Course|3663,3672|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|3663,3672|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|Hospital Course|3695,3701|false|false|false|||repeat
Finding|Functional Concept|Hospital Course|3695,3701|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Procedure|Diagnostic Procedure|Hospital Course|3703,3710|false|false|false|C0040405|X-Ray Computed Tomography|CT scan
Event|Event|Hospital Course|3706,3710|false|false|false|||scan
Procedure|Diagnostic Procedure|Hospital Course|3706,3710|false|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Finding|Intellectual Product|Hospital Course|3725,3729|false|false|false|C1561540|Transaction counts and value totals - week|week
Attribute|Clinical Attribute|Hospital Course|3746,3754|false|false|false|C0881858||CT chest
Procedure|Diagnostic Procedure|Hospital Course|3746,3754|false|false|false|C0202823|Chest CT|CT chest
Anatomy|Body Location or Region|Hospital Course|3749,3754|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|3749,3754|false|false|false|C0741025|Chest problem|chest
Finding|Finding|Hospital Course|3777,3780|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Hospital Course|3777,3780|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Disorder|Disease or Syndrome|Hospital Course|3781,3791|false|false|false|C0009450|Communicable Diseases|infectious
Event|Event|Hospital Course|3781,3791|false|false|false|||infectious
Finding|Pathologic Function|Hospital Course|3781,3799|false|false|false|C0745283|INFECTIOUS PROCESS|infectious process
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|3792,3799|false|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|Hospital Course|3792,3799|false|false|false|C1951340|Process Pharmacologic Substance|process
Event|Event|Hospital Course|3792,3799|false|false|false|||process
Finding|Functional Concept|Hospital Course|3792,3799|false|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|Hospital Course|3792,3799|false|false|false|C1522240|Process|process
Finding|Functional Concept|Hospital Course|3807,3812|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Finding|Intellectual Product|Hospital Course|3824,3830|false|false|false|C1552826|Table Cell Vertical Align - middle|middle
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|3831,3836|false|false|false|C0796494|lobe|lobes
Finding|Finding|Hospital Course|3841,3845|false|false|false|C5575035|Well (answer to question)|well
Finding|Intellectual Product|Hospital Course|3849,3855|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|Hospital Course|3856,3861|false|false|false|||areas
Disorder|Disease or Syndrome|Hospital Course|3865,3878|false|false|false|C0521530|Lung consolidation|consolidation
Event|Event|Hospital Course|3865,3878|false|false|false|||consolidation
Event|Event|Hospital Course|3892,3902|false|false|false|||consistent
Finding|Idea or Concept|Hospital Course|3892,3902|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|Hospital Course|3892,3907|false|false|false|C0332290|Consistent with|consistent with
Disorder|Neoplastic Process|Hospital Course|3908,3934|false|false|false|C0007120|Bronchioloalveolar Adenocarcinoma|bronchioalveolar carcinoma
Disorder|Neoplastic Process|Hospital Course|3925,3934|false|false|false|C0007097|Carcinoma|carcinoma
Event|Event|Hospital Course|3925,3934|false|false|false|||carcinoma
Event|Event|Hospital Course|3946,3953|false|false|false|||started
Drug|Antibiotic|Hospital Course|3957,3968|false|false|false|C0007561|ceftriaxone|ceftriaxone
Drug|Organic Chemical|Hospital Course|3957,3968|false|false|false|C0007561|ceftriaxone|ceftriaxone
Event|Event|Hospital Course|3957,3968|false|false|false|||ceftriaxone
Drug|Antibiotic|Hospital Course|3973,3985|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|Hospital Course|3973,3985|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|Hospital Course|3973,3985|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Event|Event|Hospital Course|3973,3985|false|false|false|||azithromycin
Event|Event|Hospital Course|3994,4004|false|false|false|||discharged
Drug|Antibiotic|Hospital Course|4009,4019|false|false|false|C0007562|cefuroxime|cefuroxime
Drug|Organic Chemical|Hospital Course|4009,4019|false|false|false|C0007562|cefuroxime|cefuroxime
Event|Event|Hospital Course|4009,4019|false|false|false|||cefuroxime
Drug|Antibiotic|Hospital Course|4024,4036|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|Hospital Course|4024,4036|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|Hospital Course|4024,4036|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Event|Event|Hospital Course|4024,4036|false|false|false|||azithromycin
Event|Event|Hospital Course|4052,4062|false|false|false|||discharged
Event|Event|Hospital Course|4066,4070|false|false|false|||home
Finding|Idea or Concept|Hospital Course|4066,4070|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|4066,4070|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|4066,4070|false|false|false|C1553498|home health encounter|home
Drug|Biologically Active Substance|Hospital Course|4072,4078|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|Hospital Course|4072,4078|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|Hospital Course|4072,4078|false|false|false|C0030054|oxygen|oxygen
Event|Event|Hospital Course|4072,4078|false|false|false|||oxygen
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4072,4078|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Drug|Biologically Active Substance|Hospital Course|4097,4103|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|Hospital Course|4097,4103|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|Hospital Course|4097,4103|false|false|false|C0030054|oxygen|oxygen
Event|Event|Hospital Course|4097,4103|false|false|false|||oxygen
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4097,4103|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Event|Event|Hospital Course|4104,4113|false|false|false|||sometimes
Finding|Finding|Hospital Course|4114,4121|false|false|false|C4534363|At home|at home
Event|Event|Hospital Course|4117,4121|false|false|false|||home
Finding|Idea or Concept|Hospital Course|4117,4121|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|4117,4121|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|4117,4121|false|false|false|C1553498|home health encounter|home
Event|Event|Hospital Course|4131,4141|false|false|false|||instructed
Event|Event|Hospital Course|4145,4148|false|false|false|||use
Finding|Finding|Hospital Course|4152,4161|false|false|false|C0682295|Full-time employment (finding)|full-time
Finding|Finding|Hospital Course|4157,4161|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Hospital Course|4157,4161|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Hospital Course|4157,4161|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|Hospital Course|4168,4177|false|false|false|||discharge
Finding|Body Substance|Hospital Course|4168,4177|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|4168,4177|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|4168,4177|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|4168,4177|false|false|false|C0030685|Patient Discharge|discharge
Finding|Intellectual Product|Hospital Course|4184,4189|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Disorder|Disease or Syndrome|Hospital Course|4184,4203|false|false|false|C0022660|Kidney Failure, Acute|Acute renal failure
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4190,4195|false|false|false|C0022646|Kidney|renal
Disorder|Disease or Syndrome|Hospital Course|4190,4195|false|false|false|C0042075|Urologic Diseases|renal
Disorder|Disease or Syndrome|Hospital Course|4190,4203|false|false|false|C0035078|Kidney Failure|renal failure
Event|Event|Hospital Course|4196,4203|false|false|false|||failure
Finding|Functional Concept|Hospital Course|4196,4203|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|Hospital Course|4196,4203|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|Hospital Course|4196,4203|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Drug|Biologically Active Substance|Hospital Course|4225,4235|false|false|false|C0010294|creatinine|creatinine
Drug|Organic Chemical|Hospital Course|4225,4235|false|false|false|C0010294|creatinine|creatinine
Event|Event|Hospital Course|4225,4235|false|false|false|||creatinine
Finding|Physiologic Function|Hospital Course|4225,4235|false|false|false|C4551889|Creatinine metabolic function|creatinine
Procedure|Laboratory Procedure|Hospital Course|4225,4235|false|false|false|C0201975|Creatinine measurement|creatinine
Event|Event|Hospital Course|4240,4249|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|4240,4249|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Drug|Biomedical or Dental Material|Hospital Course|4271,4279|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|Hospital Course|4271,4279|false|false|false|||baseline
Finding|Idea or Concept|Hospital Course|4271,4279|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|Hospital Course|4303,4307|false|false|false|||felt
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4314,4322|false|false|false|C1550297|Prerenal|prerenal
Disorder|Disease or Syndrome|Hospital Course|4314,4331|false|false|false|C0554309|Prerenal azotemia|prerenal azotemia
Disorder|Disease or Syndrome|Hospital Course|4323,4331|false|false|false|C0242528;C0554309|Azotemia;Prerenal azotemia|azotemia
Event|Event|Hospital Course|4323,4331|false|false|false|||azotemia
Event|Event|Hospital Course|4339,4347|false|false|false|||improved
Event|Event|Hospital Course|4356,4365|false|false|false|||hydration
Finding|Finding|Hospital Course|4356,4365|false|false|false|C1321013;C4520800|Hydration;Hydration status|hydration
Finding|Physiologic Function|Hospital Course|4356,4365|false|false|false|C1321013;C4520800|Hydration;Hydration status|hydration
Disorder|Disease or Syndrome|Hospital Course|4382,4387|false|false|false|C1410088|Still|still
Finding|Finding|Hospital Course|4392,4395|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Hospital Course|4392,4395|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4396,4401|false|false|false|C0022646|Kidney|renal
Disorder|Disease or Syndrome|Hospital Course|4396,4401|false|false|false|C0042075|Urologic Diseases|renal
Disorder|Disease or Syndrome|Hospital Course|4396,4415|false|false|false|C0035078;C1565489|Kidney Failure;Renal Insufficiency|renal insufficiency
Event|Event|Hospital Course|4402,4415|false|false|false|||insufficiency
Finding|Functional Concept|Hospital Course|4402,4415|false|false|false|C0231179|Insufficiency|insufficiency
Finding|Finding|Hospital Course|4426,4432|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|4426,4432|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|Hospital Course|4434,4441|false|false|false|||benefit
Event|Event|Hospital Course|4447,4453|false|false|false|||follow
Finding|Functional Concept|Hospital Course|4447,4453|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|Hospital Course|4447,4453|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|Hospital Course|4447,4456|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|Hospital Course|4447,4456|false|false|false|C1522577|follow-up|follow-up
Event|Event|Hospital Course|4454,4456|false|false|false|||up
Event|Event|Hospital Course|4462,4472|false|false|false|||nephrology
Event|Event|Hospital Course|4479,4488|false|false|false|||discharge
Finding|Body Substance|Hospital Course|4479,4488|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|4479,4488|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|4479,4488|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|4479,4488|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|Hospital Course|4505,4515|false|false|false|||instructed
Event|Event|Hospital Course|4519,4525|false|false|false|||follow
Finding|Finding|Hospital Course|4528,4531|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Hospital Course|4528,4531|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Finding|Hospital Course|4528,4541|false|false|false|C0860866|Potassium low|low potassium
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4528,4546|false|false|false|C0452349|Potassium restricted diet|low potassium diet
Drug|Biologically Active Substance|Hospital Course|4532,4541|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Element, Ion, or Isotope|Hospital Course|4532,4541|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Food|Hospital Course|4532,4541|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Inorganic Chemical|Hospital Course|4532,4541|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Pharmacologic Substance|Hospital Course|4532,4541|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Event|Event|Hospital Course|4532,4541|false|false|false|||potassium
Finding|Physiologic Function|Hospital Course|4532,4541|false|false|false|C4553027|Potassium metabolic function|potassium
Procedure|Laboratory Procedure|Hospital Course|4532,4541|false|false|false|C0202194|Potassium measurement|potassium
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4532,4546|false|false|false|C0301596|Potassium diet|potassium diet
Drug|Food|Hospital Course|4542,4546|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|Hospital Course|4542,4546|false|false|false|||diet
Finding|Functional Concept|Hospital Course|4542,4546|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|Hospital Course|4542,4546|false|false|false|C0012159|Diet therapy|diet
Disorder|Disease or Syndrome|Hospital Course|4552,4564|false|false|false|C0020625|Hyponatremia|Hyponatremia
Finding|Finding|Hospital Course|4574,4577|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Hospital Course|4574,4577|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Drug|Indicator, Reagent, or Diagnostic Aid|Hospital Course|4578,4583|false|false|false|C5575602|Cell Culture Serum|serum
Finding|Body Substance|Hospital Course|4578,4583|false|false|false|C0229671;C1546774;C1550100|Serum;Serum specimen|serum
Finding|Intellectual Product|Hospital Course|4578,4583|false|false|false|C0229671;C1546774;C1550100|Serum;Serum specimen|serum
Lab|Laboratory or Test Result|Hospital Course|4578,4590|false|false|false|C0587356|Serum sodium level|serum sodium
Procedure|Laboratory Procedure|Hospital Course|4578,4590|false|false|false|C0523891|Serum sodium measurement|serum sodium
Drug|Biologically Active Substance|Hospital Course|4584,4590|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|Hospital Course|4584,4590|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|Hospital Course|4584,4590|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Event|Event|Hospital Course|4584,4590|false|false|false|||sodium
Finding|Physiologic Function|Hospital Course|4584,4590|false|false|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|Hospital Course|4584,4590|false|false|false|C0337443|Sodium measurement|sodium
Event|Event|Hospital Course|4594,4603|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|4594,4603|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|Hospital Course|4605,4609|false|false|false|||felt
Drug|Organic Chemical|Hospital Course|4617,4624|false|false|false|C0163712|Relate - vinyl resin|related
Event|Event|Hospital Course|4617,4624|false|false|false|||related
Finding|Finding|Hospital Course|4617,4624|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|Hospital Course|4617,4624|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Event|Event|Hospital Course|4628,4639|false|false|false|||hypovolemia
Finding|Finding|Hospital Course|4628,4639|false|true|false|C0546884|Hypovolemia|hypovolemia
Finding|Mental Process|Hospital Course|4647,4654|false|false|false|C0542559|contextual factors|setting
Event|Event|Hospital Course|4662,4669|false|false|false|||illness
Finding|Sign or Symptom|Hospital Course|4662,4669|false|false|false|C0221423|Illness (finding)|illness
Drug|Biologically Active Substance|Hospital Course|4677,4683|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|Hospital Course|4677,4683|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|Hospital Course|4677,4683|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Event|Event|Hospital Course|4677,4683|false|false|false|||sodium
Finding|Physiologic Function|Hospital Course|4677,4683|false|false|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|Hospital Course|4677,4683|false|false|false|C0337443|Sodium measurement|sodium
Event|Event|Hospital Course|4684,4692|false|false|false|||improved
Event|Event|Hospital Course|4703,4709|false|false|false|||levels
Drug|Substance|Hospital Course|4718,4724|false|false|false|C0302908|Liquid substance|fluids
Event|Event|Hospital Course|4718,4724|false|false|false|||fluids
Finding|Body Substance|Hospital Course|4718,4724|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4718,4724|false|false|false|C0016286|Fluid Therapy|fluids
Attribute|Clinical Attribute|Hospital Course|4730,4735|false|false|false|C1300072|Tumor stage|Stage
Finding|Intellectual Product|Hospital Course|4730,4738|false|false|false|C0441772|Stage level 4|Stage IV
Disorder|Neoplastic Process|Hospital Course|4730,4758|false|false|false|C0854988|Adenocarcinoma of lung, stage IV|Stage IV Lung Adenocarcinoma
Anatomy|Body Location or Region|Hospital Course|4739,4743|false|false|false|C0024109;C4037972|Chest>Lung;Lung|Lung
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4739,4743|false|false|false|C0024109;C4037972|Chest>Lung;Lung|Lung
Disorder|Disease or Syndrome|Hospital Course|4739,4743|false|false|false|C0024115|Lung diseases|Lung
Finding|Finding|Hospital Course|4739,4743|false|false|false|C0740941|Lung Problem|Lung
Disorder|Neoplastic Process|Hospital Course|4739,4758|false|false|false|C0152013|Adenocarcinoma of lung (disorder)|Lung Adenocarcinoma
Disorder|Neoplastic Process|Hospital Course|4744,4758|false|false|false|C0001418;C5551397|Adenocarcinoma;Malignant adenomatous neoplasm|Adenocarcinoma
Event|Event|Hospital Course|4744,4758|false|false|false|||Adenocarcinoma
Event|Event|Hospital Course|4773,4779|false|false|false|||cycles
Drug|Organic Chemical|Hospital Course|4784,4794|false|false|false|C0210657|pemetrexed|pemetrexed
Drug|Pharmacologic Substance|Hospital Course|4784,4794|false|false|false|C0210657|pemetrexed|pemetrexed
Event|Event|Hospital Course|4784,4794|false|false|false|||pemetrexed
Event|Event|Hospital Course|4808,4814|false|false|false|||follow
Event|Event|Hospital Course|4859,4868|false|false|false|||treatment
Finding|Conceptual Entity|Hospital Course|4859,4868|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Hospital Course|4859,4868|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Hospital Course|4859,4868|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4859,4868|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Disorder|Disease or Syndrome|Hospital Course|4874,4880|false|false|false|C0002871|Anemia|Anemia
Event|Event|Hospital Course|4874,4880|false|false|false|||Anemia
Event|Event|Hospital Course|4890,4895|false|false|false|||given
Event|Event|Hospital Course|4898,4902|false|false|false|||unit
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4906,4911|false|false|false|C2316467|Packed red blood cells|PRBCs
Drug|Pharmacologic Substance|Hospital Course|4906,4911|false|false|false|C2316467|Packed red blood cells|PRBCs
Event|Event|Hospital Course|4906,4911|false|false|false|||PRBCs
Disorder|Disease or Syndrome|Hospital Course|4916,4922|false|false|false|C0002871|Anemia|anemia
Event|Event|Hospital Course|4916,4922|false|false|false|||anemia
Event|Event|Hospital Course|4927,4936|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|4927,4936|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Disorder|Disease or Syndrome|Hospital Course|4943,4949|false|false|false|C0002871|Anemia|anemia
Event|Event|Hospital Course|4943,4949|false|false|false|||anemia
Event|Event|Hospital Course|4954,4958|false|false|false|||felt
Drug|Organic Chemical|Hospital Course|4965,4972|false|false|false|C0163712|Relate - vinyl resin|related
Event|Event|Hospital Course|4965,4972|false|false|false|||related
Finding|Finding|Hospital Course|4965,4972|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|Hospital Course|4965,4972|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Event|Event|Hospital Course|4988,5000|false|false|false|||chemotherapy
Finding|Functional Concept|Hospital Course|4988,5000|false|false|false|C0013217|pharmacotherapeutic|chemotherapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4988,5000|false|false|false|C0013216;C0392920;C3665472|Chemotherapy;Chemotherapy Regimen;Pharmacotherapy|chemotherapy
Disorder|Disease or Syndrome|Hospital Course|5006,5009|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5006,5009|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|5006,5009|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Hospital Course|5006,5009|false|false|false|||CAD
Finding|Gene or Genome|Hospital Course|5006,5009|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|5006,5009|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|5006,5009|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5006,5009|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|Hospital Course|5019,5028|false|false|false|||continued
Drug|Organic Chemical|Hospital Course|5034,5040|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|statin
Drug|Pharmacologic Substance|Hospital Course|5034,5040|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|statin
Event|Event|Hospital Course|5034,5040|false|false|false|||statin
Finding|Gene or Genome|Hospital Course|5034,5040|false|false|false|C1414273|EEF1A2 gene|statin
Drug|Organic Chemical|Hospital Course|5042,5049|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|Hospital Course|5042,5049|false|false|false|C0004057|aspirin|aspirin
Event|Event|Hospital Course|5042,5049|false|false|false|||aspirin
Drug|Organic Chemical|Hospital Course|5055,5066|false|false|false|C0070166|clopidogrel|clopidogrel
Drug|Pharmacologic Substance|Hospital Course|5055,5066|false|false|false|C0070166|clopidogrel|clopidogrel
Event|Event|Hospital Course|5055,5066|false|false|false|||clopidogrel
Disorder|Disease or Syndrome|Hospital Course|5072,5075|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|Hospital Course|5072,5075|false|false|false|||HTN
Event|Event|Hospital Course|5085,5094|false|false|false|||continued
Drug|Organic Chemical|Hospital Course|5098,5108|false|false|false|C0051696|amlodipine|amlodipine
Drug|Pharmacologic Substance|Hospital Course|5098,5108|false|false|false|C0051696|amlodipine|amlodipine
Event|Event|Hospital Course|5098,5108|false|false|false|||amlodipine
Attribute|Clinical Attribute|Hospital Course|5112,5123|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|5112,5123|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|5112,5123|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|5112,5123|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|5112,5136|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|5127,5136|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|5127,5136|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Organic Chemical|Hospital Course|5138,5148|false|false|false|C0051696|amlodipine|amlodipine
Drug|Pharmacologic Substance|Hospital Course|5138,5148|false|false|false|C0051696|amlodipine|amlodipine
Drug|Organic Chemical|Hospital Course|5160,5172|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|Hospital Course|5160,5172|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|Hospital Course|5160,5172|false|false|false|||atorvastatin
Drug|Organic Chemical|Hospital Course|5185,5196|false|false|false|C0070166|clopidogrel|clopidogrel
Drug|Pharmacologic Substance|Hospital Course|5185,5196|false|false|false|C0070166|clopidogrel|clopidogrel
Event|Event|Hospital Course|5185,5196|false|false|false|||clopidogrel
Drug|Organic Chemical|Hospital Course|5209,5216|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|Hospital Course|5209,5216|false|false|false|C0004057|aspirin|aspirin
Event|Event|Hospital Course|5209,5216|false|false|false|||aspirin
Drug|Organic Chemical|Hospital Course|5229,5239|false|false|false|C0034665|ranitidine|ranitidine
Drug|Pharmacologic Substance|Hospital Course|5229,5239|false|false|false|C0034665|ranitidine|ranitidine
Event|Event|Hospital Course|5229,5239|false|false|false|||ranitidine
Drug|Organic Chemical|Hospital Course|5253,5259|false|false|false|C0178638|folate|folate
Drug|Pharmacologic Substance|Hospital Course|5253,5259|false|false|false|C0178638|folate|folate
Drug|Vitamin|Hospital Course|5253,5259|false|false|false|C0178638|folate|folate
Event|Event|Hospital Course|5253,5259|false|false|false|||folate
Procedure|Laboratory Procedure|Hospital Course|5253,5259|false|false|false|C0523631|Folic acid measurement|folate
Drug|Organic Chemical|Hospital Course|5260,5270|false|false|false|C0023992|loperamide|loperamide
Drug|Pharmacologic Substance|Hospital Course|5260,5270|false|false|false|C0023992|loperamide|loperamide
Finding|Gene or Genome|Hospital Course|5271,5274|false|false|false|C1422467|CIAO3 gene|prn
Drug|Organic Chemical|Hospital Course|5275,5284|false|false|false|C0024002|lorazepam|lorazepam
Drug|Pharmacologic Substance|Hospital Course|5275,5284|false|false|false|C0024002|lorazepam|lorazepam
Finding|Gene or Genome|Hospital Course|5285,5288|false|false|false|C1422467|CIAO3 gene|prn
Drug|Organic Chemical|Hospital Course|5289,5303|false|false|false|C0025853|metoclopramide|metoclopramide
Drug|Pharmacologic Substance|Hospital Course|5289,5303|false|false|false|C0025853|metoclopramide|metoclopramide
Finding|Gene or Genome|Hospital Course|5304,5307|false|false|false|C1422467|CIAO3 gene|prn
Drug|Organic Chemical|Hospital Course|5308,5319|false|false|false|C0061851|ondansetron|ondansetron
Drug|Pharmacologic Substance|Hospital Course|5308,5319|false|false|false|C0061851|ondansetron|ondansetron
Finding|Gene or Genome|Hospital Course|5320,5323|false|false|false|C1422467|CIAO3 gene|prn
Drug|Organic Chemical|Hospital Course|5324,5333|false|false|false|C0040805|trazodone|trazodone
Drug|Pharmacologic Substance|Hospital Course|5324,5333|false|false|false|C0040805|trazodone|trazodone
Event|Event|Hospital Course|5324,5333|false|false|false|||trazodone
Finding|Gene or Genome|Hospital Course|5346,5349|false|false|false|C1422467|CIAO3 gene|prn
Event|Event|Hospital Course|5353,5362|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|5353,5362|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|5353,5362|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|5353,5362|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|5353,5362|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|5353,5374|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|5363,5374|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|5363,5374|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|5363,5374|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|5363,5374|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|5379,5389|false|false|false|C0051696|amlodipine|Amlodipine
Drug|Pharmacologic Substance|Hospital Course|5379,5389|false|false|false|C0051696|amlodipine|Amlodipine
Drug|Biomedical or Dental Material|Hospital Course|5395,5401|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|5415,5421|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|5415,5421|false|false|false|||Tablet
Drug|Organic Chemical|Hospital Course|5446,5458|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|5446,5458|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Biomedical or Dental Material|Hospital Course|5465,5471|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|5472,5475|false|false|false|||Sig
Drug|Biomedical or Dental Material|Hospital Course|5485,5491|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|5485,5491|false|false|false|||Tablet
Event|Event|Hospital Course|5492,5494|false|false|false|||PO
Finding|Intellectual Product|Hospital Course|5495,5499|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|5495,5505|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|Hospital Course|5502,5505|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|5502,5505|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|5513,5524|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Pharmacologic Substance|Hospital Course|5513,5524|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Biomedical or Dental Material|Hospital Course|5531,5537|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|5551,5557|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|5551,5557|false|false|false|||Tablet
Drug|Organic Chemical|Hospital Course|5582,5589|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Hospital Course|5582,5589|false|false|false|C0004057|aspirin|Aspirin
Drug|Biomedical or Dental Material|Hospital Course|5596,5602|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|5596,5612|false|false|false|C0304290|Chewable Tablet|Tablet, Chewable
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5613,5616|false|false|false|C0262329|Short insular gyrus|Sig
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5613,5616|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Immunologic Factor|Hospital Course|5613,5616|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Finding|Receptor|Hospital Course|5613,5616|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Biomedical or Dental Material|Hospital Course|5626,5632|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|5626,5632|false|false|false|||Tablet
Drug|Biomedical or Dental Material|Hospital Course|5626,5642|false|false|false|C0304290|Chewable Tablet|Tablet, Chewable
Event|Event|Hospital Course|5634,5642|false|false|false|||Chewable
Drug|Organic Chemical|Hospital Course|5667,5677|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Pharmacologic Substance|Hospital Course|5667,5677|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Organic Chemical|Hospital Course|5667,5681|false|false|false|C0700466|ranitidine hydrochloride|Ranitidine HCl
Drug|Pharmacologic Substance|Hospital Course|5667,5681|false|false|false|C0700466|ranitidine hydrochloride|Ranitidine HCl
Disorder|Neoplastic Process|Hospital Course|5678,5681|false|false|false|C0023443|Hairy Cell Leukemia|HCl
Drug|Immunologic Factor|Hospital Course|5678,5681|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Inorganic Chemical|Hospital Course|5678,5681|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Pharmacologic Substance|Hospital Course|5678,5681|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Event|Event|Hospital Course|5678,5681|false|false|false|||HCl
Drug|Biomedical or Dental Material|Hospital Course|5689,5695|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|5709,5715|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|5709,5715|false|false|false|||Tablet
Drug|Organic Chemical|Hospital Course|5740,5750|false|false|false|C0016410|folic acid|Folic Acid
Drug|Pharmacologic Substance|Hospital Course|5740,5750|false|false|false|C0016410|folic acid|Folic Acid
Drug|Vitamin|Hospital Course|5740,5750|false|false|false|C0016410|folic acid|Folic Acid
Procedure|Laboratory Procedure|Hospital Course|5740,5750|false|false|false|C0523631|Folic acid measurement|Folic Acid
Event|Event|Hospital Course|5746,5750|false|false|false|||Acid
Drug|Biomedical or Dental Material|Hospital Course|5756,5762|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|5763,5766|false|false|false|||Sig
Drug|Biomedical or Dental Material|Hospital Course|5776,5782|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|5776,5782|false|false|false|||Tablet
Drug|Organic Chemical|Hospital Course|5807,5817|false|false|false|C0023992|loperamide|Loperamide
Drug|Pharmacologic Substance|Hospital Course|5807,5817|false|false|false|C0023992|loperamide|Loperamide
Drug|Biomedical or Dental Material|Hospital Course|5823,5829|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|5830,5833|false|false|false|||Sig
Drug|Biomedical or Dental Material|Hospital Course|5843,5849|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|5843,5849|false|false|false|||Tablet
Disorder|Disease or Syndrome|Hospital Course|5858,5863|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|Hospital Course|5867,5870|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|5867,5870|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|5874,5880|false|false|false|||needed
Event|Event|Hospital Course|5885,5893|false|false|false|||diarrhea
Finding|Finding|Hospital Course|5885,5893|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|Hospital Course|5885,5893|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Drug|Organic Chemical|Hospital Course|5900,5909|false|false|false|C0024002|lorazepam|Lorazepam
Drug|Pharmacologic Substance|Hospital Course|5900,5909|false|false|false|C0024002|lorazepam|Lorazepam
Event|Event|Hospital Course|5900,5909|false|false|false|||Lorazepam
Anatomy|Body Space or Junction|Hospital Course|5911,5915|false|false|false|C0226896|Oral cavity|Oral
Drug|Biomedical or Dental Material|Hospital Course|5911,5915|false|false|false|C1272919|Oral Dosage Form|Oral
Finding|Finding|Hospital Course|5911,5915|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Finding|Functional Concept|Hospital Course|5911,5915|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Drug|Organic Chemical|Hospital Course|5919,5933|false|false|false|C0025853|metoclopramide|Metoclopramide
Drug|Pharmacologic Substance|Hospital Course|5919,5933|false|false|false|C0025853|metoclopramide|Metoclopramide
Event|Event|Hospital Course|5919,5933|false|false|false|||Metoclopramide
Anatomy|Body Space or Junction|Hospital Course|5935,5939|false|false|false|C0226896|Oral cavity|Oral
Drug|Biomedical or Dental Material|Hospital Course|5935,5939|false|false|false|C1272919|Oral Dosage Form|Oral
Event|Event|Hospital Course|5935,5939|false|false|false|||Oral
Finding|Finding|Hospital Course|5935,5939|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Finding|Functional Concept|Hospital Course|5935,5939|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Drug|Organic Chemical|Hospital Course|5944,5950|false|false|false|C0206046|Zofran|Zofran
Drug|Pharmacologic Substance|Hospital Course|5944,5950|false|false|false|C0206046|Zofran|Zofran
Anatomy|Body Space or Junction|Hospital Course|5952,5956|false|false|false|C0226896|Oral cavity|Oral
Drug|Biomedical or Dental Material|Hospital Course|5952,5956|false|false|false|C1272919|Oral Dosage Form|Oral
Finding|Finding|Hospital Course|5952,5956|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Finding|Functional Concept|Hospital Course|5952,5956|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Drug|Organic Chemical|Hospital Course|5961,5970|false|false|false|C0040805|trazodone|Trazodone
Drug|Pharmacologic Substance|Hospital Course|5961,5970|false|false|false|C0040805|trazodone|Trazodone
Drug|Biomedical or Dental Material|Hospital Course|5977,5983|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|5997,6003|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|6004,6006|false|false|false|||PO
Event|Event|Hospital Course|6022,6028|false|false|false|||needed
Drug|Pharmacologic Substance|Hospital Course|6033,6041|false|false|false|C1950154|Insomnia homeopathic medication|insomnia
Event|Event|Hospital Course|6033,6041|false|false|false|||insomnia
Finding|Sign or Symptom|Hospital Course|6033,6041|false|false|false|C0917801|Sleeplessness|insomnia
Drug|Antibiotic|Hospital Course|6049,6061|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Drug|Clinical Drug|Hospital Course|6049,6061|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Drug|Organic Chemical|Hospital Course|6049,6061|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Drug|Biomedical or Dental Material|Hospital Course|6069,6075|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|6089,6095|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|6089,6095|false|false|false|||Tablet
Event|Event|Hospital Course|6099,6103|false|false|false|||Q24H
Event|Event|Hospital Course|6140,6144|false|false|false|||dose
Drug|Biomedical or Dental Material|Hospital Course|6161,6167|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|6161,6167|false|false|false|||Tablet
Finding|Idea or Concept|Hospital Course|6172,6179|false|false|false|C0807726|refill|Refills
Drug|Antibiotic|Hospital Course|6188,6198|false|false|false|C0007562|cefuroxime|Cefuroxime
Drug|Organic Chemical|Hospital Course|6188,6198|false|false|false|C0007562|cefuroxime|Cefuroxime
Event|Event|Hospital Course|6188,6198|false|false|false|||Cefuroxime
Drug|Antibiotic|Hospital Course|6188,6205|false|false|false|C0055015|cefuroxime axetil|Cefuroxime Axetil
Drug|Organic Chemical|Hospital Course|6188,6205|false|false|false|C0055015|cefuroxime axetil|Cefuroxime Axetil
Drug|Biomedical or Dental Material|Hospital Course|6213,6219|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|6233,6239|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|6252,6255|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|6252,6255|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|6274,6278|false|false|false|||dose
Drug|Antibiotic|Hospital Course|6309,6319|false|false|false|C0003232|Antibiotics|antibiotic
Event|Event|Hospital Course|6309,6319|false|false|false|||antibiotic
Event|Event|Hospital Course|6327,6337|false|false|false|||completion
Drug|Biomedical or Dental Material|Hospital Course|6348,6354|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|6359,6366|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|6375,6380|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|Hospital Course|6375,6380|false|false|false|C3489575|sennosides, USP|Senna
Drug|Biomedical or Dental Material|Hospital Course|6388,6394|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|6408,6414|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|6426,6429|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|6426,6429|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|6434,6440|false|false|false|||needed
Event|Event|Hospital Course|6445,6457|false|false|false|||constipation
Finding|Sign or Symptom|Hospital Course|6445,6457|false|false|false|C0009806|Constipation|constipation
Drug|Organic Chemical|Hospital Course|6465,6475|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|Hospital Course|6465,6475|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|Hospital Course|6465,6484|false|false|false|C0700548|metoprolol tartrate|Metoprolol Tartrate
Drug|Pharmacologic Substance|Hospital Course|6465,6484|false|false|false|C0700548|metoprolol tartrate|Metoprolol Tartrate
Drug|Organic Chemical|Hospital Course|6476,6484|false|false|false|C0039328;C0144544|Tartrates;tartrate|Tartrate
Drug|Pharmacologic Substance|Hospital Course|6476,6484|false|false|false|C0039328;C0144544|Tartrates;tartrate|Tartrate
Event|Event|Hospital Course|6476,6484|false|false|false|||Tartrate
Drug|Biomedical or Dental Material|Hospital Course|6491,6497|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|6511,6517|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|6511,6517|false|false|false|||Tablet
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6521,6524|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6521,6524|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|6521,6524|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|6521,6524|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|6521,6524|false|false|false|C1332410|BID gene|BID
Finding|Finding|Hospital Course|6527,6534|false|false|false|C4035627|2 times|2 times
Disorder|Disease or Syndrome|Hospital Course|6529,6534|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|Hospital Course|6537,6540|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|6537,6540|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biomedical or Dental Material|Hospital Course|6549,6561|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Drug|Organic Chemical|Hospital Course|6549,6561|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Drug|Organic Chemical|Hospital Course|6549,6568|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Pharmacologic Substance|Hospital Course|6549,6568|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Organic Chemical|Hospital Course|6549,6573|false|false|false|C0724672|polyethylene glycol 3350|Polyethylene Glycol 3350
Drug|Pharmacologic Substance|Hospital Course|6549,6573|false|false|false|C0724672|polyethylene glycol 3350|Polyethylene Glycol 3350
Drug|Hazardous or Poisonous Substance|Hospital Course|6562,6568|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Drug|Organic Chemical|Hospital Course|6562,6568|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Event|Event|Hospital Course|6562,6568|false|false|false|||Glycol
Drug|Biomedical or Dental Material|Hospital Course|6587,6593|false|false|false|C0032861;C1382110|Powder dose form;powder physical state|Powder
Drug|Substance|Hospital Course|6587,6593|false|false|false|C0032861;C1382110|Powder dose form;powder physical state|Powder
Event|Event|Hospital Course|6587,6593|false|false|false|||Powder
Event|Event|Hospital Course|6594,6597|false|false|false|||Sig
Event|Event|Hospital Course|6629,6635|false|false|false|||needed
Event|Event|Hospital Course|6640,6652|false|false|false|||constipation
Finding|Sign or Symptom|Hospital Course|6640,6652|false|false|false|C0009806|Constipation|constipation
Event|Event|Hospital Course|6658,6667|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|6658,6667|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|6658,6667|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|6658,6667|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|6658,6667|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|6658,6679|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|6658,6679|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|6668,6679|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|6668,6679|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|6668,6679|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|Hospital Course|6681,6685|false|false|false|||Home
Finding|Idea or Concept|Hospital Course|6681,6685|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|6681,6685|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|6681,6685|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|Hospital Course|6691,6698|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|Hospital Course|6691,6698|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|Hospital Course|6701,6709|false|false|false|||Facility
Finding|Intellectual Product|Hospital Course|6701,6709|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|Hospital Course|6718,6727|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|6718,6727|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|6718,6727|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|6718,6727|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|6718,6727|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|6718,6737|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|6728,6737|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|6728,6737|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|6728,6737|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|6728,6737|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|6728,6737|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Disease or Syndrome|Principle Diagnosis|6758,6786|false|false|false|C0694549|Community-Acquired Pneumonia|Community-Acquired Pneumonia
Disorder|Disease or Syndrome|Principle Diagnosis|6777,6786|false|false|false|C0032285|Pneumonia|Pneumonia
Event|Event|Principle Diagnosis|6777,6786|false|false|false|||Pneumonia
Disorder|Neoplastic Process|Principle Diagnosis|6788,6797|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Event|Event|Principle Diagnosis|6788,6797|false|false|false|||Secondary
Finding|Functional Concept|Principle Diagnosis|6788,6797|false|false|false|C1522484|metastatic qualifier|Secondary
Attribute|Clinical Attribute|Principle Diagnosis|6788,6807|false|false|false|C4255018||Secondary Diagnosis
Finding|Finding|Principle Diagnosis|6788,6807|false|false|false|C0332138|Secondary diagnosis|Secondary Diagnosis
Attribute|Clinical Attribute|Principle Diagnosis|6798,6807|false|false|false|C0945731||Diagnosis
Event|Event|Principle Diagnosis|6798,6807|false|false|false|||Diagnosis
Finding|Classification|Principle Diagnosis|6798,6807|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Principle Diagnosis|6798,6807|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Principle Diagnosis|6798,6807|false|false|false|C0011900|Diagnosis|Diagnosis
Anatomy|Cell|Principle Diagnosis|6819,6823|false|false|false|C0007634|Cells|cell
Finding|Gene or Genome|Principle Diagnosis|6819,6823|false|false|false|C1413336;C1413337|CEL gene;CELP gene|cell
Anatomy|Body Location or Region|Principle Diagnosis|6824,6828|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|6824,6828|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Principle Diagnosis|6824,6828|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Principle Diagnosis|6824,6828|false|false|false|C0740941|Lung Problem|lung
Disorder|Neoplastic Process|Principle Diagnosis|6824,6835|false|false|false|C0242379;C0684249|Carcinoma of lung;Malignant neoplasm of lung|lung cancer
Disorder|Neoplastic Process|Principle Diagnosis|6829,6835|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Principle Diagnosis|6829,6835|false|false|false|||cancer
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|6836,6844|false|false|false|C0018787|Heart|Coronary
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|6836,6851|false|false|false|C0205042|Coronary artery|Coronary Artery
Disorder|Disease or Syndrome|Principle Diagnosis|6836,6859|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|Coronary Artery Disease
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|6845,6851|false|false|false|C0003842;C0226004|Arterial system;Arteries|Artery
Anatomy|Body System|Principle Diagnosis|6845,6851|false|false|false|C0003842;C0226004|Arterial system;Arteries|Artery
Disorder|Disease or Syndrome|Principle Diagnosis|6845,6859|false|false|false|C0852949|Arteriopathic disease|Artery Disease
Disorder|Disease or Syndrome|Principle Diagnosis|6852,6859|false|false|false|C0012634|Disease|Disease
Event|Event|Principle Diagnosis|6852,6859|false|false|false|||Disease
Finding|Mental Process|Discharge Condition|6884,6890|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|6884,6897|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|6884,6897|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|6891,6897|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|6891,6897|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|6899,6904|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|6899,6904|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|6909,6917|false|false|false|||coherent
Finding|Finding|Discharge Condition|6909,6917|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|6919,6924|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|6919,6941|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|6919,6941|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|6928,6941|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|6928,6941|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|6928,6941|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|6943,6948|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|6943,6948|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|6943,6948|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|6943,6948|false|false|false|||Alert
Finding|Finding|Discharge Condition|6943,6948|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|6943,6948|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|6943,6948|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|6953,6964|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|6953,6964|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|6966,6974|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|6966,6974|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|6966,6974|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|6975,6981|false|false|false|C5889824||Status
Event|Event|Discharge Condition|6975,6981|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|6975,6981|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|6983,6993|false|false|false|||Ambulatory
Finding|Functional Concept|Discharge Condition|6983,6993|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|6983,6993|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|6983,6993|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|6983,6993|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|6996,7007|false|false|false|||Independent
Finding|Finding|Discharge Condition|6996,7007|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Condition|6996,7007|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Event|Event|Discharge Instructions|7045,7053|false|false|false|||admitted
Finding|Idea or Concept|Discharge Instructions|7061,7069|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|Discharge Instructions|7078,7083|false|false|false|||fever
Finding|Finding|Discharge Instructions|7078,7083|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|Discharge Instructions|7078,7083|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Procedure|Diagnostic Procedure|Discharge Instructions|7103,7110|false|false|false|C0040405|X-Ray Computed Tomography|CT scan
Event|Event|Discharge Instructions|7106,7110|false|false|false|||scan
Procedure|Diagnostic Procedure|Discharge Instructions|7106,7110|false|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Anatomy|Body Location or Region|Discharge Instructions|7119,7124|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Discharge Instructions|7119,7124|false|false|false|C0741025|Chest problem|chest
Event|Event|Discharge Instructions|7130,7136|false|false|false|||showed
Finding|Finding|Discharge Instructions|7146,7152|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Discharge Instructions|7146,7152|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Disorder|Disease or Syndrome|Discharge Instructions|7159,7168|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|Discharge Instructions|7159,7168|false|false|false|||pneumonia
Finding|Functional Concept|Discharge Instructions|7177,7182|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|7177,7187|false|false|false|C0225706|Right lung|right lung
Anatomy|Body Location or Region|Discharge Instructions|7183,7187|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|7183,7187|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Discharge Instructions|7183,7187|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Discharge Instructions|7183,7187|false|false|false|C0740941|Lung Problem|lung
Event|Event|Discharge Instructions|7199,7206|false|false|false|||started
Drug|Antibiotic|Discharge Instructions|7210,7221|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|Discharge Instructions|7210,7221|false|false|false|||antibiotics
Event|Event|Discharge Instructions|7226,7231|false|false|false|||treat
Disorder|Disease or Syndrome|Discharge Instructions|7237,7246|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|Discharge Instructions|7237,7246|false|false|false|||pneumonia
Drug|Biologically Active Substance|Discharge Instructions|7275,7281|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|Discharge Instructions|7275,7281|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|Discharge Instructions|7275,7281|false|false|false|C0030054|oxygen|oxygen
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|7275,7281|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Event|Event|Discharge Instructions|7282,7293|false|false|false|||requirement
Finding|Functional Concept|Discharge Instructions|7282,7293|false|false|false|C1514873|Requirement|requirement
Event|Event|Discharge Instructions|7305,7311|false|false|false|||ALWAYS
Finding|Finding|Discharge Instructions|7305,7311|false|false|false|C1549493;C3812891|All of the Time;Always - AcknowledgementCondition|ALWAYS
Finding|Idea or Concept|Discharge Instructions|7305,7311|false|false|false|C1549493;C3812891|All of the Time;Always - AcknowledgementCondition|ALWAYS
Event|Event|Discharge Instructions|7313,7317|false|false|false|||wear
Finding|Functional Concept|Discharge Instructions|7318,7330|false|false|false|C2348609|Supplement|supplemental
Finding|Finding|Discharge Instructions|7318,7337|false|false|false|C4534306|Supplemental oxygen|supplemental oxygen
Drug|Biologically Active Substance|Discharge Instructions|7331,7337|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|Discharge Instructions|7331,7337|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|Discharge Instructions|7331,7337|false|false|false|C0030054|oxygen|oxygen
Event|Event|Discharge Instructions|7331,7337|false|false|false|||oxygen
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|7331,7337|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Event|Activity|Discharge Instructions|7341,7345|false|false|false|C0871208|Rating (action)|rate
Event|Event|Discharge Instructions|7341,7345|false|false|false|||rate
Finding|Idea or Concept|Discharge Instructions|7341,7345|false|false|false|C1549480|Amount type - Rate|rate
Finding|Finding|Discharge Instructions|7386,7389|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Discharge Instructions|7386,7389|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Finding|Discharge Instructions|7386,7401|false|false|false|C0850869|blood count low|low blood count
Disorder|Disease or Syndrome|Discharge Instructions|7390,7395|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Discharge Instructions|7390,7395|false|false|false|||blood
Finding|Body Substance|Discharge Instructions|7390,7395|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Procedure|Laboratory Procedure|Discharge Instructions|7390,7401|false|false|false|C0005771|Blood Cell Count|blood count
Event|Event|Discharge Instructions|7396,7401|false|false|false|||count
Disorder|Disease or Syndrome|Discharge Instructions|7419,7424|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Discharge Instructions|7419,7424|false|false|false|||blood
Finding|Body Substance|Discharge Instructions|7419,7424|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Event|Discharge Instructions|7426,7437|false|false|false|||transfusion
Finding|Functional Concept|Discharge Instructions|7426,7437|false|false|false|C0199960||transfusion
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|7426,7437|false|false|false|C0005841;C1879316|Blood Transfusion;Transfusion (procedure)|transfusion
Event|Event|Discharge Instructions|7447,7451|false|false|false|||felt
Disorder|Disease or Syndrome|Discharge Instructions|7462,7467|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Discharge Instructions|7462,7467|false|false|false|||blood
Finding|Body Substance|Discharge Instructions|7462,7467|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Procedure|Laboratory Procedure|Discharge Instructions|7462,7473|false|false|false|C0005771|Blood Cell Count|blood count
Event|Event|Discharge Instructions|7468,7473|false|false|false|||count
Event|Event|Discharge Instructions|7478,7481|false|false|false|||low
Finding|Finding|Discharge Instructions|7478,7481|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Discharge Instructions|7478,7481|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Event|Event|Discharge Instructions|7490,7502|false|false|false|||chemotherapy
Finding|Functional Concept|Discharge Instructions|7490,7502|false|false|false|C0013217|pharmacotherapeutic|chemotherapy
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|7490,7502|false|false|false|C0013216;C0392920;C3665472|Chemotherapy;Chemotherapy Regimen;Pharmacotherapy|chemotherapy
Event|Event|Discharge Instructions|7516,7521|false|false|false|||weigh
Event|Event|Discharge Instructions|7549,7553|false|false|false|||call
Finding|Intellectual Product|Discharge Instructions|7559,7565|false|false|false|C2348314|Doctor - Title|doctor
Event|Event|Discharge Instructions|7601,7607|false|false|false|||notice
Event|Event|Discharge Instructions|7619,7628|false|false|false|||shortness
Finding|Body Substance|Discharge Instructions|7633,7639|false|false|false|C0225386|Breath|breath
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|7644,7647|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Pathologic Function|Discharge Instructions|7644,7656|false|true|false|C0581394|Swelling of lower limb|leg swelling
Event|Event|Discharge Instructions|7648,7656|false|false|false|||swelling
Finding|Finding|Discharge Instructions|7648,7656|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|Discharge Instructions|7648,7656|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Event|Event|Discharge Instructions|7659,7666|false|false|false|||Changes
Finding|Functional Concept|Discharge Instructions|7659,7666|false|false|false|C0392747|Changing|Changes
Attribute|Clinical Attribute|Discharge Instructions|7675,7686|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|7675,7686|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|7675,7686|false|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|7675,7686|false|false|false|C4284232|Medications|medications
Event|Event|Discharge Instructions|7688,7693|false|false|false|||ADDED
Finding|Idea or Concept|Discharge Instructions|7694,7704|false|false|false|C0549178|Continuous|continuous
Event|Event|Discharge Instructions|7705,7717|false|false|false|||supplemental
Finding|Functional Concept|Discharge Instructions|7705,7717|false|false|false|C2348609|Supplement|supplemental
Finding|Finding|Discharge Instructions|7705,7724|false|false|false|C4534306|Supplemental oxygen|supplemental oxygen
Drug|Biologically Active Substance|Discharge Instructions|7718,7724|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|Discharge Instructions|7718,7724|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|Discharge Instructions|7718,7724|false|false|false|C0030054|oxygen|oxygen
Event|Event|Discharge Instructions|7718,7724|false|false|false|||oxygen
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|7718,7724|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Event|Event|Discharge Instructions|7748,7753|false|false|false|||ADDED
Drug|Antibiotic|Discharge Instructions|7754,7764|false|false|false|C0007562|cefuroxime|cefuroxime
Drug|Organic Chemical|Discharge Instructions|7754,7764|false|false|false|C0007562|cefuroxime|cefuroxime
Event|Event|Discharge Instructions|7754,7764|false|false|false|||cefuroxime
Disorder|Mental or Behavioral Dysfunction|Discharge Instructions|7772,7775|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Discharge Instructions|7772,7775|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Discharge Instructions|7772,7775|false|false|false|C1530795|BID protein, human|BID
Event|Event|Discharge Instructions|7772,7775|false|false|false|||BID
Finding|Gene or Genome|Discharge Instructions|7772,7775|false|false|false|C1332410|BID gene|BID
Drug|Antibiotic|Discharge Instructions|7798,7810|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|Discharge Instructions|7798,7810|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|Discharge Instructions|7798,7810|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Event|Event|Discharge Instructions|7798,7810|false|false|false|||azithromycin
Finding|Functional Concept|Discharge Instructions|7817,7825|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Discharge Instructions|7820,7825|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Discharge Instructions|7820,7825|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Event|Discharge Instructions|7842,7847|false|false|false|||ADDED
Drug|Organic Chemical|Discharge Instructions|7848,7853|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|Discharge Instructions|7848,7853|false|false|false|C3489575|sennosides, USP|Senna
Drug|Biomedical or Dental Material|Discharge Instructions|7856,7859|false|false|false|C0039225|Tablet Dosage Form|tab
Event|Event|Discharge Instructions|7856,7859|false|false|false|||tab
Event|Event|Discharge Instructions|7875,7881|false|false|false|||needed
Event|Event|Discharge Instructions|7886,7898|false|false|false|||constipation
Finding|Sign or Symptom|Discharge Instructions|7886,7898|false|false|false|C0009806|Constipation|constipation
Event|Event|Discharge Instructions|7899,7904|false|false|false|||ADDED
Drug|Biomedical or Dental Material|Discharge Instructions|7905,7917|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Drug|Organic Chemical|Discharge Instructions|7905,7917|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Drug|Organic Chemical|Discharge Instructions|7905,7924|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Pharmacologic Substance|Discharge Instructions|7905,7924|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Hazardous or Poisonous Substance|Discharge Instructions|7918,7924|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Drug|Organic Chemical|Discharge Instructions|7918,7924|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Event|Event|Discharge Instructions|7918,7924|false|false|false|||Glycol
Drug|Organic Chemical|Discharge Instructions|7926,7933|false|false|false|C0876088|Miralax|Miralax
Drug|Pharmacologic Substance|Discharge Instructions|7926,7933|false|false|false|C0876088|Miralax|Miralax
Event|Event|Discharge Instructions|7937,7943|false|false|false|||packet
Event|Event|Discharge Instructions|7953,7959|false|false|false|||needed
Event|Event|Discharge Instructions|7965,7977|false|false|false|||constipation
Finding|Sign or Symptom|Discharge Instructions|7965,7977|false|false|false|C0009806|Constipation|constipation
Procedure|Health Care Activity|Discharge Instructions|7980,7988|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|7989,8001|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|7989,8001|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|7989,8001|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

