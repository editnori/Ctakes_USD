CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|Known|Modifier|false|false||Knownnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Adverse reaction to drug|Finding|true|false||Adverse Drug Reactionsnull|Adverse reaction to drug|Finding|true|false||Drug Reactionsnull|Pharmaceutical Preparations|Drug|false|false||Drug
null|Pharmacologic Substance|Drug|false|false||Drugnull|Drug problem|Finding|false|false||Drugnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Structure of right flank|Anatomy|false|false|C1552823;C2598155;C0009938;C2136686;C1549543;C0030193;C0085639|Right flanknull|Table Cell Horizontal Align - right|Finding|false|false|C0230171;C0733995|Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Flank (surface region)|Anatomy|false|false|C1549543;C0030193;C1552823;C2136686;C0009938|flanknull|Contusions|Disorder|false|false|C0733995;C0230171|bruisingnull|reported bruising (history)|Finding|false|false|C0230171;C0733995|bruisingnull|Administration Method - Pain|Finding|false|false|C0230171;C0733995|pain
null|Pain|Finding|false|false|C0230171;C0733995|painnull|null|Attribute|false|false|C0733995|painnull|Falls|Finding|false|false|C0733995|fallnull|Autumn|Time|false|false||fallnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Mathematical Factor|Finding|false|false||factor
null|Factor|Finding|false|false||factor
null|Feelings about Genomic Testing Results|Finding|false|false||factornull|Malnutrition|Disorder|false|false||deficiencynull|Deficiency|Finding|false|false||deficiencynull|deficiency aspects|Modifier|false|false||deficiencynull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Neck swelling|Finding|false|false|C0027530;C3159206|neck swellingnull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|neck
null|Neck problem|Finding|false|false|C0027530;C3159206|necknull|dendritic spine neck|Anatomy|false|false|C2046386;C1546397;C0812434;C0684335;C0578454|neck
null|Neck|Anatomy|false|false|C2046386;C1546397;C0812434;C0684335;C0578454|necknull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Snowboarding (activity)|Finding|false|false||snowboarding
null|snowboarding (history)|Finding|false|false||snowboardingnull|Admission Type - Accident|Finding|false|false|C0027530;C3159206|accident
null|history of accident|Finding|false|false|C0027530;C3159206|accidentnull|Accidents|Phenomenon|false|false||accidentnull|Accidental event (event)|Event|false|false||accidentnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Loss (adaptation)|Finding|false|false||lossnull|Loss (quantitative)|LabModifier|false|false||lossnull|Consciousness related finding|Finding|false|false||consciousness
null|Conscious|Finding|false|false||consciousness
null|null|Finding|false|false||consciousnessnull|Initially|Time|false|false||initiallynull|Imaging of head|Procedure|false|false|C0018670;C0152336|imaging of headnull|Imaging problem|Finding|false|false|C0018670;C0152336|imagingnull|Diagnostic Imaging|Procedure|false|false|C0018670;C0152336|imaging
null|Imaging Techniques|Procedure|false|false|C0018670;C0152336|imagingnull|Imaging Technology|Title|false|false||imagingnull|Problems with head|Disorder|false|false|C0027530;C3159206;C0018670;C0152336|headnull|Procedure on head|Procedure|false|false|C0018670;C0152336;C0027530;C3159206|headnull|Structure of head of caudate nucleus|Anatomy|false|false|C2711858;C0812434;C0684335;C0079595;C0011923;C0876917;C0362076;C0740845|head
null|Head|Anatomy|false|false|C2711858;C0812434;C0684335;C0079595;C0011923;C0876917;C0362076;C0740845|headnull|Head Device|Device|false|false||headnull|Passive joint movement of neck (finding)|Finding|false|false|C0018670;C0152336;C0027530;C3159206|neck
null|Neck problem|Finding|false|false|C0018670;C0152336;C0027530;C3159206|necknull|dendritic spine neck|Anatomy|false|false|C0362076;C0812434;C0684335;C0876917|neck
null|Neck|Anatomy|false|false|C0362076;C0812434;C0684335;C0876917|necknull|Intracranial Hemorrhage|Finding|false|false|C0524466|intracranial hemorrhagenull|Intracranial Route of Administration|Finding|false|false|C0524466|intracranialnull|Intracranial|Anatomy|false|false|C0019080;C0151699;C1522213|intracranialnull|Hemorrhage|Finding|false|false|C0524466|hemorrhagenull|Cancer/Testis Antigen|Drug|false|false|C0027530;C3159206|CTAnull|PCYT1A wt Allele|Finding|false|false|C0027530;C3159206|CTA
null|CERNA3 gene|Finding|false|false|C0027530;C3159206|CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false|C0027530;C3159206|CTAnull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|neck
null|Neck problem|Finding|false|false|C0027530;C3159206|necknull|dendritic spine neck|Anatomy|false|false|C3813556;C1552823;C3272310;C0812434;C0684335;C3540513;C4554671|neck
null|Neck|Anatomy|false|false|C3813556;C1552823;C3272310;C0812434;C0684335;C3540513;C4554671|necknull|Table Cell Horizontal Align - right|Finding|false|false|C0027530;C3159206|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Structure of platysma muscle|Anatomy|false|false|C1285542;C0018944|platysma musclenull|Structure of platysma muscle|Anatomy|false|false||platysmanull|Pterostichus (Platysma)|Entity|false|false||platysmanull|Muscle (organ)|Anatomy|false|false|C0018944;C1285542|muscle
null|Muscle Tissue|Anatomy|false|false|C0018944;C1285542|musclenull|Hematoma|Finding|false|false|C4083049;C0026845;C0224176|hematomanull|Has focus|Finding|false|false|C0224176;C4083049;C0026845|focusnull|Focal|Modifier|false|false||focusnull|Contrast Media|Drug|false|false|C0224176;C0921006|contrastnull|Contrast|Modifier|false|false||contrastnull|Extravasation of Diagnostic and Therapeutic Materials|Disorder|false|false|C0921006;C0224176;C4083049;C0026845;C0921006;C0224176|extravasationnull|Extravasation|Finding|false|false|C0921006;C4083049;C0026845;C0224176;C0921006|extravasationnull|Right platysma|Anatomy|false|false|C0015376;C0009924;C0015379;C1552823|right platysma musclenull|Right platysma|Anatomy|false|false|C1552823;C0015379;C0015376|right platysmanull|Table Cell Horizontal Align - right|Finding|false|false|C0921006;C4083049;C0026845;C0921006;C0224176|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Structure of platysma muscle|Anatomy|false|false|C0009924;C0015379;C0015376;C1552823|platysma musclenull|Structure of platysma muscle|Anatomy|false|false|C0015379|platysmanull|Pterostichus (Platysma)|Entity|false|false||platysmanull|Muscle (organ)|Anatomy|false|false|C0015376;C0015379;C1552823|muscle
null|Muscle Tissue|Anatomy|false|false|C0015376;C0015379;C1552823|musclenull|Structure of right shoulder region|Anatomy|false|false|C0869975;C0221590;C0018944;C1552823|right shouldernull|Table Cell Horizontal Align - right|Finding|false|false|C0524468|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Examination of shoulder(s)|Procedure|false|false|C0524468;C0037004;C4299050|shoulder
null|Procedures on Shoulder|Procedure|false|false|C0524468;C0037004;C4299050|shouldernull|Upper extremity>Shoulder|Anatomy|false|false|C0869975;C0221590|shoulder
null|Shoulder|Anatomy|false|false|C0869975;C0221590|shouldernull|Hematoma|Finding|false|false|C0524468|hematomanull|Examination of shoulder(s)|Procedure|false|false|C0037004;C4299050|shoulder
null|Procedures on Shoulder|Procedure|false|false|C0037004;C4299050|shouldernull|Upper extremity>Shoulder|Anatomy|false|false|C0869975;C0221590|shoulder
null|Shoulder|Anatomy|false|false|C0869975;C0221590|shouldernull|null|Finding|false|false||filmsnull|film (photographic)|Device|false|false||filmsnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Congenital Abnormality|Disorder|false|false||abnormalitynull|Abnormality|Finding|false|false||abnormalitynull|Diagnostic Service Section ID - Hematology|Finding|false|false||Hematologynull|diagnostic service sources hematology (procedure)|Procedure|false|false||Hematology
null|Hematology procedure|Procedure|false|false||Hematology
null|Hematologic Tests|Procedure|false|false||Hematologynull|hematology (field)|Title|false|false||Hematologynull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|DDAVP|Drug|false|false||DDAVP
null|DDAVP|Drug|false|false||DDAVP
null|DDAVP|Drug|false|false||DDAVPnull|Mathematical Factor|Finding|false|false||factor
null|Factor|Finding|false|false||factor
null|Feelings about Genomic Testing Results|Finding|false|false||factornull|Biological Assay|Procedure|false|false||assay
null|Assay|Procedure|false|false||assaynull|assay qualifier|Modifier|false|false||assaynull|Report (document)|Finding|false|false||reportnull|Reporting|Procedure|false|false||reportnull|null|Attribute|false|false||reportnull|Report (document)|Finding|false|false||reportnull|Reporting|Procedure|false|false||reportnull|null|Attribute|false|false||reportnull|Hemoglobin below reference range|Finding|false|false||hemoglobin decreasednull|Hemoglobin|Drug|false|false||hemoglobin
null|chrysarobin|Drug|false|false||hemoglobin
null|chrysarobin|Drug|false|false||hemoglobin
null|Hemoglobin|Drug|false|false||hemoglobinnull|Hemoglobin finding|Finding|false|false||hemoglobinnull|Hemoglobin measurement|Procedure|false|false||hemoglobinnull|Repeat Object|Finding|false|false||Repeat
null|Repeat|Finding|false|false||Repeatnull|Repeat Pattern|Time|false|false||Repeatnull|Imaging problem|Finding|false|false||imagingnull|Diagnostic Imaging|Procedure|false|false||imaging
null|Imaging Techniques|Procedure|false|false||imagingnull|Imaging Technology|Title|false|false||imagingnull|Morning|Time|false|false||in the morningnull|Morning|Time|false|false||morningnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Female genital injuries|Disorder|false|false||injuries
null|Male Genital Injuries|Disorder|false|false||injuries
null|Traumatic injury|Disorder|false|false||injuries
null|urologic injuries|Disorder|false|false||injuriesnull|trauma qualifier|Modifier|false|false||injuriesnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Hematologist|Subject|false|false||hematologistnull|Hemoglobin|Drug|false|false||hemoglobin
null|chrysarobin|Drug|false|false||hemoglobin
null|chrysarobin|Drug|false|false||hemoglobin
null|Hemoglobin|Drug|false|false||hemoglobinnull|Hemoglobin finding|Finding|false|false||hemoglobinnull|Hemoglobin measurement|Procedure|false|false||hemoglobinnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Reduced|Finding|false|false||decreasenull|Decrease|LabModifier|false|false||decreasenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Hemoglobin|Drug|false|false||hemoglobin
null|chrysarobin|Drug|false|false||hemoglobin
null|chrysarobin|Drug|false|false||hemoglobin
null|Hemoglobin|Drug|false|false||hemoglobinnull|Hemoglobin finding|Finding|false|false||hemoglobinnull|Hemoglobin measurement|Procedure|false|false||hemoglobinnull|Flank (surface region)|Anatomy|false|false||flanknull|Hematoma|Finding|false|false||hematomanull|Concern|Finding|false|false|C0035359|concernnull|Retroperitoneal Space|Anatomy|false|false|C2699424|retroperitonealnull|Hemorrhage|Finding|false|false||bleednull|Has patient|Finding|false|false||patient hasnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|DDAVP|Drug|false|false||DDAVP
null|DDAVP|Drug|false|false||DDAVP
null|DDAVP|Drug|false|false||DDAVPnull|Admission Type - Accident|Finding|false|false||accident
null|history of accident|Finding|false|false||accidentnull|Accidents|Phenomenon|false|false||accidentnull|Accidental event (event)|Event|false|false||accidentnull|Lightheadedness|Finding|true|false||lightheadednessnull|Palpitations|Finding|false|false||palpitationsnull|Increase|Finding|true|false||increasenull|Neck swelling|Finding|false|false|C0027530;C3159206|neck swellingnull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|neck
null|Neck problem|Finding|false|false|C0027530;C3159206|necknull|dendritic spine neck|Anatomy|false|false|C0812434;C0684335;C0578454|neck
null|Neck|Anatomy|false|false|C0812434;C0684335;C0578454|necknull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Course|Time|false|false||coursenull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Administration Method - Pain|Finding|false|false|C0524468;C0037004;C4299050|pain
null|Pain|Finding|false|false|C0524468;C0037004;C4299050|painnull|null|Attribute|false|false||painnull|Structure of right shoulder region|Anatomy|false|false|C0869975;C0221590;C1552823;C1549543;C0030193|right shouldernull|Table Cell Horizontal Align - right|Finding|false|false|C0524468;C0037004;C4299050|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Examination of shoulder(s)|Procedure|false|false|C0524468;C0037004;C4299050|shoulder
null|Procedures on Shoulder|Procedure|false|false|C0524468;C0037004;C4299050|shouldernull|Upper extremity>Shoulder|Anatomy|false|false|C0869975;C0221590;C1552823;C1549543;C0030193|shoulder
null|Shoulder|Anatomy|false|false|C0869975;C0221590;C1552823;C1549543;C0030193|shouldernull|Course|Time|false|false||coursenull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Initial (abbreviation)|Finding|false|false||initialnull|Initially|Time|false|false||initialnull|Firstly|Modifier|false|false||initialnull|Taking vital signs|Procedure|false|false||vital signsnull|null|Attribute|false|false||vital signs
null|Vital signs|Attribute|false|false||vital signsnull|Vital High Nitrogen Enteral Nutrition|Drug|false|false||vitalnull|Vital (qualifier value)|Modifier|false|false||vitalnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Initial (abbreviation)|Finding|false|false||Initialnull|Initially|Time|false|false||Initialnull|Firstly|Modifier|false|false||Initialnull|Laboratory test finding|Lab|false|false||labsnull|Hemoglobin|Drug|false|false||hemoglobin
null|chrysarobin|Drug|false|false||hemoglobin
null|chrysarobin|Drug|false|false||hemoglobin
null|Hemoglobin|Drug|false|false||hemoglobinnull|Hemoglobin finding|Finding|false|false||hemoglobinnull|Hemoglobin measurement|Procedure|false|false||hemoglobinnull|Repeat Object|Finding|false|false||repeat
null|Repeat|Finding|false|false||repeatnull|Repeat Pattern|Time|false|false||repeatnull|null|Modifier|false|false||unremarkablenull|antihemophilic factor, human recombinant|Drug|false|false||FVIII
null|antihemophilic factor, human recombinant|Drug|false|false||FVIIInull|F8 wt Allele|Finding|false|false||FVIII
null|F8 gene|Finding|false|false||FVIIInull|Activity (animal life circumstance)|Finding|false|false||activity
null|Physical activity|Finding|false|false||activitynull|Activities|Event|false|false||activitynull|null|Modifier|false|false||activitynull|Muscle (organ)|Anatomy|false|false||muscularnull|Muscular|Modifier|false|false||muscularnull|Hemorrhage|Finding|false|false||hemorrhagenull|Flank (surface region)|Anatomy|false|false||flanknull|Retroperitoneal Hemorrhage|Finding|true|false|C0035359|retroperitoneal bleednull|Retroperitoneal Space|Anatomy|false|false|C0019080;C0151705|retroperitonealnull|Hemorrhage|Finding|true|false|C0035359|bleednull|Preliminary|Time|false|false||preliminarynull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Patient Class - Outpatient|Finding|false|false||outpatient
null|Referral category - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Hematologist|Subject|false|false||hematologistnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|desmopressin|Drug|false|false||desmopressin
null|desmopressin|Drug|false|false||desmopressin
null|desmopressin|Drug|false|false||desmopressinnull|ug/g|LabModifier|false|false||mg/kgnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Disease Management|Procedure|false|false||managementnull|Management Occupations|Subject|false|false||managementnull|Management procedure|Event|false|false||management
null|Administration occupational activities|Event|false|false||managementnull|Review of|Finding|false|false||review ofnull|Review (Publication Type)|Finding|false|false||review
null|Act Class - review|Finding|false|false||reviewnull|Quantity limited request - Records|Finding|false|false||records
null|Records|Finding|false|false||recordsnull|Query Quantity Unit - Records|Modifier|false|false||recordsnull|Has patient|Finding|false|false||patient hasnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Hemorrhage|Finding|false|false||bleedingnull|Male Circumcision|Procedure|false|false||circumcisionnull|Blood Transfusion|Procedure|false|false||blood transfusionnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|null|Finding|false|false||transfusionnull|Blood Transfusion|Procedure|false|false||transfusion
null|Transfusion (procedure)|Procedure|false|false||transfusionnull|Childhood|Time|false|false||childhoodnull|Tendency to bruise easily|Finding|false|false||tendency to bruise easilynull|Easy|Finding|false|false||easilynull|Disease|Disorder|false|false||diseasenull|Late|Time|false|false||Laternull|Extraction of wisdom tooth|Procedure|false|false|C0026369;C1305762;C0040426|wisdom tooth extractionnull|Structure of wisdom tooth|Anatomy|false|false|C0185115;C0684295;C0204147;C0871611;C0040440;C1879715|wisdom tooth
null|null|Anatomy|false|false|C0185115;C0684295;C0204147;C0871611;C0040440;C1879715|wisdom toothnull|wisdom|Finding|false|false|C0040426;C0026369;C1305762|wisdomnull|Tooth Extraction|Procedure|false|false|C0026369;C1305762;C0040426|tooth extraction
null|Apical Endodontic Surgery|Procedure|false|false|C0026369;C1305762;C0040426|tooth extractionnull|Tooth structure|Anatomy|false|false|C0871611;C0040440;C1879715;C0204147|toothnull|Chemical extraction|Procedure|false|false|C0026369;C1305762|extraction
null|Extraction|Procedure|false|false|C0026369;C1305762|extractionnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Late|Time|false|false||latenull|day|Time|false|false||daysnull|Late|Time|false|false||laternull|Hemorrhage|Finding|false|false||bleedingnull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|DDAVP|Drug|false|false||DDAVP
null|DDAVP|Drug|false|false||DDAVP
null|DDAVP|Drug|false|false||DDAVPnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Hematologist|Subject|false|false||hematologistnull|Hemophilia A|Disorder|false|false||hemophilia
null|null|Disorder|false|false||hemophilianull|null|Title|false|false||hemophilianull|antihemophilic factor, human recombinant|Drug|false|false||FVIII
null|antihemophilic factor, human recombinant|Drug|false|false||FVIIInull|F8 wt Allele|Finding|false|false||FVIII
null|F8 gene|Finding|false|false||FVIIInull|Activity (animal life circumstance)|Finding|false|false||activity
null|Physical activity|Finding|false|false||activitynull|Activities|Event|false|false||activitynull|null|Modifier|false|false||activitynull|Numerous|LabModifier|false|false||multiplenull|Sometimes|Time|false|false||sometimesnull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|arrival - ActRelationshipType|Finding|false|false||arrivalnull|null|Event|false|false||arrivalnull|Floor (anatomic)|Anatomy|false|false||floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Feeling comfortable|Finding|false|false||comfortablenull|Complaint (finding)|Finding|false|false||complaintnull|null|Attribute|false|false||complaintnull|Review of systems (procedure)|Procedure|false|false||Review of Systemsnull|null|Attribute|false|false||Review of Systems
null|null|Attribute|false|false||Review of Systemsnull|Review of|Finding|false|false||Review ofnull|Review (Publication Type)|Finding|false|false||Review
null|Act Class - review|Finding|false|false||Reviewnull|System|Finding|false|false||Systemsnull|Proline dehydrogenase deficiency|Disorder|false|false||HPInull|History of present illness (finding)|Finding|false|false||HPI
null|allene oxide synthase activity|Finding|false|false||HPInull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Chills|Finding|false|false||chillsnull|Night sweats|Finding|false|false||night sweatsnull|Night time|Time|false|false||nightnull|Sweating|Finding|false|false||sweats
null|Sweat|Finding|false|false||sweatsnull|Headache|Finding|false|false||headachenull|Vision|Finding|false|false||visionnull|null|Attribute|false|false||visionnull|Specialized Stand Alone Plan - Vision|Entity|false|false||visionnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Rhinorrhea|Finding|false|false||rhinorrheanull|Congestion|Finding|false|false||congestionnull|Sore Throat brand of benzocaine & menthol|Drug|false|false|C0230069;C3665375;C0031354|sore throat
null|Sore Throat brand of Phenol|Drug|false|false|C0230069;C3665375;C0031354|sore throat
null|Sore Throat brand of Phenol|Drug|false|false|C0230069;C3665375;C0031354|sore throat
null|Sore Throat brand of benzocaine & menthol|Drug|false|false|C0230069;C3665375;C0031354|sore throatnull|Pharyngitis|Disorder|false|false|C0230069;C3665375;C0031354|sore throatnull|Sore Throat|Finding|false|false|C0230069;C3665375;C0031354|sore throatnull|Sore to touch|Finding|false|false||sore
null|Sore skin|Finding|false|false||sorenull|Sore sensation quality|Modifier|false|false||sorenull|Throat Homeopathic Medication|Drug|false|false|C0230069;C3665375;C0031354|throatnull|Specimen Type - Throat|Finding|false|false|C0230069;C3665375;C0031354|throat
null|null|Finding|false|false|C0230069;C3665375;C0031354|throatnull|Anterior portion of neck|Anatomy|false|false|C0010200;C1550663;C1547926;C1950455;C0242429;C3244654;C0723402;C0031350|throat
null|Throat|Anatomy|false|false|C0010200;C1550663;C1547926;C1950455;C0242429;C3244654;C0723402;C0031350|throat
null|Pharyngeal structure|Anatomy|false|false|C0010200;C1550663;C1547926;C1950455;C0242429;C3244654;C0723402;C0031350|throatnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false|C0230069;C3665375;C0031354|coughnull|Dyspnea|Finding|false|false||shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false||breathnull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C2926613;C1549543;C0030193;C0741025;C0008031|chest
null|Anterior thoracic region|Anatomy|false|false|C2926613;C1549543;C0030193;C0741025;C0008031|chestnull|Abdominal Pain|Finding|false|false|C0000726|pain, abdominalnull|Administration Method - Pain|Finding|false|false|C1527391;C0817096|pain
null|Pain|Finding|false|false|C1527391;C0817096|painnull|null|Attribute|false|false||painnull|Abdominal Pain|Finding|false|false|C0000726|abdominal painnull|Abdomen|Anatomy|false|false|C1549543;C0030193;C0000737;C0000737|abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Administration Method - Pain|Finding|false|false|C0000726|pain
null|Pain|Finding|false|false|C0000726|painnull|null|Attribute|false|false||painnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Vomiting|Finding|false|false||vomitingnull|rectal discharge diarrhea (physical finding)|Finding|false|false||diarrhea
null|Diarrhea|Finding|false|false||diarrheanull|Constipation|Finding|false|false||constipationnull|Hematochezia|Disorder|false|false||BRBPRnull|Melena|Finding|false|false||melenanull|Hematochezia|Disorder|false|false||hematochezianull|Blood in stool|Finding|false|false||hematochezianull|Dysuria|Finding|false|false||dysurianull|Hematuria|Disorder|false|false||hematurianull|Factor VIII Deficiency|Disorder|false|false|C2327388;C0228488|Factor VIII deficiency
null|Hemophilia A|Disorder|false|false|C2327388;C0228488|Factor VIII deficiencynull|Human Coagulation Factor VIII/Von Willebrand Factor Complex|Drug|false|false|C2327388;C0228488|Factor VIII
null|factor VIII|Drug|false|false|C2327388;C0228488|Factor VIII
null|factor VIII|Drug|false|false|C2327388;C0228488|Factor VIII
null|factor VIII|Drug|false|false|C2327388;C0228488|Factor VIII
null|factor VIII, human|Drug|false|false|C2327388;C0228488|Factor VIII
null|factor VIII, human|Drug|false|false|C2327388;C0228488|Factor VIII
null|factor VIII, human|Drug|false|false|C2327388;C0228488|Factor VIII
null|Factor viii (antihemophilic factor, human) per i.u.|Drug|false|false|C2327388;C0228488|Factor VIII
null|Human Coagulation Factor VIII/Von Willebrand Factor Complex|Drug|false|false|C2327388;C0228488|Factor VIII
null|antihemophilic factor, human recombinant|Drug|false|false|C2327388;C0228488|Factor VIII
null|antihemophilic factor, human recombinant|Drug|false|false|C2327388;C0228488|Factor VIIInull|F8 gene|Finding|false|false|C2327388;C0228488|Factor VIIInull|Mathematical Factor|Finding|false|false|C2327388;C0228488|Factor
null|Factor|Finding|false|false|C2327388;C0228488|Factor
null|Feelings about Genomic Testing Results|Finding|false|false|C2327388;C0228488|Factornull|Roman numeral VIII|Finding|false|false|C2327388;C0228488|VIII
null|COX8A gene|Finding|false|false|C2327388;C0228488|VIIInull|Lamina VIII of gray matter of spinal cord|Anatomy|false|false|C1366370;C0011155;C4520835;C2732016;C0015506;C1307126;C2732002;C5400797;C1521761;C2827422;C0445599;C1413661;C0162429;C3494187;C0019069|VIII
null|Cerebellar pyramis|Anatomy|false|false|C1366370;C0011155;C4520835;C2732016;C0015506;C1307126;C2732002;C5400797;C1521761;C2827422;C0445599;C1413661;C0162429;C3494187;C0019069|VIIInull|Malnutrition|Disorder|false|false|C2327388;C0228488|deficiencynull|Deficiency|Finding|false|false|C2327388;C0228488|deficiencynull|deficiency aspects|Modifier|false|false||deficiencynull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Relationship - Mother|Finding|false|false||mothernull|Mother (person)|Subject|false|false||mothernull|Bleeding tendency|Finding|false|false||tendency to bleednull|On admission|Time|false|false||ON ADMISSIONnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GENERALnull|General medical service|Procedure|false|false||GENERALnull|Generalized|Modifier|false|false||GENERALnull|Residential flat|Device|false|false||flatnull|Flat shape|Modifier|false|false||flatnull|BORNHOLM EYE DISEASE|Disorder|false|false||bednull|Bachelor of Education|Finding|false|false||bednull|Beds|Device|false|false||bednull|Patient Location - Bed|Modifier|false|false||bednull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|false|false||acutenull|Emotional distress|Finding|true|false||distress
null|Distress|Finding|true|false||distressnull|HEENT|Anatomy|false|false||HEENTnull|Myelofibrosis|Disorder|false|false|C0694605|MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false|C0026987|MMMnull|Remote control command - Clear|Finding|false|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|NECK
null|Neck problem|Finding|false|false|C0027530;C3159206|NECKnull|dendritic spine neck|Anatomy|false|false|C0812434;C0684335|NECK
null|Neck|Anatomy|false|false|C0812434;C0684335|NECKnull|Supple|Finding|false|false||Supplenull|Cardiac attachment|Finding|false|false|C0018787|CARDIACnull|Heart|Anatomy|false|false|C1314974|CARDIACnull|Cardiac - anatomy qualifier|Modifier|false|false||CARDIACnull|Heart murmur|Finding|true|false||murmursnull|Pericardial friction rub|Finding|true|false||rubsnull|Lung diseases|Disorder|false|false|C4037972;C0024109|LUNGnull|Lung Problem|Finding|false|false|C4037972;C0024109|LUNGnull|Chest>Lung|Anatomy|false|false|C0740941;C0024115|LUNG
null|Lung|Anatomy|false|false|C0740941;C0024115|LUNGnull|Cancer/Testis Antigen|Drug|false|false||CTAnull|PCYT1A wt Allele|Finding|false|false||CTA
null|CERNA3 gene|Finding|false|false||CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false||CTAnull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|ABDOMENnull|Abdomen problem|Finding|false|false|C0230168;C0000726|ABDOMENnull|Abdomen|Anatomy|false|false|C0153662;C0941288|ABDOMEN
null|Abdominal Cavity|Anatomy|false|false|C0153662;C0941288|ABDOMENnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|All extremities|Anatomy|false|false||EXTREMITIES
null|Limb structure|Anatomy|false|false||EXTREMITIESnull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|null|Drug|false|false||PULSESnull|Physiologic pulse|Finding|false|false||PULSESnull|Pulse taking|Procedure|false|false||PULSESnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Neurology speciality|Title|false|false||NEUROnull|Neurologic (qualifier value)|Modifier|false|false||NEUROnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765|SKIN
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765|SKINnull|Skin Specimen Source Code|Finding|false|false|C1123023;C4520765|SKIN
null|Skin Specimen|Finding|false|false|C1123023;C4520765|SKINnull|Skin, Human|Anatomy|false|false|C1546781;C0444099;C0178298;C0496955|SKIN
null|Skin|Anatomy|false|false|C1546781;C0444099;C0178298;C0496955|SKINnull|Hematoma|Finding|false|false|C0230171;C0027530;C3159206|Hematomasnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Aspect (characteristic)|Modifier|false|false||aspectnull|Aspect - Kind of quantity|LabModifier|false|false||aspectnull|Passive joint movement of neck (finding)|Finding|false|false|C0230171;C0027530;C3159206|neck
null|Neck problem|Finding|false|false|C0230171;C0027530;C3159206|necknull|dendritic spine neck|Anatomy|false|false|C0018944;C0812434;C0684335|neck
null|Neck|Anatomy|false|false|C0018944;C0812434;C0684335|necknull|Flank (surface region)|Anatomy|false|false|C0018944;C0812434;C0684335|flanknull|On discharge|Time|false|false||ON DISCHARGEnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GENERALnull|General medical service|Procedure|false|false||GENERALnull|Generalized|Modifier|false|false||GENERALnull|Residential flat|Device|false|false||flatnull|Flat shape|Modifier|false|false||flatnull|BORNHOLM EYE DISEASE|Disorder|false|false||bednull|Bachelor of Education|Finding|false|false||bednull|Beds|Device|false|false||bednull|Patient Location - Bed|Modifier|false|false||bednull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|false|false||acutenull|Emotional distress|Finding|true|false||distress
null|Distress|Finding|true|false||distressnull|HEENT|Anatomy|false|false||HEENTnull|Myelofibrosis|Disorder|false|false|C0694605|MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false|C0026987|MMMnull|Remote control command - Clear|Finding|false|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|NECK
null|Neck problem|Finding|false|false|C0027530;C3159206|NECKnull|dendritic spine neck|Anatomy|false|false|C0812434;C0684335|NECK
null|Neck|Anatomy|false|false|C0812434;C0684335|NECKnull|Supple|Finding|false|false||Supplenull|Cardiac attachment|Finding|false|false|C0018787|CARDIACnull|Heart|Anatomy|false|false|C1314974|CARDIACnull|Cardiac - anatomy qualifier|Modifier|false|false||CARDIACnull|Heart murmur|Finding|true|false||murmursnull|Pericardial friction rub|Finding|true|false||rubsnull|Lung diseases|Disorder|false|false|C4037972;C0024109|LUNGnull|Lung Problem|Finding|false|false|C4037972;C0024109|LUNGnull|Chest>Lung|Anatomy|false|false|C0740941;C0024115|LUNG
null|Lung|Anatomy|false|false|C0740941;C0024115|LUNGnull|Cancer/Testis Antigen|Drug|false|false||CTAnull|PCYT1A wt Allele|Finding|false|false||CTA
null|CERNA3 gene|Finding|false|false||CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false||CTAnull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|ABDOMENnull|Abdomen problem|Finding|false|false|C0230168;C0000726|ABDOMENnull|Abdomen|Anatomy|false|false|C0153662;C0941288|ABDOMEN
null|Abdominal Cavity|Anatomy|false|false|C0153662;C0941288|ABDOMENnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|All extremities|Anatomy|false|false||EXTREMITIES
null|Limb structure|Anatomy|false|false||EXTREMITIESnull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|null|Drug|false|false||PULSESnull|Physiologic pulse|Finding|false|false||PULSESnull|Pulse taking|Procedure|false|false||PULSESnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Neurology speciality|Title|false|false||NEUROnull|Neurologic (qualifier value)|Modifier|false|false||NEUROnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765|SKIN
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765|SKINnull|Skin Specimen Source Code|Finding|false|false|C1123023;C4520765|SKIN
null|Skin Specimen|Finding|false|false|C1123023;C4520765|SKINnull|Skin, Human|Anatomy|false|false|C0178298;C0496955;C1546781;C0444099|SKIN
null|Skin|Anatomy|false|false|C0178298;C0496955;C1546781;C0444099|SKINnull|Hematoma|Finding|false|false|C0027530;C3159206;C0230171|Hematomasnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Aspect (characteristic)|Modifier|false|false||aspectnull|Aspect - Kind of quantity|LabModifier|false|false||aspectnull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206;C0230171|neck
null|Neck problem|Finding|false|false|C0027530;C3159206;C0230171|necknull|dendritic spine neck|Anatomy|false|false|C0812434;C0684335;C0018944|neck
null|Neck|Anatomy|false|false|C0812434;C0684335;C0018944|necknull|Flank (surface region)|Anatomy|false|false|C0812434;C0684335;C0018944|flanknull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0851353;C0005768;C0229664;C0005767|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Monos|Drug|false|false||Monos
null|Mono-S|Drug|false|false||Monos
null|Monos|Drug|false|false||Monosnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||Eos
null|Familial eosinophilia|Disorder|false|false||Eosnull|PRSS33 gene|Finding|false|false||Eos
null|IKZF4 gene|Finding|false|false||Eosnull|Eos <Loriini>|Entity|false|false||Eosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0851353;C0005768;C0229664;C0005767|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0851353;C0005768;C0229664;C0005767|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Mandibular right central incisor mesial prosthesis|Device|false|false||25PMnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0005768;C0229664;C0005767;C0851353|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Color of urine|Finding|false|false||URINE Colornull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|color additive|Drug|false|false||Color
null|Coloring Excipient|Drug|false|false||Colornull|color - solid dosage form|Modifier|false|false||Color
null|Color|Modifier|false|false||Colornull|Color quantity|LabModifier|false|false||Colornull|Yellow color|Modifier|false|false||Yellownull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Hematuria|Disorder|false|false||URINE Bloodnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Blood and lymphatic system disorders|Disorder|false|false||Bloodnull|peripheral blood|Finding|false|false||Blood
null|Blood|Finding|false|false||Blood
null|In Blood|Finding|false|false||Bloodnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|nitrite ion|Drug|false|false||Nitrite
null|Nitrites|Drug|false|false||Nitrite
null|Nitrites|Drug|false|false||Nitrite
null|Nitrites|Drug|false|false||Nitrite
null|nitrite ion|Drug|false|false||Nitrite
null|nitrite ion|Drug|false|false||Nitritenull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Proteins|Drug|false|false||Protein
null|Proteins|Drug|false|false||Proteinnull|Protein Info|Finding|false|false||Proteinnull|Protein measurement|Procedure|false|false||Proteinnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Ketones|Drug|false|false||Ketonenull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|null|Lab|false|false|C0014792|URINE RBC
null|Red blood cells urine positive|Lab|false|false|C0014792|URINE RBCnull|Portion of urine|Finding|false|false|C0014792|URINE
null|null|Finding|false|false|C0014792|URINE
null|Urine|Finding|false|false|C0014792|URINE
null|In Urine|Finding|false|false|C0014792|URINE
null|Urine specimen|Finding|false|false|C0014792|URINEnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C0221752;C2188659;C0042036;C2963137;C0042037;C1547942;C1610733;C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Leukocytes|Anatomy|false|false||WBCnull|Yeast, Dried|Drug|false|false||Yeast
null|Candida albicans allergenic extract|Drug|false|false||Yeast
null|Candida albicans allergenic extract|Drug|false|false||Yeast
null|Candida albicans allergenic extract|Drug|false|false||Yeastnull|Saccharomyces cerevisiae|Entity|false|false||Yeast
null|Yeasts|Entity|false|false||Yeastnull|Tissue Factor Pathway Inhibitor, human|Drug|false|false||Epi
null|epinephrine|Drug|false|false||Epi
null|epinephrine|Drug|false|false||Epi
null|epinephrine|Drug|false|false||Epi
null|Tissue Factor Pathway Inhibitor, human|Drug|false|false||Epinull|Exocrine pancreatic insufficiency|Disorder|false|false||Epinull|Eysenck personality inventory|Finding|false|false||Epi
null|TFPI wt Allele|Finding|false|false||Epi
null|TFPI gene|Finding|false|false||Epinull|Electronic Portal Imaging|Procedure|false|false||Epi
null|Echo-Planar Imaging|Procedure|false|false||Epinull|Mucus in urine (finding)|Finding|false|false||URINE Mucousnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Mucus (substance)|Finding|false|false||Mucous
null|mucus layer|Finding|false|false||Mucousnull|Mucous appearance|Modifier|false|false||Mucousnull|Retinoic Acid Response Element|Finding|false|false||RAREnull|Infrequent|Time|false|false||RAREnull|Rare|Modifier|false|false||RAREnull|Imaging problem|Finding|false|false||IMAGINGnull|Diagnostic Imaging|Procedure|false|false||IMAGING
null|Imaging Techniques|Procedure|false|false||IMAGINGnull|Imaging Technology|Title|false|false||IMAGINGnull|Scientific Study|Procedure|false|false||STUDIESnull|Choline-Phosphate Cytidylyltransferase A|Drug|false|false||CT A
null|Choline-Phosphate Cytidylyltransferase A|Drug|false|false||CT Anull|Acute hemorrhage|Finding|false|false|C0446499;C0230171|Acute hemorrhagenull|Admission Level of Care Code - Acute|Finding|false|false||Acute
null|Acute - Triage Code|Finding|false|false||Acutenull|acute|Time|false|false||Acutenull|Hemorrhage|Finding|false|false||hemorrhagenull|Right posterior|Modifier|false|false||right posteriornull|Table Cell Horizontal Align - right|Finding|false|false|C0446499|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Posterior abdominal surface region|Anatomy|false|false|C0751438;C0333276;C1552823|posterior flanknull|Posterior pituitary disease|Disorder|false|false|C0446499;C0230171|posteriornull|Dorsal|Modifier|false|false||posteriornull|Flank (surface region)|Anatomy|false|false|C0333276;C0751438|flanknull|Set of muscles|Anatomy|false|false||musculaturenull|Probably|Finding|false|false|C0934502|probably
null|Probable diagnosis|Finding|false|false|C0934502|probablynull|anatomical layer|Anatomy|false|false|C0332148;C0750492|layeringnull|Hardness|Modifier|false|false||hardnull|Set of muscles|Anatomy|false|false|C0019080|musculaturenull|Hemorrhage|Finding|false|false|C1995013|hemorrhagenull|Extravasation of Diagnostic and Therapeutic Materials|Disorder|true|false||extravasationnull|Extravasation|Finding|true|false||extravasationnull|Probable diagnosis|Finding|false|false|C0733996|Probablenull|Probability|LabModifier|false|false||Probablenull|Old|Time|false|false||oldnull|Hematoma|Finding|false|false|C0733996;C0230171|hematomanull|Posterior pituitary disease|Disorder|false|false|C0733996;C0230171|posteriornull|Dorsal|Modifier|false|false||posteriornull|Structure of left flank|Anatomy|false|false|C0332148;C1552822;C0751438;C0018944|left flanknull|Table Cell Horizontal Align - left|Finding|false|false|C0733996;C0230171|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Flank (surface region)|Anatomy|false|false|C0751438;C1552822;C0018944|flanknull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|antihemophilic factor, human recombinant|Drug|false|false||FVIII
null|antihemophilic factor, human recombinant|Drug|false|false||FVIIInull|F8 wt Allele|Finding|false|false||FVIII
null|F8 gene|Finding|false|false||FVIIInull|Malnutrition|Disorder|false|false||deficiencynull|Deficiency|Finding|false|false||deficiencynull|deficiency aspects|Modifier|false|false||deficiencynull|Snowboarding (activity)|Finding|false|false||snowboarding
null|snowboarding (history)|Finding|false|false||snowboardingnull|Admission Type - Accident|Finding|false|false||accident
null|history of accident|Finding|false|false||accidentnull|Accidents|Phenomenon|false|false||accidentnull|Accidental event (event)|Event|false|false||accidentnull|Numerous|LabModifier|false|false||multiplenull|Hematoma|Finding|false|false||hematomasnull|Hemoglobin|Drug|false|false||hemoglobin
null|chrysarobin|Drug|false|false||hemoglobin
null|chrysarobin|Drug|false|false||hemoglobin
null|Hemoglobin|Drug|false|false||hemoglobinnull|Hemoglobin finding|Finding|false|false||hemoglobinnull|Hemoglobin measurement|Procedure|false|false||hemoglobinnull|Continuous|Finding|false|false||ongoingnull|Hemorrhage|Finding|false|false||bleedingnull|Factor VIII Deficiency|Disorder|false|false|C2327388;C0228488|FACTOR VIII DEFICIENCY
null|Hemophilia A|Disorder|false|false|C2327388;C0228488|FACTOR VIII DEFICIENCYnull|Human Coagulation Factor VIII/Von Willebrand Factor Complex|Drug|false|false|C2327388;C0228488|FACTOR VIII
null|factor VIII|Drug|false|false|C2327388;C0228488|FACTOR VIII
null|factor VIII|Drug|false|false|C2327388;C0228488|FACTOR VIII
null|factor VIII|Drug|false|false|C2327388;C0228488|FACTOR VIII
null|factor VIII, human|Drug|false|false|C2327388;C0228488|FACTOR VIII
null|factor VIII, human|Drug|false|false|C2327388;C0228488|FACTOR VIII
null|factor VIII, human|Drug|false|false|C2327388;C0228488|FACTOR VIII
null|Factor viii (antihemophilic factor, human) per i.u.|Drug|false|false|C2327388;C0228488|FACTOR VIII
null|Human Coagulation Factor VIII/Von Willebrand Factor Complex|Drug|false|false|C2327388;C0228488|FACTOR VIII
null|antihemophilic factor, human recombinant|Drug|false|false|C2327388;C0228488|FACTOR VIII
null|antihemophilic factor, human recombinant|Drug|false|false|C2327388;C0228488|FACTOR VIIInull|F8 gene|Finding|false|false|C2327388;C0228488|FACTOR VIIInull|Mathematical Factor|Finding|false|false||FACTOR
null|Factor|Finding|false|false||FACTOR
null|Feelings about Genomic Testing Results|Finding|false|false||FACTORnull|Roman numeral VIII|Finding|false|false|C2327388;C0228488|VIII
null|COX8A gene|Finding|false|false|C2327388;C0228488|VIIInull|Lamina VIII of gray matter of spinal cord|Anatomy|false|false|C0162429;C3494187;C0019069;C0445599;C1413661;C4520835;C2732016;C0015506;C1307126;C2732002;C1366370;C0011155|VIII
null|Cerebellar pyramis|Anatomy|false|false|C0162429;C3494187;C0019069;C0445599;C1413661;C4520835;C2732016;C0015506;C1307126;C2732002;C1366370;C0011155|VIIInull|Malnutrition|Disorder|false|false|C2327388;C0228488|DEFICIENCYnull|Deficiency|Finding|false|false|C2327388;C0228488|DEFICIENCYnull|deficiency aspects|Modifier|false|false||DEFICIENCYnull|Numerous|LabModifier|false|false||MULTIPLEnull|Hematoma|Finding|false|false||HEMATOMASnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Presentation|Finding|false|false||presentednull|Recent|Time|false|false||recentnull|Snowboarding (activity)|Finding|false|false||snowboarding
null|snowboarding (history)|Finding|false|false||snowboardingnull|Admission Type - Accident|Finding|false|false||accident
null|history of accident|Finding|false|false||accidentnull|Accidents|Phenomenon|false|false||accidentnull|Accidental event (event)|Event|false|false||accidentnull|Imaging problem|Finding|false|false||imagingnull|Diagnostic Imaging|Procedure|false|false||imaging
null|Imaging Techniques|Procedure|false|false||imagingnull|Imaging Technology|Title|false|false||imagingnull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|neck
null|Neck problem|Finding|false|false|C0027530;C3159206|necknull|dendritic spine neck|Anatomy|false|false|C0812434;C0684335;C0018944;C0869975;C0221590|neck
null|Neck|Anatomy|false|false|C0812434;C0684335;C0018944;C0869975;C0221590|necknull|Examination of shoulder(s)|Procedure|false|false|C0037004;C4299050;C0027530;C3159206|shoulder
null|Procedures on Shoulder|Procedure|false|false|C0037004;C4299050;C0027530;C3159206|shouldernull|Upper extremity>Shoulder|Anatomy|false|false|C0869975;C0221590;C0018944|shoulder
null|Shoulder|Anatomy|false|false|C0869975;C0221590;C0018944|shouldernull|Hematoma|Finding|false|false|C0037004;C4299050;C0027530;C3159206|hematomasnull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Flank (surface region)|Anatomy|false|false|C0018944|flanknull|Hematoma|Finding|false|false|C0230171|hematomanull|Accidental Falls|Disorder|false|false||fallingnull|Falls|Finding|false|false||fallingnull|Hemoglobin|Drug|false|false||hemoglobin
null|chrysarobin|Drug|false|false||hemoglobin
null|chrysarobin|Drug|false|false||hemoglobin
null|Hemoglobin|Drug|false|false||hemoglobinnull|Hemoglobin finding|Finding|false|false||hemoglobinnull|Hemoglobin measurement|Procedure|false|false||hemoglobinnull|Concern|Finding|false|false||concernnull|Retroperitoneal Hemorrhage|Finding|false|false|C0035359|retroperitoneal bleednull|Retroperitoneal Space|Anatomy|false|false|C0019080;C0151705|retroperitonealnull|Hemorrhage|Finding|false|false|C0035359|bleednull|Hematoma|Finding|false|false||hematomanull|Flank (surface region)|Anatomy|false|false|C0015376;C0015379|flanknull|Set of muscles|Anatomy|false|false|C0015376;C0015379|musculaturenull|Extravasation of Diagnostic and Therapeutic Materials|Disorder|true|false|C1995013;C0230171|extravasationnull|Extravasation|Finding|true|false|C1995013;C0230171|extravasationnull|DDAVP|Drug|false|false||DDAVP
null|DDAVP|Drug|false|false||DDAVP
null|DDAVP|Drug|false|false||DDAVPnull|antihemophilic factor, human recombinant|Drug|false|false||FVIII
null|antihemophilic factor, human recombinant|Drug|false|false||FVIIInull|F8 wt Allele|Finding|false|false||FVIII
null|F8 gene|Finding|false|false||FVIIInull|Activity (animal life circumstance)|Finding|false|false||activity
null|Physical activity|Finding|false|false||activitynull|Activities|Event|false|false||activitynull|null|Modifier|false|false||activitynull|Complete Blood Count|Procedure|false|false|C2263086|CBCnull|Nuclear cap binding complex location|Anatomy|false|false|C0009555|CBCnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Further|Modifier|false|false||furthernull|Patient Class - Inpatient|Finding|false|false||inpatient
null|Referral category - Inpatient|Finding|false|false||inpatientnull|inpatient encounter|Procedure|false|false||inpatientnull|inpatient|Subject|false|false||inpatientnull|Preventive monitoring|Procedure|false|false||monitoringnull|null|Event|false|false||monitoringnull|Diagnostic Service Section ID - Hematology|Finding|false|false||hematologynull|diagnostic service sources hematology (procedure)|Procedure|false|false||hematology
null|Hematology procedure|Procedure|false|false||hematology
null|Hematologic Tests|Procedure|false|false||hematologynull|hematology (field)|Title|false|false||hematologynull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Hemoglobin|Drug|false|false||hemoglobin
null|chrysarobin|Drug|false|false||hemoglobin
null|chrysarobin|Drug|false|false||hemoglobin
null|Hemoglobin|Drug|false|false||hemoglobinnull|Hemoglobin finding|Finding|false|false||hemoglobinnull|Hemoglobin measurement|Procedure|false|false||hemoglobinnull|Preventive monitoring|Procedure|false|false||monitoringnull|null|Event|false|false||monitoringnull|Further|Modifier|false|false||furthernull|DDAVP|Drug|true|false||DDAVP
null|DDAVP|Drug|true|false||DDAVP
null|DDAVP|Drug|true|false||DDAVPnull|antihemophilic factor, human recombinant|Drug|false|false||FVIII
null|antihemophilic factor, human recombinant|Drug|false|false||FVIIInull|F8 wt Allele|Finding|false|false||FVIII
null|F8 gene|Finding|false|false||FVIIInull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Complete Blood Count|Procedure|false|false|C2263086|CBCnull|Nuclear cap binding complex location|Anatomy|false|false|C0009555|CBCnull|Activity (animal life circumstance)|Finding|false|false||activity
null|Physical activity|Finding|false|false||activitynull|Activities|Event|false|false||activitynull|null|Modifier|false|false||activitynull|MDF Attribute Type - Code|Finding|false|false||Code
null|A Codes|Finding|false|false||Code
null|Code|Finding|false|false||Codenull|Coding|Event|false|false||Codenull|Full|Modifier|false|false||fullnull|emergency contact|Finding|false|false||Emergency Contactnull|Consent Non-Disclosure Reason - Emergency|Finding|false|false||Emergency
null|Admission Type - Emergency|Finding|false|false||Emergency
null|Referral category - Emergency|Finding|false|false||Emergency
null|Emergencies [Disease/Finding]|Finding|false|false||Emergency
null|Consent Bypass Reason - Emergency|Finding|false|false||Emergency
null|Level of Care - Emergency|Finding|false|false||Emergency
null|Certification patient type - Emergency|Finding|false|false||Emergency
null|Encounter Admission Source - emergency|Finding|false|false||Emergency
null|Patient Class - Emergency|Finding|false|false||Emergency
null|Visit Priority Code - Emergency|Finding|false|false||Emergencynull|emergency encounter|Procedure|false|false||Emergencynull|Emergency Situation|Phenomenon|false|false||Emergencynull|Specialty Type - Emergency|Title|false|false||Emergencynull|Bale out|Time|false|false||Emergencynull|Contact - HL7 Attribution|Finding|false|false||Contact
null|Contact with|Finding|false|false||Contact
null|Communication Contact|Finding|false|false||Contactnull|contact person|Subject|false|false||Contactnull|Physical contact|Phenomenon|false|false||Contactnull|Personal Contact|Event|false|false||Contactnull|wife|Subject|false|false||wifenull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Accurate (qualifier value)|Modifier|false|false||accuratenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|null|Drug|false|false|C0028429|Desmopressin Nasalnull|desmopressin|Drug|false|false||Desmopressin
null|desmopressin|Drug|false|false||Desmopressin
null|desmopressin|Drug|false|false||Desmopressinnull|Nasal brand of oxymetazoline|Drug|false|false|C0028429|Nasal
null|Nasal brand of oxymetazoline|Drug|false|false|C0028429|Nasal
null|Nasal dosage form|Drug|false|false|C0028429|Nasalnull|Nasal Route of Administration|Finding|false|false|C0028429|Nasal
null|Nasal (intended site)|Finding|false|false|C0028429|Nasalnull|null|Anatomy|false|false|C5552704;C4520890;C1522019;C1272939;C0721966;C3212180;C0027609|Nasalnull|microgram|LabModifier|false|false||mcgnull|Tobacco containing mixture|Drug|false|false||NAS
null|N-acetylserotonin|Drug|false|false||NASnull|Neonatal Abstinence Syndrome|Disorder|false|false|C0028429|NASnull|null|Finding|false|false|C0028429|NASnull|National Academy of Sciences (U.S.)|Entity|false|false||NASnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Hemorrhage|Finding|false|false||bleedingnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every eight hours|Time|false|false||Q8Hnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|null|Drug|false|false|C0028429|Desmopressin Nasalnull|desmopressin|Drug|false|false||Desmopressin
null|desmopressin|Drug|false|false||Desmopressin
null|desmopressin|Drug|false|false||Desmopressinnull|Nasal brand of oxymetazoline|Drug|false|false|C0028429|Nasal
null|Nasal brand of oxymetazoline|Drug|false|false|C0028429|Nasal
null|Nasal dosage form|Drug|false|false|C0028429|Nasalnull|Nasal Route of Administration|Finding|false|false|C0028429|Nasal
null|Nasal (intended site)|Finding|false|false|C0028429|Nasalnull|null|Anatomy|false|false|C3212180;C4520890;C1522019;C1272939;C0721966;C5552704;C0027609|Nasalnull|microgram|LabModifier|false|false||mcgnull|Tobacco containing mixture|Drug|false|false||NAS
null|N-acetylserotonin|Drug|false|false||NASnull|Neonatal Abstinence Syndrome|Disorder|false|false|C0028429|NASnull|null|Finding|false|false|C0028429|NASnull|National Academy of Sciences (U.S.)|Entity|false|false||NASnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Hemorrhage|Finding|false|false||bleedingnull|Referral category - Outpatient|Finding|false|false||Outpatient
null|Patient Class - Outpatient|Finding|false|false||Outpatientnull|Outpatients|Subject|false|false||Outpatientnull|AML Lab Table|Finding|false|false||Lab
null|LAT2 gene|Finding|false|false||Lab
null|EWS Lab Table|Finding|false|false||Labnull|Laboratory|Device|false|false||Labnull|Labrador retriever|Entity|false|false||Lab
null|Laboratory|Entity|false|false||Labnull|Work|Event|false|false||Worknull|Complete Blood Count|Procedure|false|false|C2263086|CBCnull|Nuclear cap binding complex location|Anatomy|false|false|C0009555|CBCnull|Last|Modifier|false|false||Lastnull|Hemoglobin|Drug|false|false||hemoglobin
null|chrysarobin|Drug|false|false||hemoglobin
null|chrysarobin|Drug|false|false||hemoglobin
null|Hemoglobin|Drug|false|false||hemoglobinnull|Hemoglobin finding|Finding|false|false||hemoglobinnull|Hemoglobin measurement|Procedure|false|false||hemoglobinnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|True primary (qualifier value)|Time|false|false||PRIMARYnull|Primary|Modifier|false|false||PRIMARYnull|Admission Level of Care Code - Acute|Finding|false|false||Acute
null|Acute - Triage Code|Finding|false|false||Acutenull|acute|Time|false|false||Acutenull|Muscle (organ)|Anatomy|false|false||muscularnull|Muscular|Modifier|false|false||muscularnull|Hematoma|Finding|false|false||hematomanull|Structure of right flank|Anatomy|false|false|C1552823|right flanknull|Table Cell Horizontal Align - right|Finding|false|false|C0230171;C0733995|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Flank (surface region)|Anatomy|false|false|C1552823|flanknull|Hemophilia A|Disorder|false|false||Hemophilia
null|null|Disorder|false|false||Hemophilianull|null|Title|false|false||Hemophilianull|Mathematical Factor|Finding|false|false||factor
null|Factor|Finding|false|false||factor
null|Feelings about Genomic Testing Results|Finding|false|false||factornull|Malnutrition|Disorder|false|false||deficiencynull|Deficiency|Finding|false|false||deficiencynull|deficiency aspects|Modifier|false|false||deficiencynull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|Production Class Code - Pleasure|Finding|false|false||pleasure
null|pleasurable emotion|Finding|false|false||pleasurenull|Pleasure - Animals raised for recreation|Entity|false|false||pleasurenull|Contusions|Disorder|false|false||bruisingnull|reported bruising (history)|Finding|false|false||bruisingnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Side|Modifier|false|false||sidenull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|counts|LabModifier|false|false||countsnull|Snowboarding (activity)|Finding|false|false||snowboarding
null|snowboarding (history)|Finding|false|false||snowboardingnull|Falls|Finding|false|false||fallnull|Autumn|Time|false|false||fallnull|null|Attribute|false|false||history of hemophilianull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Hemophilia A|Disorder|false|false||hemophilia
null|null|Disorder|false|false||hemophilianull|null|Title|false|false||hemophilianull|Important|Modifier|false|false||importantnull|Code System Type - Internal|Modifier|false|false||internal
null|Internal Surface|Modifier|false|false||internal
null|Internal|Modifier|false|false||internalnull|Hemorrhage|Finding|false|false|C0230171|bleedingnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Muscle (organ)|Anatomy|false|false|C1516698;C0600644;C1704815;C1704814|muscularnull|Muscular|Modifier|false|false||muscularnull|Flank (surface region)|Anatomy|false|false|C0851353;C1516698;C0600644;C1704815;C1704814;C0019080;C0005768;C0229664;C0005767|flanknull|Blood and lymphatic system disorders|Disorder|false|false|C0230171|bloodnull|peripheral blood|Finding|false|false|C0230171|blood
null|Blood|Finding|false|false|C0230171|blood
null|In Blood|Finding|false|false|C0230171|bloodnull|Collection Object - UML Entity|Finding|false|false|C4083049;C0230171|collection
null|Item Collection|Finding|false|false|C4083049;C0230171|collection
null|Collections (publication)|Finding|false|false|C4083049;C0230171|collection
null|Collection (action)|Finding|false|false|C4083049;C0230171|collectionnull|Roman numeral VIII|Finding|false|false|C2327388;C0228488|VIII
null|COX8A gene|Finding|false|false|C2327388;C0228488|VIIInull|Lamina VIII of gray matter of spinal cord|Anatomy|false|false|C0445599;C1413661|VIII
null|Cerebellar pyramis|Anatomy|false|false|C0445599;C1413661|VIIInull|DDAVP|Drug|false|false||DDAVP
null|DDAVP|Drug|false|false||DDAVP
null|DDAVP|Drug|false|false||DDAVPnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|counts|LabModifier|false|false||countsnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Improved - answer to question|Finding|false|false||improved
null|Admission Level of Care Code - Improved|Finding|false|false||improved
null|Improved|Finding|false|false||improvednull|Better|Modifier|false|false||improvednull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Important|Modifier|false|false||importantnull|activities (history)|Finding|false|false||activitiesnull|Activities|Event|false|false||activitiesnull|Recent|Time|false|false||recentnull|Hemorrhage|Finding|false|false||bleednull|Hemophilia A|Disorder|false|false||hemophilia
null|null|Disorder|false|false||hemophilianull|null|Title|false|false||hemophilianull|Hemorrhage|Finding|false|false||Bleedingnull|Hemophiliacs|Subject|false|false||hemophiliacsnull|More|LabModifier|false|false||morenull|Potential|Modifier|false|false||potentialnull|Life|Finding|false|false||lifenull|Laser-Induced Fluorescence Endoscopy|Procedure|false|false||lifenull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|counts|LabModifier|false|false||countsnull|null|Finding|false|false|C1515974|sitenull|Anatomic Site|Anatomy|false|false|C1546778|sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Regular|Modifier|false|false||regularnull|Doctor - Title|Finding|false|false||doctornull|Physicians|Subject|false|false||doctornull|Early|Time|false|false||earlynull|next - HtmlLinkType|Finding|false|false||nextnull|Following|Time|false|false||next
null|Then|Time|false|false||nextnull|Adjacent|Modifier|false|false||nextnull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Care team|Finding|false|false||Care Teamnull|null|Attribute|false|false||Care Teamnull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|Team|Subject|false|false||Teamnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions