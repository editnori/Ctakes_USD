 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Procedure|Health Care Activity|SIMPLE_SEGMENT|46,55|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|46,60|false|false|false|C2598112||Admission Date
Finding|Body Substance|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|80,89|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|80,94|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|136,139|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|147,154|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|147,154|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Finding|Finding|SIMPLE_SEGMENT|156,163|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Finding|Functional Concept|SIMPLE_SEGMENT|156,163|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Finding|Idea or Concept|SIMPLE_SEGMENT|156,163|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|156,163|false|false|false|C0543467|Operative Surgical Procedures|SURGERY
Finding|Functional Concept|Allergies|184,193|false|false|false|C1999232|Attending (action)|Attending
Attribute|Clinical Attribute|Chief Complaint|219,225|false|false|false|C4255480||Nausea
Finding|Sign or Symptom|Chief Complaint|219,225|false|false|false|C0027497|Nausea|Nausea
Finding|Sign or Symptom|Chief Complaint|219,234|false|false|false|C0027498|Nausea and vomiting|Nausea/Vomiting
Finding|Sign or Symptom|Chief Complaint|226,234|false|false|false|C0042963|Vomiting|Vomiting
Finding|Classification|Chief Complaint|237,242|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|243,251|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|243,251|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|255,273|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|264,273|false|false|false|C0945766||Procedure
Event|Occupational Activity|Chief Complaint|264,273|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|264,273|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|264,273|false|false|false|C0184661|Interventional procedure|Procedure
Finding|Classification|Chief Complaint|280,290|false|false|false|C0376209;C0456081;C0678219;C0683269;C1546424|Adjustment - classification term;Personal Adjustment;Psychological adjustment;Transaction Type - Adjustment|adjustment
Finding|Functional Concept|Chief Complaint|280,290|false|false|false|C0376209;C0456081;C0678219;C0683269;C1546424|Adjustment - classification term;Personal Adjustment;Psychological adjustment;Transaction Type - Adjustment|adjustment
Finding|Idea or Concept|Chief Complaint|280,290|false|false|false|C0376209;C0456081;C0678219;C0683269;C1546424|Adjustment - classification term;Personal Adjustment;Psychological adjustment;Transaction Type - Adjustment|adjustment
Finding|Individual Behavior|Chief Complaint|280,290|false|false|false|C0376209;C0456081;C0678219;C0683269;C1546424|Adjustment - classification term;Personal Adjustment;Psychological adjustment;Transaction Type - Adjustment|adjustment
Disorder|Disease or Syndrome|History of Present Illness|343,346|false|false|false|C0396060|Congenital laryngeal adductor palsy|lap
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|343,346|false|false|false|C1870042|ACP2 protein, human|lap
Drug|Enzyme|History of Present Illness|343,346|false|false|false|C1870042|ACP2 protein, human|lap
Finding|Finding|History of Present Illness|343,346|false|false|false|C0456170;C1412132;C1413323;C1423544;C1424863;C1425522;C2827449;C3540509;C5575443;C5890955|ACP2 gene;ACP2 wt Allele;CEBPB gene;CEBPB wt Allele;CENPJ gene;LAP3 gene;LAP3 wt Allele;Left atrial pressure;PICALM gene;PICALM wt Allele|lap
Finding|Gene or Genome|History of Present Illness|343,346|false|false|false|C0456170;C1412132;C1413323;C1423544;C1424863;C1425522;C2827449;C3540509;C5575443;C5890955|ACP2 gene;ACP2 wt Allele;CEBPB gene;CEBPB wt Allele;CENPJ gene;LAP3 gene;LAP3 wt Allele;Left atrial pressure;PICALM gene;PICALM wt Allele|lap
Procedure|Diagnostic Procedure|History of Present Illness|343,346|false|false|false|C0031150|Laparoscopy|lap
Finding|Intellectual Product|History of Present Illness|380,384|false|false|false|C1561540|Transaction counts and value totals - week|week
Finding|Conceptual Entity|History of Present Illness|385,392|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|385,392|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|385,392|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|385,395|false|false|false|C0262926|Medical History|history of
Attribute|Clinical Attribute|History of Present Illness|396,402|false|false|false|C4255480||nausea
Finding|Sign or Symptom|History of Present Illness|396,402|false|false|false|C0027497|Nausea|nausea
Finding|Body Substance|History of Present Illness|427,433|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Physiologic Function|History of Present Illness|427,433|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Sign or Symptom|History of Present Illness|427,433|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Body Substance|History of Present Illness|437,452|false|false|false|C0558301|Undigested food|undigested food
Drug|Food|History of Present Illness|448,452|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Drug|Immunologic Factor|History of Present Illness|448,452|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Drug|Pharmacologic Substance|History of Present Illness|448,452|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Finding|Organism Function|History of Present Illness|459,465|false|false|false|C0013470|Eating|eating
Finding|Finding|History of Present Illness|467,478|false|false|false|C0231199;C1547317;C1547543;C1744706|Charge Type Reason - Intolerance;Sensitivity to Causative Agent Code - Intolerance;intolerance to substance|intolerance
Finding|Idea or Concept|History of Present Illness|467,478|false|false|false|C0231199;C1547317;C1547543;C1744706|Charge Type Reason - Intolerance;Sensitivity to Causative Agent Code - Intolerance;intolerance to substance|intolerance
Finding|Intellectual Product|History of Present Illness|467,478|false|false|false|C0231199;C1547317;C1547543;C1744706|Charge Type Reason - Intolerance;Sensitivity to Causative Agent Code - Intolerance;intolerance to substance|intolerance
Finding|Organism Function|History of Present Illness|467,478|false|false|false|C0231199;C1547317;C1547543;C1744706|Charge Type Reason - Intolerance;Sensitivity to Causative Agent Code - Intolerance;intolerance to substance|intolerance
Drug|Biomedical or Dental Material|History of Present Illness|482,488|false|false|false|C0302909;C1378566|Solid Dose Form;solid substance|solids
Drug|Substance|History of Present Illness|482,488|false|false|false|C0302909;C1378566|Solid Dose Form;solid substance|solids
Disorder|Disease or Syndrome|History of Present Illness|496,511|false|false|false|C0037036|Sialorrhea|hypersalivation
Finding|Finding|History of Present Illness|517,525|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|History of Present Illness|517,525|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Anatomy|Body Location or Region|History of Present Illness|540,550|false|false|false|C0521440|Epigastric|epigastric
Finding|Sign or Symptom|History of Present Illness|551,561|false|false|false|C2364135|Discomfort|discomfort
Finding|Finding|History of Present Illness|574,579|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|History of Present Illness|574,579|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|History of Present Illness|581,587|false|false|false|C0085593|Chills|chills
Finding|Sign or Symptom|History of Present Illness|589,600|true|false|false|C0018926|Hematemesis|hematemesis
Disorder|Disease or Syndrome|History of Present Illness|602,607|false|false|false|C0018932|Hematochezia|BRBPR
Finding|Pathologic Function|History of Present Illness|610,616|false|false|false|C0025222|Melena|melena
Finding|Finding|History of Present Illness|618,626|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|History of Present Illness|618,626|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Disorder|Disease or Syndrome|History of Present Illness|644,655|false|false|false|C0011175;C2062903|Dehydration;dehydration (Na, H2O)|dehydration
Disorder|Injury or Poisoning|History of Present Illness|644,655|false|false|false|C0011175;C2062903|Dehydration;dehydration (Na, H2O)|dehydration
Procedure|Laboratory Procedure|History of Present Illness|644,655|false|false|false|C4284399|Dehydration procedure|dehydration
Finding|Sign or Symptom|History of Present Illness|689,698|false|false|false|C0012833;C0042571|Dizziness;Vertigo|dizziness
Attribute|Clinical Attribute|History of Present Illness|715,724|false|false|false|C0945731||diagnosis
Finding|Classification|History of Present Illness|715,724|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|History of Present Illness|715,724|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|History of Present Illness|715,724|false|false|false|C0011900|Diagnosis|diagnosis
Disorder|Disease or Syndrome|History of Present Illness|734,738|false|false|false|C0155502|Benign Paroxysmal Positional Vertigo|BPPV
Finding|Body Substance|History of Present Illness|753,760|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|753,760|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|753,760|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|History of Present Illness|830,838|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|History of Present Illness|830,838|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Disorder|Disease or Syndrome|Past Medical History|971,985|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|Hyperlipidemia
Finding|Finding|Past Medical History|971,985|false|false|false|C0428465|Serum lipids high (finding)|Hyperlipidemia
Drug|Biologically Active Substance|Past Medical History|1004,1016|false|false|false|C0041004|Triglycerides|triglyceride
Drug|Organic Chemical|Past Medical History|1004,1016|false|false|false|C0041004|Triglycerides|triglyceride
Drug|Biologically Active Substance|Past Medical History|1018,1022|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|Past Medical History|1018,1022|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|Past Medical History|1018,1022|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Procedure|Laboratory Procedure|Past Medical History|1018,1022|false|false|false|C0337439|Iron measurement|iron
Disorder|Disease or Syndrome|Past Medical History|1023,1033|false|false|false|C0162429|Malnutrition|deficiency
Finding|Functional Concept|Past Medical History|1023,1033|false|false|false|C0011155|Deficiency|deficiency
Disorder|Disease or Syndrome|Past Medical History|1023,1040|false|false|false|C0041782|Deficiency anemias|deficiency anemia
Disorder|Disease or Syndrome|Past Medical History|1034,1040|false|false|false|C0002871|Anemia|anemia
Finding|Finding|Past Medical History|1042,1051|false|false|false|C0022107;C2700617|Irritability - emotion;Irritable Mood|irritable
Finding|Mental Process|Past Medical History|1042,1051|false|false|false|C0022107;C2700617|Irritability - emotion;Irritable Mood|irritable
Disorder|Disease or Syndrome|Past Medical History|1042,1057|false|false|false|C0022104|Irritable Bowel Syndrome|irritable bowel
Disorder|Disease or Syndrome|Past Medical History|1042,1066|false|false|false|C0022104|Irritable Bowel Syndrome|irritable bowel syndrome
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1052,1057|false|false|false|C0021853|Intestines|bowel
Disorder|Disease or Syndrome|Past Medical History|1058,1066|false|false|false|C0039082|Syndrome|syndrome
Finding|Functional Concept|Past Medical History|1068,1076|false|false|false|C0700624|Allergic|allergic
Disorder|Disease or Syndrome|Past Medical History|1068,1085|false|false|false|C2607914|Allergic rhinitis (disorder)|allergic rhinitis
Finding|Gene or Genome|Past Medical History|1068,1085|false|false|false|C1334103|IL13 gene|allergic rhinitis
Disorder|Disease or Syndrome|Past Medical History|1077,1085|false|false|false|C0035455|Rhinitis|rhinitis
Disorder|Disease or Syndrome|Past Medical History|1087,1099|false|false|false|C0013390|Dysmenorrhea|dysmenorrhea
Drug|Organic Chemical|Past Medical History|1101,1108|false|false|false|C0042890|Vitamins|vitamin
Drug|Pharmacologic Substance|Past Medical History|1101,1108|false|false|false|C0042890|Vitamins|vitamin
Drug|Vitamin|Past Medical History|1101,1108|false|false|false|C0042890|Vitamins|vitamin
Drug|Hormone|Past Medical History|1101,1110|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|vitamin D
Drug|Organic Chemical|Past Medical History|1101,1110|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|vitamin D
Drug|Pharmacologic Substance|Past Medical History|1101,1110|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|vitamin D
Drug|Vitamin|Past Medical History|1101,1110|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|vitamin D
Procedure|Laboratory Procedure|Past Medical History|1101,1110|false|false|false|C0919758|Vitamin D measurement|vitamin D
Disorder|Disease or Syndrome|Past Medical History|1101,1121|false|false|false|C0042870|Vitamin D Deficiency|vitamin D deficiency
Finding|Finding|Past Medical History|1101,1121|false|false|false|C5886864|Decreased circulating vitamin D concentration|vitamin D deficiency
Disorder|Disease or Syndrome|Past Medical History|1111,1121|false|false|false|C0162429|Malnutrition|deficiency
Finding|Functional Concept|Past Medical History|1111,1121|false|false|false|C0011155|Deficiency|deficiency
Finding|Intellectual Product|Past Medical History|1123,1131|false|false|false|C1522634|Question (inquiry)|question
Disorder|Disease or Syndrome|Past Medical History|1135,1149|false|false|false|C0020676|Hypothyroidism|hypothyroidism
Finding|Finding|Past Medical History|1155,1167|false|false|false|C0586553|Raised TSH level|elevated TSH
Attribute|Clinical Attribute|Past Medical History|1164,1167|false|false|false|C2708739||TSH
Drug|Amino Acid, Peptide, or Protein|Past Medical History|1164,1167|false|false|false|C0040160|thyrotropin|TSH
Drug|Hormone|Past Medical History|1164,1167|false|false|false|C0040160|thyrotropin|TSH
Drug|Pharmacologic Substance|Past Medical History|1164,1167|false|false|false|C0040160|thyrotropin|TSH
Procedure|Laboratory Procedure|Past Medical History|1164,1167|false|false|false|C0202230|Thyroid stimulating hormone measurement|TSH
Procedure|Laboratory Procedure|Past Medical History|1164,1173|false|false|false|C0202230|Thyroid stimulating hormone measurement|TSH level
Disorder|Disease or Syndrome|Past Medical History|1175,1186|false|false|false|C0039730|Thalassemia|thalassemia
Disorder|Disease or Syndrome|Past Medical History|1175,1192|false|false|false|C0702157|Thalassemia trait|thalassemia trait
Disorder|Disease or Syndrome|Past Medical History|1194,1205|false|false|false|C0015695;C2711227|Fatty Liver;Steatohepatitis|fatty liver
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1200,1205|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Past Medical History|1200,1205|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Past Medical History|1200,1205|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Past Medical History|1200,1205|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Past Medical History|1200,1205|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Past Medical History|1200,1205|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Finding|Finding|Past Medical History|1200,1205|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Past Medical History|1200,1205|false|false|false|C0872387|Procedures on liver|liver
Disorder|Disease or Syndrome|Past Medical History|1210,1224|false|false|false|C0008350|Cholelithiasis|cholelithiasis
Finding|Functional Concept|Past Medical History|1228,1238|false|false|false|C0220934|Ultrasonic|ultrasound
Phenomenon|Natural Phenomenon or Process|Past Medical History|1228,1238|false|false|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|ultrasound
Procedure|Diagnostic Procedure|Past Medical History|1228,1238|false|false|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|ultrasound
Finding|Intellectual Product|Past Medical History|1239,1244|false|false|false|C1705923|Study Object|study
Procedure|Research Activity|Past Medical History|1239,1244|false|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|study
Finding|Conceptual Entity|Past Medical History|1248,1255|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Past Medical History|1248,1255|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Past Medical History|1248,1255|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Past Medical History|1248,1258|false|false|false|C0262926|Medical History|history of
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1267,1274|false|false|false|C0040421;C0836921|Palatine Tonsil;Tonsil|tonsils
Procedure|Health Care Activity|Past Medical History|1267,1274|false|false|false|C2239123|examination of tonsils|tonsils
Finding|Functional Concept|Past Medical History|1300,1311|false|false|false|C0549186|Obstructed|obstructive
Disorder|Disease or Syndrome|Past Medical History|1300,1323|false|false|false|C0520679|Sleep Apnea, Obstructive|obstructive sleep apnea
Drug|Organic Chemical|Past Medical History|1312,1317|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Drug|Pharmacologic Substance|Past Medical History|1312,1317|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Finding|Organism Function|Past Medical History|1312,1317|false|false|false|C0037313|Sleep|sleep
Disorder|Disease or Syndrome|Past Medical History|1312,1323|false|false|false|C0037315|Sleep Apnea Syndromes|sleep apnea
Finding|Sign or Symptom|Past Medical History|1318,1323|false|false|false|C0003578|Apnea|apnea
Anatomy|Body Location or Region|Past Medical History|1328,1344|false|false|false|C0744316|gastroesophageal|gastroesophageal
Disorder|Disease or Syndrome|Past Medical History|1328,1351|false|false|false|C0017168|Gastroesophageal reflux disease|gastroesophageal reflux
Finding|Finding|Past Medical History|1328,1351|false|false|false|C3813607;C4317146|Acid reflux;Infantile Gastroesophageal Reflux|gastroesophageal reflux
Finding|Pathologic Function|Past Medical History|1345,1351|false|false|false|C0232483|Reflux|reflux
Finding|Conceptual Entity|Past Medical History|1364,1372|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolved
Finding|Pathologic Function|Past Medical History|1364,1372|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolved
Finding|Finding|Past Medical History|1364,1383|false|false|false|C5419890|Completely Resolved|resolved completely
Finding|Intellectual Product|Past Medical History|1373,1383|false|false|false|C4554154|Completely - dosing instruction fragment|completely
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1395,1408|false|false|false|C0040423|Tonsillectomy|tonsillectomy
Finding|Conceptual Entity|Past Medical History|1417,1424|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|Past Medical History|1417,1424|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|Past Medical History|1417,1424|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|Past Medical History|1417,1427|false|false|false|C0262926|Medical History|History of
Disorder|Disease or Syndrome|Past Medical History|1428,1444|false|false|false|C0032460|Polycystic Ovary Syndrome|polycystic ovary
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1439,1444|false|false|false|C0029939;C0227898;C4266530|Both ovaries;Ovary;Pelvis>Ovary|ovary
Disorder|Disease or Syndrome|Past Medical History|1439,1444|false|false|false|C0029928;C0496920|Neoplasm of uncertain or unknown behavior of ovary;Ovarian Diseases|ovary
Disorder|Neoplastic Process|Past Medical History|1439,1444|false|false|false|C0029928;C0496920|Neoplasm of uncertain or unknown behavior of ovary;Ovarian Diseases|ovary
Disorder|Disease or Syndrome|Past Medical History|1445,1453|false|false|false|C0039082|Syndrome|syndrome
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1492,1499|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|Family Medical History|1492,1499|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Procedure|Therapeutic or Preventive Procedure|Family Medical History|1492,1499|false|false|false|C0872388|Procedures on bladder|bladder
Disorder|Neoplastic Process|Family Medical History|1492,1502|false|true|false|C0005684|Malignant neoplasm of urinary bladder|bladder CA
Disorder|Disease or Syndrome|Family Medical History|1509,1517|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|diabetes
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1519,1525|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|Family Medical History|1519,1525|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Finding|Finding|Family Medical History|1519,1525|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|Family Medical History|1519,1525|false|false|false|C0191838|Procedures on breast|breast
Disorder|Neoplastic Process|Family Medical History|1526,1535|false|false|false|C0027651;C1882062|Neoplasms;Neoplastic disease|neoplasia
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1537,1542|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|Family Medical History|1537,1542|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|Family Medical History|1537,1542|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Finding|Finding|Family Medical History|1537,1542|false|false|false|C0750873|COLON PROBLEM|colon
Disorder|Neoplastic Process|Family Medical History|1537,1545|false|false|false|C0007102|Malignant tumor of colon|colon CA
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1547,1554|false|false|false|C0205065|Ovarian|ovarian
Disorder|Neoplastic Process|Family Medical History|1563,1570|false|false|false|C1261473;C4551686|Malignant neoplasm of soft tissue;Sarcoma|sarcoma
Finding|Gene or Genome|General Exam|1592,1596|false|false|false|C1823816|C1orf210 gene|Temp
Procedure|Therapeutic or Preventive Procedure|General Exam|1592,1596|false|false|false|C0279848|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Temp
Finding|Classification|General Exam|1648,1651|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|GEN
Finding|Gene or Genome|General Exam|1648,1651|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|GEN
Disorder|Disease or Syndrome|General Exam|1658,1661|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|1658,1661|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|1658,1661|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|1658,1661|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|1658,1661|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Finding|Finding|General Exam|1658,1661|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|General Exam|1662,1667|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|General Exam|1672,1679|false|false|false|C0036410|Sclera|scleral
Finding|Finding|General Exam|1672,1687|true|false|false|C0240962|Scleral icterus|scleral icterus
Finding|Sign or Symptom|General Exam|1680,1687|true|false|false|C0022346|Icterus|icterus
Anatomy|Body Part, Organ, or Organ Component|General Exam|1689,1692|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|General Exam|1689,1692|false|false|false|C0026987|Myelofibrosis|MMM
Procedure|Health Care Activity|General Exam|1701,1705|false|false|false|C1315068|Pulmonary ventilator management|PULM
Finding|Finding|General Exam|1720,1729|true|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Functional Concept|General Exam|1720,1729|true|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Sign or Symptom|General Exam|1720,1747|true|false|false|C0859927|Increased work of breathing|increased work of breathing
Event|Occupational Activity|General Exam|1730,1734|true|false|false|C0043227|Work|work
Finding|Organ or Tissue Function|General Exam|1730,1747|true|false|false|C0043229|Work of Breathing|work of breathing
Attribute|Clinical Attribute|General Exam|1738,1747|false|false|false|C5885990||breathing
Finding|Finding|General Exam|1738,1747|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|General Exam|1738,1747|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|General Exam|1738,1747|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|General Exam|1738,1747|false|false|false|C1160636|respiratory system process|breathing
Anatomy|Body Location or Region|General Exam|1748,1751|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|ABD
Disorder|Cell or Molecular Dysfunction|General Exam|1748,1751|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|ABD
Disorder|Disease or Syndrome|General Exam|1753,1757|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Procedure|Diagnostic Procedure|General Exam|1787,1796|false|false|false|C0030247|Palpation|palpation
Anatomy|Body Location or Region|General Exam|1800,1810|false|false|false|C0521440|Epigastric|epigastric
Drug|Amino Acid Sequence|General Exam|1812,1818|false|false|false|C1514562|Protein Domain|region
Finding|Finding|General Exam|1834,1842|true|false|false|C0427198|Protective muscle spasm|guarding
Drug|Food|General Exam|1853,1857|false|false|false|C0452253|Port - alcoholic beverage|port
Disorder|Congenital Abnormality|General Exam|1858,1861|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Finding|Gene or Genome|General Exam|1858,1861|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Attribute|Clinical Attribute|General Exam|1870,1875|false|false|false|C1717255||edema
Finding|Pathologic Function|General Exam|1870,1875|false|false|false|C0013604|Edema|edema
Finding|Finding|General Exam|1877,1881|false|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|General Exam|1877,1881|false|false|false|C0687712|warming process|warm
Finding|Finding|General Exam|1886,1890|false|false|false|C5575035|Well (answer to question)|well
Procedure|Laboratory Procedure|General Exam|1936,1939|false|false|false|C0201617|Primed lymphocyte test|PLT
Drug|Antibiotic|General Exam|1979,1984|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Biomedical or Dental Material|General Exam|1979,1984|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Organic Chemical|General Exam|1979,1984|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Disorder|Disease or Syndrome|General Exam|1989,1992|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|EOS
Finding|Gene or Genome|General Exam|1989,1992|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|EOS
Finding|Body Substance|General Exam|2125,2130|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|2125,2130|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|2125,2130|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Finding|General Exam|2125,2138|false|false|false|C0455910|Mucus in urine (finding)|URINE  MUCOUS
Finding|Body Substance|General Exam|2132,2138|false|false|false|C0026727;C2753459|Mucus (substance);mucus layer|MUCOUS
Finding|Gene or Genome|General Exam|2139,2143|false|false|false|C1514917|Retinoic Acid Response Element|RARE
Finding|Body Substance|General Exam|2156,2161|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|2156,2161|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|2156,2161|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Body Substance|General Exam|2163,2170|false|false|false|C0020191|Hyalin Substance|HYALINE
Finding|Body Substance|General Exam|2186,2191|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|2186,2191|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|2186,2191|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Lab|Laboratory or Test Result|General Exam|2186,2196|false|false|false|C0221752;C2188659|Red blood cells urine positive|URINE  RBC
Anatomy|Cell|General Exam|2193,2196|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|2193,2196|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|2193,2196|false|false|false|C0014792|Erythrocytes|RBC
Anatomy|Cell|General Exam|2200,2203|false|false|false|C0023516|Leukocytes|WBC
Finding|Functional Concept|General Exam|2206,2214|false|false|false|C1510439|bacteria aspects|BACTERIA
Disorder|Disease or Syndrome|General Exam|2215,2218|false|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|MOD
Drug|Food|General Exam|2219,2224|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Immunologic Factor|General Exam|2219,2224|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|2219,2224|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Pharmacologic Substance|General Exam|2219,2224|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Disorder|Disease or Syndrome|General Exam|2231,2234|false|false|false|C0267963|Exocrine pancreatic insufficiency|EPI
Drug|Amino Acid, Peptide, or Protein|General Exam|2231,2234|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Biologically Active Substance|General Exam|2231,2234|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Hormone|General Exam|2231,2234|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Organic Chemical|General Exam|2231,2234|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Pharmacologic Substance|General Exam|2231,2234|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Finding|Gene or Genome|General Exam|2231,2234|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|EPI
Finding|Intellectual Product|General Exam|2231,2234|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|EPI
Procedure|Diagnostic Procedure|General Exam|2231,2234|false|false|false|C0162734;C3641909|Echo-Planar Imaging;Electronic Portal Imaging|EPI
Finding|Body Substance|General Exam|2250,2255|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|2250,2255|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|2250,2255|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Disorder|Disease or Syndrome|General Exam|2250,2262|false|false|false|C0018965|Hematuria|URINE  BLOOD
Disorder|Disease or Syndrome|General Exam|2257,2262|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|2257,2262|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Finding|General Exam|2263,2266|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|General Exam|2267,2274|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Drug|Inorganic Chemical|General Exam|2267,2274|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Drug|Pharmacologic Substance|General Exam|2267,2274|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Finding|Finding|General Exam|2275,2278|false|false|false|C5848551|Neg - answer|NEG
Drug|Amino Acid, Peptide, or Protein|General Exam|2279,2286|false|false|false|C0033684|Proteins|PROTEIN
Drug|Biologically Active Substance|General Exam|2279,2286|false|false|false|C0033684|Proteins|PROTEIN
Finding|Conceptual Entity|General Exam|2279,2286|false|false|false|C1521746|Protein Info|PROTEIN
Procedure|Laboratory Procedure|General Exam|2279,2286|false|false|false|C0202202|Protein measurement|PROTEIN
Drug|Biologically Active Substance|General Exam|2291,2298|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|General Exam|2291,2298|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|General Exam|2291,2298|false|false|false|C0017725|glucose|GLUCOSE
Lab|Laboratory or Test Result|General Exam|2291,2298|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|General Exam|2291,2298|false|false|false|C0337438|Glucose measurement|GLUCOSE
Finding|Finding|General Exam|2299,2302|false|false|false|C5848551|Neg - answer|NEG
Drug|Organic Chemical|General Exam|2303,2309|false|false|false|C0022634|Ketones|KETONE
Finding|Finding|General Exam|2310,2313|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|General Exam|2314,2323|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Drug|Organic Chemical|General Exam|2314,2323|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Drug|Pharmacologic Substance|General Exam|2314,2323|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Procedure|Laboratory Procedure|General Exam|2314,2323|false|false|false|C0201913;C0863174|Bilirubin, total measurement;blood bilirubin level test|BILIRUBIN
Finding|Finding|General Exam|2324,2327|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|General Exam|2338,2341|false|false|false|C5848551|Neg - answer|NEG
Finding|Body Substance|General Exam|2370,2375|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|2370,2375|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|2370,2375|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Finding|General Exam|2370,2382|false|false|false|C0278030|Color of urine|URINE  COLOR
Drug|Biomedical or Dental Material|General Exam|2377,2382|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|COLOR
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|2377,2382|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|COLOR
Finding|Body Substance|General Exam|2421,2426|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|2421,2426|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|2421,2426|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Classification|General Exam|2432,2440|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Finding|Finding|General Exam|2432,2440|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Lab|Laboratory or Test Result|General Exam|2432,2440|false|false|false|C5237010|Expression Negative|NEGATIVE
Finding|Body Substance|General Exam|2453,2458|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|2453,2458|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|2453,2458|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Body Substance|General Exam|2485,2490|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|2485,2490|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|2485,2490|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Attribute|Clinical Attribute|Hospital Course|2566,2572|false|false|false|C4255480||nausea
Finding|Sign or Symptom|Hospital Course|2566,2572|false|false|false|C0027497|Nausea|nausea
Finding|Sign or Symptom|Hospital Course|2578,2586|false|false|false|C0042963|Vomiting|vomiting
Finding|Functional Concept|Hospital Course|2600,2606|false|false|false|C1512806|Intake|intake
Procedure|Health Care Activity|Hospital Course|2600,2606|false|false|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|intake
Finding|Idea or Concept|Hospital Course|2653,2657|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|Hospital Course|2653,2657|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Finding|Hospital Course|2675,2680|false|false|false|C3714655|On IV|on IV
Drug|Substance|Hospital Course|2681,2687|false|false|false|C0302908|Liquid substance|fluids
Finding|Body Substance|Hospital Course|2681,2687|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2681,2687|false|false|false|C0016286|Fluid Therapy|fluids
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2693,2704|false|false|false|C0034997|Rehydration|rehydration
Attribute|Clinical Attribute|Hospital Course|2710,2720|false|false|false|C2598148||laboratory
Finding|Functional Concept|Hospital Course|2710,2720|false|false|false|C1548427;C1571737;C3244292|Diagnostic Service Section ID - Laboratory;Laboratory domain;Referral type - Laboratory|laboratory
Finding|Intellectual Product|Hospital Course|2710,2720|false|false|false|C1548427;C1571737;C3244292|Diagnostic Service Section ID - Laboratory;Laboratory domain;Referral type - Laboratory|laboratory
Lab|Laboratory or Test Result|Hospital Course|2710,2720|false|false|false|C4283904|Laboratory observation|laboratory
Procedure|Health Care Activity|Hospital Course|2750,2759|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Functional Concept|Hospital Course|2768,2776|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Hospital Course|2768,2776|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Drug|Pharmacologic Substance|Hospital Course|2801,2812|false|false|false|C0003297;C3536993|Antiemetic [EPC];Antiemetics|anti-emetic
Attribute|Clinical Attribute|Hospital Course|2814,2825|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Hospital Course|2814,2825|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|Hospital Course|2814,2825|false|false|false|C4284232|Medications|medications
Drug|Substance|Hospital Course|2830,2838|false|false|false|C1289919|Intravenous fluid|IV fluid
Drug|Substance|Hospital Course|2833,2838|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|2833,2838|false|false|false|C1546638|Fluid Specimen Code|fluid
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2833,2846|false|false|false|C0016286;C0522792|Administration of intravenous fluids;Fluid Therapy|fluid therapy
Finding|Finding|Hospital Course|2839,2846|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|Hospital Course|2839,2846|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2839,2846|false|false|false|C0087111|Therapeutic procedure|therapy
Drug|Biomedical or Dental Material|Hospital Course|2868,2876|false|false|false|C0168634|BaseLine dental cement|baseline
Finding|Idea or Concept|Hospital Course|2868,2876|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Intellectual Product|Hospital Course|2878,2886|false|false|false|C1315013|Clinical NEC (not elsewhere classified in LNC)|clinical
Attribute|Clinical Attribute|Hospital Course|2878,2893|false|false|false|C0449440;C5890498|Clinical status|clinical status
Attribute|Clinical Attribute|Hospital Course|2887,2893|false|false|false|C5889824||status
Finding|Idea or Concept|Hospital Course|2887,2893|false|false|false|C1546481|What subject filter - Status|status
Drug|Inorganic Chemical|Hospital Course|2929,2934|false|false|false|C0043047;C1550678|Water Specimen;water|Water
Drug|Pharmacologic Substance|Hospital Course|2929,2934|false|false|false|C0043047;C1550678|Water Specimen;water|Water
Finding|Intellectual Product|Hospital Course|2929,2934|false|false|false|C1547961|Water - Specimen Source Codes|Water
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2929,2934|false|false|false|C0020311|Hydrotherapy|Water
Attribute|Clinical Attribute|Hospital Course|2936,2945|false|false|false|C0798503||challenge
Finding|Conceptual Entity|Hospital Course|2936,2945|false|false|false|C3274764|Proficiency Testing Challenge|challenge
Procedure|Health Care Activity|Hospital Course|2936,2945|false|false|false|C0805586|Challenge|challenge
Procedure|Laboratory Procedure|Hospital Course|2936,2950|false|false|false|C1315011|Challenge tests|challenge test
Anatomy|Body Location or Region|Hospital Course|2946,2950|false|false|false|C4318744|Test - temporal region|test
Finding|Functional Concept|Hospital Course|2946,2950|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|Hospital Course|2946,2950|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|Hospital Course|2946,2950|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|Hospital Course|2946,2950|false|false|false|C0022885|Laboratory Procedures|test
Finding|Classification|Hospital Course|2971,2981|false|false|false|C0376209;C0456081;C0678219;C0683269;C1546424|Adjustment - classification term;Personal Adjustment;Psychological adjustment;Transaction Type - Adjustment|adjustment
Finding|Functional Concept|Hospital Course|2971,2981|false|false|false|C0376209;C0456081;C0678219;C0683269;C1546424|Adjustment - classification term;Personal Adjustment;Psychological adjustment;Transaction Type - Adjustment|adjustment
Finding|Idea or Concept|Hospital Course|2971,2981|false|false|false|C0376209;C0456081;C0678219;C0683269;C1546424|Adjustment - classification term;Personal Adjustment;Psychological adjustment;Transaction Type - Adjustment|adjustment
Finding|Individual Behavior|Hospital Course|2971,2981|false|false|false|C0376209;C0456081;C0678219;C0683269;C1546424|Adjustment - classification term;Personal Adjustment;Psychological adjustment;Transaction Type - Adjustment|adjustment
Finding|Classification|Hospital Course|2990,2998|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|2990,2998|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|2990,2998|false|false|false|C5237010|Expression Negative|negative
Attribute|Clinical Attribute|Hospital Course|3008,3012|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|3008,3012|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|3008,3012|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|Hospital Course|3014,3020|false|false|false|C4255480||nausea
Finding|Sign or Symptom|Hospital Course|3014,3020|false|false|false|C0027497|Nausea|nausea
Finding|Finding|Hospital Course|3014,3032|false|false|false|C3843946|Nausea or vomiting|nausea or vomiting
Finding|Sign or Symptom|Hospital Course|3024,3032|true|false|false|C0042963|Vomiting|vomiting
Finding|Idea or Concept|Hospital Course|3056,3060|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Attribute|Clinical Attribute|Hospital Course|3062,3071|false|false|false|C3864998||condition
Disorder|Disease or Syndrome|Hospital Course|3062,3071|false|false|false|C0012634|Disease|condition
Finding|Conceptual Entity|Hospital Course|3062,3071|false|false|false|C1705253|Logical Condition|condition
Attribute|Clinical Attribute|Hospital Course|3077,3089|false|false|false|C3263700||instructions
Finding|Intellectual Product|Hospital Course|3077,3089|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|instructions
Finding|Body Substance|Hospital Course|3134,3143|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|3134,3143|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|3134,3143|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|3134,3143|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|3134,3155|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|3144,3155|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|3144,3155|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Hospital Course|3144,3155|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|3160,3169|false|false|false|C0024002|lorazepam|Lorazepam
Drug|Pharmacologic Substance|Hospital Course|3160,3169|false|false|false|C0024002|lorazepam|Lorazepam
Disorder|Mental or Behavioral Dysfunction|Hospital Course|3180,3183|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|3180,3183|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|3180,3183|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|3180,3183|false|false|false|C1332410|BID gene|BID
Finding|Gene or Genome|Hospital Course|3184,3187|false|false|false|C1422467|CIAO3 gene|PRN
Disorder|Mental or Behavioral Dysfunction|Hospital Course|3188,3195|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Finding|Sign or Symptom|Hospital Course|3188,3195|false|false|false|C0860603|Anxiety symptoms|anxiety
Drug|Organic Chemical|Hospital Course|3200,3209|false|false|false|C0006462|buspirone|BusPIRone
Drug|Pharmacologic Substance|Hospital Course|3200,3209|false|false|false|C0006462|buspirone|BusPIRone
Finding|Body Substance|Hospital Course|3226,3235|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|3226,3235|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|3226,3235|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|3226,3235|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|3226,3247|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|3226,3247|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|3236,3247|false|false|false|C2926604||Disposition
Procedure|Health Care Activity|Hospital Course|3236,3247|false|false|false|C0184758|Patient disposition|Disposition
Finding|Idea or Concept|Hospital Course|3249,3253|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|3249,3253|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|3249,3253|false|false|false|C1553498|home health encounter|Home
Finding|Body Substance|Hospital Course|3256,3265|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|3256,3265|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|3256,3265|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|3256,3265|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|3256,3275|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|3266,3275|false|false|false|C0945731||Diagnosis
Finding|Classification|Hospital Course|3266,3275|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|3266,3275|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|3266,3275|false|false|false|C0011900|Diagnosis|Diagnosis
Attribute|Clinical Attribute|Hospital Course|3277,3283|false|false|false|C4255480||nausea
Finding|Sign or Symptom|Hospital Course|3277,3283|false|false|false|C0027497|Nausea|nausea
Finding|Sign or Symptom|Hospital Course|3277,3296|false|false|false|C0027498|Nausea and vomiting|nausea and vomiting
Finding|Sign or Symptom|Hospital Course|3288,3296|false|false|false|C0042963|Vomiting|vomiting
Finding|Mental Process|Discharge Condition|3339,3345|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|3339,3352|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|3339,3352|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|3346,3352|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|3346,3352|false|false|false|C1546481|What subject filter - Status|Status
Finding|Idea or Concept|Discharge Condition|3354,3359|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Finding|Discharge Condition|3364,3372|false|false|false|C4068804|Coherent|coherent
Attribute|Clinical Attribute|Discharge Condition|3374,3396|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|3374,3396|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Finding|Finding|Discharge Condition|3383,3396|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|3383,3396|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|3398,3403|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|3398,3403|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|3398,3403|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|Discharge Condition|3398,3403|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|3398,3403|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|3398,3403|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|3408,3419|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|3421,3429|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|3421,3429|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|3421,3429|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|3430,3436|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|3430,3436|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|Discharge Condition|3438,3448|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|3438,3448|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|3438,3448|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|3438,3448|false|false|false|C1561560|ambulatory encounter|Ambulatory
Finding|Finding|Discharge Condition|3451,3462|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Condition|3451,3462|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Attribute|Clinical Attribute|Discharge Instructions|3525,3531|false|false|false|C4255480||Nausea
Finding|Sign or Symptom|Discharge Instructions|3525,3531|false|false|false|C0027497|Nausea|Nausea
Finding|Sign or Symptom|Discharge Instructions|3525,3544|false|false|false|C0027498|Nausea and vomiting|Nausea and vomiting
Finding|Sign or Symptom|Discharge Instructions|3536,3544|false|false|false|C0042963|Vomiting|vomiting
Attribute|Clinical Attribute|Discharge Instructions|3588,3594|false|false|false|C4255480||nausea
Finding|Sign or Symptom|Discharge Instructions|3588,3594|false|false|false|C0027497|Nausea|nausea
Finding|Sign or Symptom|Discharge Instructions|3588,3607|false|false|false|C0027498|Nausea and vomiting|nausea and vomiting
Finding|Sign or Symptom|Discharge Instructions|3599,3607|false|false|false|C0042963|Vomiting|vomiting
Finding|Functional Concept|Discharge Instructions|3672,3676|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Drug|Inorganic Chemical|Discharge Instructions|3708,3713|false|false|false|C0043047;C1550678|Water Specimen;water|water
Drug|Pharmacologic Substance|Discharge Instructions|3708,3713|false|false|false|C0043047;C1550678|Water Specimen;water|water
Finding|Intellectual Product|Discharge Instructions|3708,3713|false|false|false|C1547961|Water - Specimen Source Codes|water
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|3708,3713|false|false|false|C0020311|Hydrotherapy|water
Finding|Body Substance|Discharge Instructions|3714,3719|false|false|false|C1186706;C1550436|Bolus of ingested food;Response Modality - Bolus|bolus
Finding|Intellectual Product|Discharge Instructions|3714,3719|false|false|false|C1186706;C1550436|Bolus of ingested food;Response Modality - Bolus|bolus
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|3714,3719|false|false|false|C1511237|bolus infusion|bolus
Anatomy|Body Location or Region|Discharge Instructions|3720,3724|false|false|false|C4318744|Test - temporal region|test
Finding|Functional Concept|Discharge Instructions|3720,3724|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|Discharge Instructions|3720,3724|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|Discharge Instructions|3720,3724|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|Discharge Instructions|3720,3724|false|false|false|C0022885|Laboratory Procedures|test
Finding|Idea or Concept|Discharge Instructions|3778,3786|false|false|false|C1547192|Organization unit type - Hospital|hospital
Attribute|Clinical Attribute|Discharge Instructions|3811,3817|false|false|false|C4255480||nausea
Finding|Sign or Symptom|Discharge Instructions|3811,3817|false|false|false|C0027497|Nausea|nausea
Finding|Sign or Symptom|Discharge Instructions|3851,3859|false|false|false|C0042963|Vomiting|vomiting
Finding|Idea or Concept|Discharge Instructions|3896,3900|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Discharge Instructions|3896,3900|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Discharge Instructions|3896,3900|false|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|Discharge Instructions|3901,3912|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|3901,3912|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|Discharge Instructions|3901,3912|false|false|false|C4284232|Medications|medications
Procedure|Health Care Activity|Discharge Instructions|3959,3969|false|false|false|C0086388|Health Care|healthcare
Procedure|Health Care Activity|Discharge Instructions|3975,3983|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|3984,3996|false|false|false|C3263700||Instructions
Finding|Intellectual Product|Discharge Instructions|3984,3996|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

