 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|22,26
No|27,29
:|29,30
_|33,34
_|34,35
_|35,36
<EOL>|36,37
<EOL>|38,39
Admission|39,48
Date|49,53
:|53,54
_|56,57
_|57,58
_|58,59
Discharge|73,82
Date|83,87
:|87,88
_|91,92
_|92,93
_|93,94
<EOL>|94,95
<EOL>|96,97
Date|97,101
of|102,104
Birth|105,110
:|110,111
_|113,114
_|114,115
_|115,116
Sex|129,132
:|132,133
F|136,137
<EOL>|137,138
<EOL>|139,140
Service|140,147
:|147,148
MEDICINE|149,157
<EOL>|157,158
<EOL>|159,160
Allergies|160,169
:|169,170
<EOL>|171,172
No|172,174
Known|175,180
Allergies|181,190
/|191,192
Adverse|193,200
Drug|201,205
Reactions|206,215
<EOL>|215,216
<EOL>|217,218
Attending|218,227
:|227,228
_|229,230
_|230,231
_|231,232
.|232,233
<EOL>|233,234
<EOL>|235,236
Chief|236,241
Complaint|242,251
:|251,252
<EOL>|252,253
shortness|253,262
of|263,265
breath|266,272
<EOL>|272,273
<EOL>|274,275
Major|275,280
Surgical|281,289
or|290,292
Invasive|293,301
Procedure|302,311
:|311,312
<EOL>|312,313
None|313,317
<EOL>|317,318
<EOL>|318,319
<EOL>|320,321
History|321,328
of|329,331
Present|332,339
Illness|340,347
:|347,348
<EOL>|348,349
Patient|349,356
is|357,359
a|360,361
_|362,363
_|363,364
_|364,365
with|366,370
history|371,378
of|379,381
coronary|382,390
artery|391,397
disease|398,405
c|406,407
/|407,408
b|408,409
<EOL>|409,410
ischemic|410,418
MR|419,421
_|422,423
_|423,424
_|424,425
DES|426,429
to|430,432
LCX|433,436
_|437,438
_|438,439
_|439,440
,|440,441
TTE|442,445
_|446,447
_|447,448
_|448,449
with|450,454
mild|455,459
regional|460,468
LV|469,471
<EOL>|471,472
systolic|472,480
dysfunction|481,492
)|492,493
,|493,494
heart|495,500
failure|501,508
with|509,513
preserved|514,523
ejection|524,532
<EOL>|532,533
fraction|533,541
(|542,543
LVEF|543,547
50|548,550
%|550,551
_|552,553
_|553,554
_|554,555
,|555,556
peripheral|557,567
vascular|568,576
disease|577,584
,|584,585
chronic|586,593
<EOL>|593,594
kidney|594,600
disease|601,608
(|609,610
stage|610,615
IV|616,618
)|618,619
,|619,620
prior|621,626
unprovoked|627,637
DVT|638,641
c|642,643
/|643,644
b|644,645
severe|646,652
UGIB|653,657
<EOL>|657,658
while|658,663
on|664,666
AC|667,669
,|669,670
HTN|671,674
,|674,675
dyslipidemia|676,688
,|688,689
and|690,693
T2DM|694,698
who|699,702
presents|703,711
with|712,716
<EOL>|716,717
several|717,724
days|725,729
of|730,732
shortness|733,742
of|743,745
breath|746,752
.|752,753
<EOL>|758,759
<EOL>|759,760
Patients|760,768
says|769,773
that|774,778
she|779,782
first|783,788
noticed|789,796
rather|797,803
acute|804,809
onset|810,815
dyspnea|816,823
<EOL>|823,824
starting|824,832
_|833,834
_|834,835
_|835,836
when|837,841
trying|842,848
to|849,851
walk|852,856
up|857,859
the|860,863
stairs|864,870
in|871,873
her|874,877
home|878,882
.|882,883
<EOL>|884,885
<EOL>|885,886
She|886,889
had|890,893
to|894,896
sit|897,900
down|901,905
and|906,909
catch|910,915
her|916,919
breath|920,926
,|926,927
whereas|928,935
just|936,940
days|941,945
<EOL>|946,947
prior|947,952
<EOL>|952,953
she|953,956
was|957,960
able|961,965
to|966,968
mount|969,974
_|975,976
_|976,977
_|977,978
of|979,981
stairs|982,988
without|989,996
difficulty|997,1007
.|1007,1008
<EOL>|1009,1010
Patient|1010,1017
denies|1018,1024
any|1025,1028
associated|1029,1039
chest|1040,1045
pain|1046,1050
or|1051,1053
palpitations|1054,1066
.|1066,1067
No|1069,1071
<EOL>|1071,1072
dizziness|1072,1081
or|1082,1084
lightheadedness|1085,1100
.|1100,1101
Patient|1103,1110
further|1111,1118
denies|1119,1125
any|1126,1129
cough|1130,1135
,|1135,1136
<EOL>|1136,1137
fevers|1137,1143
/|1143,1144
chills|1144,1150
,|1150,1151
or|1152,1154
pleuritic|1155,1164
chest|1165,1170
discomfort|1171,1181
.|1181,1182
She|1184,1187
has|1188,1191
not|1192,1195
<EOL>|1195,1196
experienced|1196,1207
any|1208,1211
symptoms|1212,1220
consistent|1221,1231
with|1232,1236
orthopnea|1237,1246
or|1247,1249
PND|1250,1253
.|1253,1254
No|1256,1258
<EOL>|1258,1259
increased|1259,1268
_|1269,1270
_|1270,1271
_|1271,1272
swelling|1273,1281
,|1281,1282
patient|1283,1290
notes|1291,1296
that|1297,1301
she|1302,1305
has|1306,1309
experienced|1310,1321
<EOL>|1321,1322
this|1322,1326
in|1327,1329
the|1330,1333
past|1334,1338
.|1338,1339
<EOL>|1341,1342
<EOL>|1342,1343
Patient|1343,1350
takes|1351,1356
her|1357,1360
weight|1361,1367
nearly|1368,1374
every|1375,1380
day|1381,1384
,|1384,1385
7lbs|1386,1390
reported|1391,1399
weight|1400,1406
<EOL>|1406,1407
gain|1407,1411
over|1412,1416
the|1417,1420
past|1421,1425
week|1426,1430
(|1431,1432
154lbs|1432,1438
-|1439,1440
>|1440,1441
161lbs|1442,1448
)|1448,1449
,|1449,1450
which|1451,1456
she|1457,1460
attributes|1461,1471
<EOL>|1471,1472
to|1472,1474
eating|1475,1481
more|1482,1486
over|1487,1491
the|1492,1495
_|1496,1497
_|1497,1498
_|1498,1499
.|1499,1500
She|1502,1505
is|1506,1508
currently|1509,1518
<EOL>|1518,1519
taking|1519,1525
torsemide|1526,1535
40mg|1536,1540
qd|1541,1543
,|1543,1544
no|1545,1547
missed|1548,1554
doses|1555,1560
.|1560,1561
No|1563,1565
issues|1566,1572
with|1573,1577
<EOL>|1577,1578
abdominal|1578,1587
bloating|1588,1596
or|1597,1599
constipation|1600,1612
.|1612,1613
No|1615,1617
recent|1618,1624
travel|1625,1631
.|1631,1632
<EOL>|1634,1635
Patient|1635,1642
's|1642,1644
<EOL>|1644,1645
husband|1645,1652
just|1653,1657
recovered|1658,1667
from|1668,1672
a|1673,1674
viral|1675,1680
URI|1681,1684
.|1684,1685
<EOL>|1692,1693
<EOL>|1693,1694
In|1694,1696
the|1697,1700
ED|1701,1703
,|1703,1704
initial|1705,1712
VS|1713,1715
were|1716,1720
:|1720,1721
97.2|1722,1726
90|1727,1729
186|1730,1733
/|1733,1734
87|1734,1736
22|1737,1739
100|1740,1743
%|1743,1744
RA|1745,1747
<EOL>|1750,1751
<EOL>|1751,1752
Exam|1752,1756
notable|1757,1764
for|1765,1768
:|1768,1769
<EOL>|1769,1770
Obvious|1770,1777
bilateral|1778,1787
wheezing|1788,1796
.|1796,1797
<EOL>|1797,1798
No|1798,1800
overt|1801,1806
volume|1807,1813
overload|1814,1822
.|1822,1823
<EOL>|1825,1826
<EOL>|1826,1827
EKG|1827,1830
:|1830,1831
NSR|1832,1835
(|1836,1837
92bpm|1837,1842
)|1842,1843
,|1843,1844
normal|1845,1851
axis|1852,1856
,|1856,1857
normal|1858,1864
PR|1865,1867
/|1867,1868
QRS|1868,1871
intervals|1872,1881
,|1881,1882
QTc|1883,1886
479|1887,1890
,|1890,1891
<EOL>|1891,1892
q|1892,1893
-|1893,1894
waves|1894,1899
III|1900,1903
/|1903,1904
aVF|1904,1907
,|1907,1908
TWIs|1909,1913
III|1914,1917
/|1917,1918
aVF|1918,1921
/|1921,1922
V3|1922,1924
/|1924,1925
V6|1925,1927
,|1927,1928
submm|1929,1934
lateral|1935,1942
STDs|1943,1947
,|1947,1948
no|1949,1951
<EOL>|1952,1953
STEs|1953,1957
.|1957,1958
<EOL>|1958,1959
<EOL>|1959,1960
Labs|1960,1964
showed|1965,1971
:|1971,1972
<EOL>|1974,1975
CBC|1975,1978
6.0|1979,1982
>|1982,1983
9.0|1983,1986
/|1986,1987
27|1987,1989
.|1989,1990
8|1990,1991
<|1991,1992
176|1992,1995
(|1996,1997
PMNs|1997,2001
75.2|2002,2006
%|2006,2007
,|2007,2008
MCV|2009,2012
97|2013,2015
)|2015,2016
<EOL>|2016,2017
BMP|2017,2020
142|2021,2024
/|2024,2025
4.8|2025,2028
/|2028,2029
105|2029,2032
/|2032,2033
_|2033,2034
_|2034,2035
_|2035,2036
/|2036,2037
2|2037,2038
.|2038,2039
4|2039,2040
/|2040,2041
189|2041,2044
<EOL>|2044,2045
Trop|2045,2049
<|2050,2051
.01|2051,2054
<EOL>|2054,2055
proBNP|2055,2061
4512|2062,2066
<EOL>|2066,2067
VBG|2067,2070
7.33|2071,2075
/|2075,2076
40|2076,2078
<EOL>|2078,2079
UA|2079,2081
:|2081,2082
1.010|2083,2088
SG|2089,2091
,|2091,2092
pH|2093,2095
6.0|2096,2099
,|2099,2100
urobilinogen|2101,2113
NEG|2114,2117
,|2117,2118
bilirubin|2119,2128
NEG|2129,2132
,|2132,2133
leuk|2134,2138
NEG|2139,2142
,|2142,2143
<EOL>|2143,2144
blood|2144,2149
NEG|2150,2153
,|2153,2154
nitrite|2155,2162
NEG|2163,2166
,|2166,2167
protein|2168,2175
100|2176,2179
,|2179,2180
glucose|2181,2188
NEG|2189,2192
,|2192,2193
ketones|2194,2201
NEG|2202,2205
,|2205,2206
<EOL>|2206,2207
RBC|2207,2210
1|2211,2212
,|2212,2213
WBC|2214,2217
1|2218,2219
,|2219,2220
few|2221,2224
bacteria|2225,2233
<EOL>|2233,2234
<EOL>|2234,2235
Imaging|2235,2242
showed|2243,2249
:|2249,2250
<EOL>|2251,2252
CXR|2252,2255
_|2256,2257
_|2257,2258
_|2258,2259
<EOL>|2259,2260
FINDINGS|2260,2268
:|2268,2269
<EOL>|2271,2272
Lungs|2272,2277
are|2278,2281
moderately|2282,2292
well|2293,2297
-|2297,2298
expanded|2298,2306
.|2306,2307
There|2308,2313
is|2314,2316
an|2317,2319
asymmetric|2320,2330
right|2331,2336
<EOL>|2336,2337
lower|2337,2342
lung|2343,2347
opacity|2348,2355
,|2355,2356
new|2357,2360
from|2361,2365
_|2366,2367
_|2367,2368
_|2368,2369
.|2369,2370
The|2371,2374
heart|2375,2380
appears|2381,2388
mildly|2389,2395
<EOL>|2395,2396
enlarged|2396,2404
and|2405,2408
there|2409,2414
is|2415,2417
mild|2418,2422
pulmonary|2423,2432
vascular|2433,2441
congestion|2442,2452
.|2452,2453
No|2454,2456
<EOL>|2456,2457
pleural|2457,2464
effusion|2465,2473
or|2474,2476
pneumothorax|2477,2489
.|2489,2490
<EOL>|2491,2492
IMPRESSION|2492,2502
:|2502,2503
<EOL>|2505,2506
Right|2506,2511
lower|2512,2517
lobe|2518,2522
opacity|2523,2530
could|2531,2536
represent|2537,2546
pneumonia|2547,2556
in|2557,2559
the|2560,2563
right|2564,2569
<EOL>|2569,2570
clinical|2570,2578
setting|2579,2586
,|2586,2587
although|2588,2596
atelectasis|2597,2608
or|2609,2611
asymmetric|2612,2622
pulmonary|2623,2632
<EOL>|2632,2633
edema|2633,2638
could|2639,2644
account|2645,2652
for|2653,2656
this|2657,2661
finding|2662,2669
.|2669,2670
Dedicated|2671,2680
PA|2681,2683
and|2684,2687
lateral|2688,2695
<EOL>|2695,2696
views|2696,2701
could|2702,2707
be|2708,2710
helpful|2711,2718
for|2719,2722
further|2723,2730
assessment|2731,2741
.|2741,2742
<EOL>|2743,2744
<EOL>|2745,2746
Consults|2746,2754
:|2754,2755
NONE|2756,2760
<EOL>|2762,2763
<EOL>|2763,2764
Patient|2764,2771
received|2772,2780
:|2780,2781
<EOL>|2783,2784
_|2784,2785
_|2785,2786
_|2786,2787
21|2788,2790
:|2790,2791
45|2791,2793
IH|2794,2796
Albuterol|2797,2806
0.083|2807,2812
%|2812,2813
Neb|2814,2817
Soln|2818,2822
1|2823,2824
NEB|2825,2828
<EOL>|2830,2831
_|2831,2832
_|2832,2833
_|2833,2834
22|2835,2837
:|2837,2838
08|2838,2840
IH|2841,2843
Albuterol|2844,2853
0.083|2854,2859
%|2859,2860
Neb|2861,2864
Soln|2865,2869
1|2870,2871
NEB|2872,2875
<EOL>|2877,2878
_|2878,2879
_|2879,2880
_|2880,2881
22|2882,2884
:|2884,2885
08|2885,2887
IH|2888,2890
Ipratropium|2891,2902
Bromide|2903,2910
Neb|2911,2914
1|2915,2916
NEB|2917,2920
<EOL>|2922,2923
_|2923,2924
_|2924,2925
_|2925,2926
22|2927,2929
:|2929,2930
47|2930,2932
IH|2933,2935
Albuterol|2936,2945
0.083|2946,2951
%|2951,2952
Neb|2953,2956
Soln|2957,2961
1|2962,2963
NEB|2964,2967
<EOL>|2968,2969
_|2969,2970
_|2970,2971
_|2971,2972
22|2973,2975
:|2975,2976
47|2976,2978
IH|2979,2981
Ipratropium|2982,2993
Bromide|2994,3001
Neb|3002,3005
1|3006,3007
NEB|3008,3011
<EOL>|3012,3013
_|3013,3014
_|3014,3015
_|3015,3016
22|3017,3019
:|3019,3020
51|3020,3022
IV|3023,3025
Azithromycin|3026,3038
<EOL>|3039,3040
_|3040,3041
_|3041,3042
_|3042,3043
22|3044,3046
:|3046,3047
51|3047,3049
IV|3050,3052
CefTRIAXone|3053,3064
<EOL>|3064,3065
_|3065,3066
_|3066,3067
_|3067,3068
22|3069,3071
:|3071,3072
51|3072,3074
PO|3075,3077
PredniSONE|3078,3088
60|3089,3091
mg|3092,3094
<EOL>|3094,3095
_|3095,3096
_|3096,3097
_|3097,3098
22|3099,3101
:|3101,3102
51|3102,3104
IV|3105,3107
Furosemide|3108,3118
80|3119,3121
mg|3122,3124
<EOL>|3125,3126
_|3126,3127
_|3127,3128
_|3128,3129
23|3130,3132
:|3132,3133
01|3133,3135
IV|3136,3138
CefTRIAXone|3139,3150
1|3151,3152
gm|3153,3155
<EOL>|3157,3158
_|3158,3159
_|3159,3160
_|3160,3161
00|3162,3164
:|3164,3165
13|3165,3167
IV|3168,3170
Azithromycin|3171,3183
500|3184,3187
mg|3188,3190
<EOL>|3190,3191
_|3191,3192
_|3192,3193
_|3193,3194
00|3195,3197
:|3197,3198
23|3198,3200
PO|3201,3203
/|3203,3204
NG|3204,3206
Atorvastatin|3207,3219
80|3220,3222
mg|3223,3225
<EOL>|3225,3226
_|3226,3227
_|3227,3228
_|3228,3229
00|3230,3232
:|3232,3233
23|3233,3235
PO|3236,3238
/|3238,3239
NG|3239,3241
Carvedilol|3242,3252
25|3253,3255
mg|3256,3258
<EOL>|3258,3259
_|3259,3260
_|3260,3261
_|3261,3262
00|3263,3265
:|3265,3266
23|3266,3268
PO|3269,3271
NIFEdipine|3272,3282
(|3283,3284
Extended|3284,3292
Release|3293,3300
)|3300,3301
60|3302,3304
mg|3305,3307
<EOL>|3308,3309
_|3309,3310
_|3310,3311
_|3311,3312
00|3313,3315
:|3315,3316
23|3316,3318
IH|3319,3321
Albuterol|3322,3331
0.083|3332,3337
%|3337,3338
Neb|3339,3342
Soln|3343,3347
1|3348,3349
NEB|3350,3353
<EOL>|3354,3355
_|3355,3356
_|3356,3357
_|3357,3358
00|3359,3361
:|3361,3362
23|3362,3364
IH|3365,3367
Ipratropium|3368,3379
Bromide|3380,3387
Neb|3388,3391
1|3392,3393
NEB|3394,3397
<EOL>|3397,3398
_|3398,3399
_|3399,3400
_|3400,3401
00|3402,3404
:|3404,3405
26|3405,3407
PO|3408,3410
/|3410,3411
NG|3411,3413
Gabapentin|3414,3424
100|3425,3428
mg|3429,3431
<EOL>|3431,3432
_|3432,3433
_|3433,3434
_|3434,3435
00|3436,3438
:|3438,3439
44|3439,3441
SC|3442,3444
Insulin|3445,3452
4|3453,3454
Units|3455,3460
<EOL>|3460,3461
<EOL>|3461,3462
Transfer|3462,3470
VS|3471,3473
were|3474,3478
:|3478,3479
98.2|3480,3484
77|3485,3487
141|3488,3491
/|3491,3492
76|3492,3494
18|3495,3497
100|3498,3501
%|3501,3502
2L|3503,3505
NC|3506,3508
<EOL>|3509,3510
<EOL>|3513,3514
On|3514,3516
arrival|3517,3524
to|3525,3527
the|3528,3531
floor|3532,3537
,|3537,3538
patient|3539,3546
recounts|3547,3555
the|3556,3559
history|3560,3567
as|3568,3570
above|3571,3576
.|3576,3577
<EOL>|3578,3579
She|3579,3582
says|3583,3587
that|3588,3592
she|3593,3596
feels|3597,3602
improved|3603,3611
after|3612,3617
treatment|3618,3627
in|3628,3630
the|3631,3634
ED|3635,3637
,|3637,3638
no|3639,3641
<EOL>|3641,3642
ongoing|3642,3649
SOB|3650,3653
.|3653,3654
<EOL>|3655,3656
<EOL>|3657,3658
10|3658,3660
-|3660,3661
point|3661,3666
ROS|3667,3670
is|3671,3673
otherwise|3674,3683
NEGATIVE|3684,3692
.|3692,3693
<EOL>|3693,3694
<EOL>|3694,3695
<EOL>|3696,3697
Past|3697,3701
Medical|3702,3709
History|3710,3717
:|3717,3718
<EOL>|3718,3719
Coronary|3719,3727
artery|3728,3734
disease|3735,3742
<EOL>|3742,3743
Peripheral|3743,3753
vascular|3754,3762
disease|3763,3770
<EOL>|3770,3771
Type|3771,3775
II|3776,3778
Diabetes|3779,3787
Mellitus|3788,3796
c|3797,3798
/|3798,3799
b|3799,3800
diabetic|3801,3809
retinopathy|3810,3821
<EOL>|3821,3822
Obesity|3822,3829
<EOL>|3829,3830
Esophageal|3830,3840
ring|3841,3845
<EOL>|3845,3846
Hypertension|3846,3858
<EOL>|3858,3859
Dyslipidemia|3859,3871
<EOL>|3871,3872
Bilateral|3872,3881
unprovoked|3882,3892
posterior|3893,3902
tibial|3903,3909
DVTs|3910,3914
(|3915,3916
_|3916,3917
_|3917,3918
_|3918,3919
)|3919,3920
off|3921,3924
AC|3925,3927
given|3928,3933
<EOL>|3933,3934
severe|3934,3940
UGIB|3941,3945
<EOL>|3945,3946
CKD|3946,3949
Stage|3950,3955
IV|3956,3958
iso|3959,3962
DM|3963,3965
/|3965,3966
HTN|3966,3969
,|3969,3970
secondary|3971,3980
hyperparathyroidism|3981,4000
<EOL>|4000,4001
Anemia|4001,4007
<EOL>|4007,4008
Gout|4008,4012
<EOL>|4012,4013
<EOL>|4014,4015
Social|4015,4021
History|4022,4029
:|4029,4030
<EOL>|4030,4031
_|4031,4032
_|4032,4033
_|4033,4034
<EOL>|4034,4035
Family|4035,4041
History|4042,4049
:|4049,4050
<EOL>|4050,4051
Niece|4051,4056
had|4057,4060
some|4061,4065
sort|4066,4070
of|4071,4073
cancer|4074,4080
.|4080,4081
Father|4082,4088
died|4089,4093
in|4094,4096
his|4097,4100
_|4101,4102
_|4102,4103
_|4103,4104
due|4105,4108
to|4109,4111
<EOL>|4112,4113
lung|4113,4117
disease|4118,4125
.|4125,4126
Mother|4127,4133
died|4134,4138
in|4139,4141
her|4142,4145
_|4146,4147
_|4147,4148
_|4148,4149
due|4150,4153
to|4154,4156
an|4157,4159
unknown|4160,4167
cause|4168,4173
.|4173,4174
<EOL>|4175,4176
No|4176,4178
early|4179,4184
CAD|4185,4188
or|4189,4191
sudden|4192,4198
cardiac|4199,4206
death|4207,4212
.|4212,4213
No|4214,4216
other|4217,4222
known|4223,4228
history|4229,4236
of|4237,4239
<EOL>|4240,4241
cancer|4241,4247
.|4247,4248
<EOL>|4249,4250
<EOL>|4251,4252
Physical|4252,4260
Exam|4261,4265
:|4265,4266
<EOL>|4266,4267
=|4267,4268
=|4268,4269
=|4269,4270
=|4270,4271
=|4271,4272
=|4272,4273
=|4273,4274
=|4274,4275
=|4275,4276
=|4276,4277
=|4277,4278
=|4278,4279
=|4279,4280
=|4280,4281
=|4281,4282
=|4282,4283
=|4283,4284
=|4284,4285
=|4285,4286
=|4286,4287
=|4287,4288
=|4288,4289
=|4289,4290
=|4290,4291
=|4291,4292
=|4292,4293
=|4293,4294
=|4294,4295
=|4295,4296
=|4296,4297
<EOL>|4297,4298
ADMISSION|4299,4308
PHYSICAL|4309,4317
EXAM|4318,4322
<EOL>|4322,4323
=|4323,4324
=|4324,4325
=|4325,4326
=|4326,4327
=|4327,4328
=|4328,4329
=|4329,4330
=|4330,4331
=|4331,4332
=|4332,4333
=|4333,4334
=|4334,4335
=|4335,4336
=|4336,4337
=|4337,4338
=|4338,4339
=|4339,4340
=|4340,4341
=|4341,4342
=|4342,4343
=|4343,4344
=|4344,4345
=|4345,4346
=|4346,4347
=|4347,4348
=|4348,4349
=|4349,4350
=|4350,4351
=|4351,4352
=|4352,4353
<EOL>|4353,4354
VS|4354,4356
:|4356,4357
97.5|4358,4362
162|4363,4366
/|4366,4367
93|4367,4369
78|4370,4372
16|4373,4375
100RA|4376,4381
<EOL>|4384,4385
GENERAL|4385,4392
:|4392,4393
Pleasant|4394,4402
female|4403,4409
appearing|4410,4419
younger|4420,4427
than|4428,4432
her|4433,4436
stated|4437,4443
age|4444,4447
,|4447,4448
<EOL>|4448,4449
taking|4449,4455
deep|4456,4460
breaths|4461,4468
while|4469,4474
speaking|4475,4483
<EOL>|4485,4486
HEENT|4486,4491
:|4491,4492
EOMI|4493,4497
,|4497,4498
PERRL|4499,4504
,|4504,4505
anicteric|4506,4515
sclera|4516,4522
,|4522,4523
pink|4524,4528
conjunctiva|4529,4540
,|4540,4541
MMM|4542,4545
.|4545,4546
<EOL>|4548,4549
NECK|4549,4553
:|4553,4554
JVD|4555,4558
10|4559,4561
CM|4562,4564
.|4564,4565
<EOL>|4566,4567
HEART|4567,4572
:|4572,4573
RRR|4574,4577
,|4577,4578
S1|4579,4581
/|4581,4582
S2|4582,4584
,|4584,4585
no|4586,4588
murmurs|4589,4596
,|4596,4597
gallops|4598,4605
,|4605,4606
or|4607,4609
rubs|4610,4614
.|4614,4615
<EOL>|4617,4618
LUNGS|4618,4623
:|4623,4624
CTAB|4625,4629
,|4629,4630
no|4631,4633
wheezes|4634,4641
.|4641,4642
<EOL>|4643,4644
ABDOMEN|4644,4651
:|4651,4652
Obese|4653,4658
abdomen|4659,4666
,|4666,4667
normoactive|4668,4679
BS|4680,4682
throughout|4683,4693
,|4693,4694
nondistended|4695,4707
,|4707,4708
<EOL>|4708,4709
nontender|4709,4718
in|4719,4721
all|4722,4725
quadrants|4726,4735
,|4735,4736
no|4737,4739
rebound|4740,4747
/|4747,4748
guarding|4748,4756
,|4756,4757
no|4758,4760
<EOL>|4760,4761
hepatosplenomegaly|4761,4779
.|4779,4780
<EOL>|4782,4783
EXTREMITIES|4783,4794
:|4794,4795
No|4796,4798
cyanosis|4799,4807
,|4807,4808
clubbing|4809,4817
,|4817,4818
or|4819,4821
edema|4822,4827
.|4827,4828
<EOL>|4830,4831
PULSES|4831,4837
:|4837,4838
2|4839,4840
+|4840,4841
radial|4842,4848
pulses|4849,4855
bilaterally|4856,4867
.|4867,4868
<EOL>|4870,4871
NEURO|4871,4876
:|4876,4877
A|4878,4879
&|4879,4880
Ox3|4880,4883
,|4883,4884
moving|4885,4891
all|4892,4895
4|4896,4897
extremities|4898,4909
with|4910,4914
purpose|4915,4922
.|4922,4923
<EOL>|4925,4926
SKIN|4926,4930
:|4930,4931
Warm|4932,4936
and|4937,4940
well|4941,4945
perfused|4946,4954
,|4954,4955
no|4956,4958
excoriations|4959,4971
or|4972,4974
lesions|4975,4982
,|4982,4983
no|4984,4986
<EOL>|4986,4987
rashes|4987,4993
.|4993,4994
<EOL>|4996,4997
<EOL>|4998,4999
=|4999,5000
=|5000,5001
=|5001,5002
=|5002,5003
=|5003,5004
=|5004,5005
=|5005,5006
=|5006,5007
=|5007,5008
=|5008,5009
=|5009,5010
=|5010,5011
=|5011,5012
=|5012,5013
=|5013,5014
=|5014,5015
=|5015,5016
=|5016,5017
=|5017,5018
=|5018,5019
=|5019,5020
=|5020,5021
=|5021,5022
=|5022,5023
=|5023,5024
=|5024,5025
=|5025,5026
=|5026,5027
=|5027,5028
=|5028,5029
<EOL>|5029,5030
DISCHARGE|5030,5039
PHYSICAL|5040,5048
EXAM|5049,5053
<EOL>|5053,5054
=|5054,5055
=|5055,5056
=|5056,5057
=|5057,5058
=|5058,5059
=|5059,5060
=|5060,5061
=|5061,5062
=|5062,5063
=|5063,5064
=|5064,5065
=|5065,5066
=|5066,5067
=|5067,5068
=|5068,5069
=|5069,5070
=|5070,5071
=|5071,5072
=|5072,5073
=|5073,5074
=|5074,5075
=|5075,5076
=|5076,5077
=|5077,5078
=|5078,5079
=|5079,5080
=|5080,5081
=|5081,5082
=|5082,5083
=|5083,5084
<EOL>|5084,5085
VS|5085,5087
:|5087,5088
Afeb|5089,5093
,|5093,5094
144|5095,5098
/|5098,5099
78|5099,5101
,|5101,5102
HR|5103,5105
57|5106,5108
,|5108,5109
97|5110,5112
%|5112,5113
RA|5114,5116
,|5116,5117
RR|5118,5120
12|5121,5123
<EOL>|5123,5124
GEN|5124,5127
:|5127,5128
Well|5129,5133
appearing|5134,5143
in|5144,5146
NAD|5147,5150
<EOL>|5150,5151
Neck|5151,5155
:|5155,5156
No|5158,5160
JVD|5161,5164
appreciated|5165,5176
<EOL>|5176,5177
CV|5177,5179
:|5179,5180
RRR|5181,5184
no|5185,5187
m|5188,5189
/|5189,5190
r|5190,5191
/|5191,5192
g|5192,5193
,|5193,5194
no|5195,5197
carotid|5198,5205
bruits|5206,5212
appreciated|5213,5224
<EOL>|5224,5225
PULM|5225,5229
:|5229,5230
CTAB|5231,5235
no|5236,5238
wheezes|5239,5246
,|5246,5247
rales|5248,5253
,|5253,5254
or|5255,5257
crackles|5258,5266
.|5266,5267
Symmetric|5269,5278
expansion|5279,5288
<EOL>|5288,5289
EXT|5289,5292
:|5292,5293
warm|5294,5298
well|5299,5303
perfused|5304,5312
,|5312,5313
no|5314,5316
pitting|5317,5324
edema|5325,5330
<EOL>|5331,5332
<EOL>|5333,5334
Pertinent|5334,5343
Results|5344,5351
:|5351,5352
<EOL>|5352,5353
=|5353,5354
=|5354,5355
=|5355,5356
=|5356,5357
=|5357,5358
=|5358,5359
=|5359,5360
=|5360,5361
=|5361,5362
=|5362,5363
=|5363,5364
=|5364,5365
=|5365,5366
=|5366,5367
=|5367,5368
=|5368,5369
=|5369,5370
=|5370,5371
=|5371,5372
=|5372,5373
=|5373,5374
=|5374,5375
=|5375,5376
=|5376,5377
=|5377,5378
=|5378,5379
=|5379,5380
=|5380,5381
=|5381,5382
=|5382,5383
<EOL>|5383,5384
ADMISSION|5385,5394
LABS|5395,5399
<EOL>|5399,5400
=|5400,5401
=|5401,5402
=|5402,5403
=|5403,5404
=|5404,5405
=|5405,5406
=|5406,5407
=|5407,5408
=|5408,5409
=|5409,5410
=|5410,5411
=|5411,5412
=|5412,5413
=|5413,5414
=|5414,5415
=|5415,5416
=|5416,5417
=|5417,5418
=|5418,5419
=|5419,5420
=|5420,5421
=|5421,5422
=|5422,5423
=|5423,5424
=|5424,5425
=|5425,5426
=|5426,5427
=|5427,5428
=|5428,5429
=|5429,5430
<EOL>|5430,5431
_|5431,5432
_|5432,5433
_|5433,5434
09|5435,5437
:|5437,5438
37PM|5438,5442
BLOOD|5443,5448
WBC|5449,5452
-|5452,5453
6.0|5453,5456
RBC|5457,5460
-|5460,5461
2|5461,5462
.|5462,5463
88|5463,5465
*|5465,5466
Hgb|5467,5470
-|5470,5471
9|5471,5472
.|5472,5473
0|5473,5474
*|5474,5475
Hct|5476,5479
-|5479,5480
27|5480,5482
.|5482,5483
8|5483,5484
*|5484,5485
<EOL>|5486,5487
MCV|5487,5490
-|5490,5491
97|5491,5493
MCH|5494,5497
-|5497,5498
31.3|5498,5502
MCHC|5503,5507
-|5507,5508
32.4|5508,5512
RDW|5513,5516
-|5516,5517
15.1|5517,5521
RDWSD|5522,5527
-|5527,5528
52|5528,5530
.|5530,5531
0|5531,5532
*|5532,5533
Plt|5534,5537
_|5538,5539
_|5539,5540
_|5540,5541
<EOL>|5541,5542
_|5542,5543
_|5543,5544
_|5544,5545
09|5546,5548
:|5548,5549
37PM|5549,5553
BLOOD|5554,5559
Neuts|5560,5565
-|5565,5566
75|5566,5568
.|5568,5569
2|5569,5570
*|5570,5571
Lymphs|5572,5578
-|5578,5579
17|5579,5581
.|5581,5582
6|5582,5583
*|5583,5584
Monos|5585,5590
-|5590,5591
4|5591,5592
.|5592,5593
4|5593,5594
*|5594,5595
<EOL>|5596,5597
Eos|5597,5600
-|5600,5601
1.8|5601,5604
Baso|5605,5609
-|5609,5610
0.3|5610,5613
Im|5614,5616
_|5617,5618
_|5618,5619
_|5619,5620
AbsNeut|5621,5628
-|5628,5629
4|5629,5630
.|5630,5631
49|5631,5633
AbsLymp|5634,5641
-|5641,5642
1|5642,5643
.|5643,5644
05|5644,5646
*|5646,5647
<EOL>|5648,5649
AbsMono|5649,5656
-|5656,5657
0|5657,5658
.|5658,5659
26|5659,5661
AbsEos|5662,5668
-|5668,5669
0|5669,5670
.|5670,5671
11|5671,5673
AbsBaso|5674,5681
-|5681,5682
0|5682,5683
.|5683,5684
02|5684,5686
<EOL>|5686,5687
_|5687,5688
_|5688,5689
_|5689,5690
06|5691,5693
:|5693,5694
40AM|5694,5698
BLOOD|5699,5704
_|5705,5706
_|5706,5707
_|5707,5708
PTT|5709,5712
-|5712,5713
25.9|5713,5717
_|5718,5719
_|5719,5720
_|5720,5721
<EOL>|5721,5722
_|5722,5723
_|5723,5724
_|5724,5725
09|5726,5728
:|5728,5729
37PM|5729,5733
BLOOD|5734,5739
Glucose|5740,5747
-|5747,5748
189|5748,5751
*|5751,5752
UreaN|5753,5758
-|5758,5759
38|5759,5761
*|5761,5762
Creat|5763,5768
-|5768,5769
2|5769,5770
.|5770,5771
4|5771,5772
*|5772,5773
Na|5774,5776
-|5776,5777
142|5777,5780
<EOL>|5781,5782
K|5782,5783
-|5783,5784
4.8|5784,5787
Cl|5788,5790
-|5790,5791
105|5791,5794
HCO3|5795,5799
-|5799,5800
20|5800,5802
*|5802,5803
AnGap|5804,5809
-|5809,5810
17|5810,5812
<EOL>|5812,5813
_|5813,5814
_|5814,5815
_|5815,5816
09|5817,5819
:|5819,5820
37PM|5820,5824
BLOOD|5825,5830
proBNP|5831,5837
-|5837,5838
4512|5838,5842
*|5842,5843
<EOL>|5843,5844
_|5844,5845
_|5845,5846
_|5846,5847
09|5848,5850
:|5850,5851
37PM|5851,5855
BLOOD|5856,5861
cTropnT|5862,5869
-|5869,5870
<|5870,5871
0|5871,5872
.|5872,5873
01|5873,5875
<EOL>|5875,5876
_|5876,5877
_|5877,5878
_|5878,5879
06|5880,5882
:|5882,5883
40AM|5883,5887
BLOOD|5888,5893
CK|5894,5896
-|5896,5897
MB|5897,5899
-|5899,5900
6|5900,5901
cTropnT|5902,5909
-|5909,5910
0|5910,5911
.|5911,5912
05|5912,5914
*|5914,5915
<EOL>|5915,5916
_|5916,5917
_|5917,5918
_|5918,5919
02|5920,5922
:|5922,5923
01PM|5923,5927
BLOOD|5928,5933
CK|5934,5936
-|5936,5937
MB|5937,5939
-|5939,5940
5|5940,5941
cTropnT|5942,5949
-|5949,5950
0|5950,5951
.|5951,5952
04|5952,5954
*|5954,5955
<EOL>|5955,5956
_|5956,5957
_|5957,5958
_|5958,5959
09|5960,5962
:|5962,5963
37PM|5963,5967
BLOOD|5968,5973
Calcium|5974,5981
-|5981,5982
9.4|5982,5985
Phos|5986,5990
-|5990,5991
4.1|5991,5994
Mg|5995,5997
-|5997,5998
2.3|5998,6001
<EOL>|6001,6002
_|6002,6003
_|6003,6004
_|6004,6005
09|6006,6008
:|6008,6009
41PM|6009,6013
BLOOD|6014,6019
_|6020,6021
_|6021,6022
_|6022,6023
pO2|6024,6027
-|6027,6028
30|6028,6030
*|6030,6031
pCO2|6032,6036
-|6036,6037
40|6037,6039
pH|6040,6042
-|6042,6043
7|6043,6044
.|6044,6045
33|6045,6047
*|6047,6048
<EOL>|6049,6050
calTCO2|6050,6057
-|6057,6058
22|6058,6060
Base|6061,6065
XS|6066,6068
-|6068,6069
-|6069,6070
5|6070,6071
<EOL>|6071,6072
<EOL>|6073,6074
=|6074,6075
=|6075,6076
=|6076,6077
=|6077,6078
=|6078,6079
=|6079,6080
=|6080,6081
=|6081,6082
=|6082,6083
=|6083,6084
=|6084,6085
=|6085,6086
=|6086,6087
=|6087,6088
=|6088,6089
=|6089,6090
=|6090,6091
=|6091,6092
=|6092,6093
=|6093,6094
=|6094,6095
=|6095,6096
=|6096,6097
=|6097,6098
=|6098,6099
=|6099,6100
=|6100,6101
=|6101,6102
=|6102,6103
=|6103,6104
<EOL>|6104,6105
IMAGING|6106,6113
<EOL>|6113,6114
=|6114,6115
=|6115,6116
=|6116,6117
=|6117,6118
=|6118,6119
=|6119,6120
=|6120,6121
=|6121,6122
=|6122,6123
=|6123,6124
=|6124,6125
=|6125,6126
=|6126,6127
=|6127,6128
=|6128,6129
=|6129,6130
=|6130,6131
=|6131,6132
=|6132,6133
=|6133,6134
=|6134,6135
=|6135,6136
=|6136,6137
=|6137,6138
=|6138,6139
=|6139,6140
=|6140,6141
=|6141,6142
=|6142,6143
=|6143,6144
<EOL>|6144,6145
TTE|6145,6148
_|6149,6150
_|6150,6151
_|6151,6152
:|6152,6153
The|6154,6157
left|6158,6162
atrial|6163,6169
volume|6170,6176
index|6177,6182
is|6183,6185
mildly|6186,6192
increased|6193,6202
.|6202,6203
<EOL>|6204,6205
The|6205,6208
estimated|6209,6218
right|6219,6224
atrial|6225,6231
pressure|6232,6240
is|6241,6243
_|6244,6245
_|6245,6246
_|6246,6247
mmHg|6248,6252
.|6252,6253
Left|6254,6258
<EOL>|6259,6260
ventricular|6260,6271
wall|6272,6276
thicknesses|6277,6288
and|6289,6292
cavity|6293,6299
size|6300,6304
are|6305,6308
normal|6309,6315
.|6315,6316
There|6317,6322
<EOL>|6323,6324
is|6324,6326
mild|6327,6331
regional|6332,6340
left|6341,6345
ventricular|6346,6357
systolic|6358,6366
dysfunction|6367,6378
with|6379,6383
<EOL>|6384,6385
basal|6385,6390
inferoseptal|6391,6403
,|6403,6404
inferior|6405,6413
,|6413,6414
inferolateral|6415,6428
as|6429,6431
well|6432,6436
as|6437,6439
mid|6440,6443
<EOL>|6444,6445
inferior|6445,6453
/|6453,6454
inferoseptal|6454,6466
wall|6467,6471
motion|6472,6478
abnormalities|6479,6492
.|6492,6493
Doppler|6494,6501
<EOL>|6502,6503
parameters|6503,6513
are|6514,6517
most|6518,6522
consistent|6523,6533
with|6534,6538
Grade|6539,6544
II|6545,6547
(|6548,6549
moderate|6549,6557
)|6557,6558
left|6559,6563
<EOL>|6564,6565
ventricular|6565,6576
diastolic|6577,6586
dysfunction|6587,6598
.|6598,6599
Right|6600,6605
ventricular|6606,6617
chamber|6618,6625
<EOL>|6626,6627
size|6627,6631
and|6632,6635
free|6636,6640
wall|6641,6645
motion|6646,6652
are|6653,6656
normal|6657,6663
.|6663,6664
The|6665,6668
diameters|6669,6678
of|6679,6681
aorta|6682,6687
at|6688,6690
<EOL>|6691,6692
the|6692,6695
sinus|6696,6701
,|6701,6702
ascending|6703,6712
and|6713,6716
arch|6717,6721
levels|6722,6728
are|6729,6732
normal|6733,6739
.|6739,6740
The|6741,6744
aortic|6745,6751
<EOL>|6752,6753
valve|6753,6758
leaflets|6759,6767
(|6768,6769
3|6769,6770
)|6770,6771
are|6772,6775
mildly|6776,6782
thickened|6783,6792
but|6793,6796
aortic|6797,6803
stenosis|6804,6812
is|6813,6815
<EOL>|6816,6817
not|6817,6820
present|6821,6828
.|6828,6829
There|6830,6835
is|6836,6838
no|6839,6841
aortic|6842,6848
valve|6849,6854
stenosis|6855,6863
.|6863,6864
Trace|6865,6870
aortic|6871,6877
<EOL>|6878,6879
regurgitation|6879,6892
is|6893,6895
seen|6896,6900
.|6900,6901
The|6902,6905
mitral|6906,6912
valve|6913,6918
leaflets|6919,6927
are|6928,6931
moderately|6932,6942
<EOL>|6943,6944
thickened|6944,6953
.|6953,6954
Mild|6955,6959
(|6960,6961
1|6961,6962
+|6962,6963
)|6963,6964
mitral|6965,6971
regurgitation|6972,6985
is|6986,6988
seen|6989,6993
.|6993,6994
The|6995,6998
tricuspid|6999,7008
<EOL>|7009,7010
valve|7010,7015
leaflets|7016,7024
are|7025,7028
mildly|7029,7035
thickened|7036,7045
.|7045,7046
There|7047,7052
is|7053,7055
mild|7056,7060
pulmonary|7061,7070
<EOL>|7071,7072
artery|7072,7078
systolic|7079,7087
hypertension|7088,7100
.|7100,7101
There|7102,7107
is|7108,7110
no|7111,7113
pericardial|7114,7125
effusion|7126,7134
.|7134,7135
<EOL>|7136,7137
<EOL>|7137,7138
IMPRESSION|7139,7149
:|7149,7150
1|7153,7154
)|7154,7155
Mild|7156,7160
regional|7161,7169
LV|7170,7172
systolic|7173,7181
dysfunction|7182,7193
c|7194,7195
/|7195,7196
w|7196,7197
<EOL>|7198,7199
prior|7199,7204
myocardial|7205,7215
infarction|7216,7226
in|7227,7229
the|7230,7233
RCA|7234,7237
territory|7238,7247
.|7247,7248
2|7251,7252
)|7252,7253
Grade|7254,7259
II|7260,7262
<EOL>|7263,7264
LV|7264,7266
diastolic|7267,7276
dysfunction|7277,7288
.|7288,7289
<EOL>|7289,7290
Compared|7291,7299
with|7300,7304
the|7305,7308
prior|7309,7314
study|7315,7320
(|7321,7322
images|7322,7328
reviewed|7329,7337
)|7337,7338
of|7339,7341
_|7342,7343
_|7343,7344
_|7344,7345
,|7345,7346
LV|7347,7349
<EOL>|7350,7351
sytolic|7351,7358
function|7359,7367
appears|7368,7375
mildly|7376,7382
less|7383,7387
vigorous|7388,7396
.|7396,7397
Regional|7398,7406
wall|7407,7411
<EOL>|7412,7413
motion|7413,7419
abnormalities|7420,7433
encompassess|7434,7446
slightly|7447,7455
greater|7456,7463
territory|7464,7473
.|7473,7474
<EOL>|7476,7477
<EOL>|7477,7478
CXR|7478,7481
PA|7482,7484
&|7485,7486
LAT|7487,7490
_|7491,7492
_|7492,7493
_|7493,7494
:|7494,7495
No|7496,7498
focal|7499,7504
consolidation|7505,7518
or|7519,7521
pulmonary|7522,7531
<EOL>|7532,7533
edema|7533,7538
.|7538,7539
<EOL>|7539,7540
<EOL>|7540,7541
BILATERAL|7541,7550
LOWER|7551,7556
EXTREMITY|7557,7566
DOPPLER|7567,7574
ULTRASOUND|7575,7585
_|7586,7587
_|7587,7588
_|7588,7589
:|7589,7590
<EOL>|7593,7594
1.|7594,7596
Nonocclusive|7597,7609
thrombosis|7610,7620
of|7621,7623
one|7624,7627
of|7628,7630
the|7631,7634
paired|7635,7641
posterior|7642,7651
tibial|7652,7658
<EOL>|7659,7660
veins|7660,7665
in|7666,7668
the|7669,7672
bilateral|7673,7682
lower|7683,7688
extremities|7689,7700
which|7701,7706
appears|7707,7714
grossly|7715,7722
<EOL>|7723,7724
unchanged|7724,7733
compared|7734,7742
to|7743,7745
bilateral|7746,7755
lower|7756,7761
extremity|7762,7771
ultrasound|7772,7782
_|7783,7784
_|7784,7785
_|7785,7786
.|7786,7787
No|7789,7791
new|7792,7795
deep|7796,7800
venous|7801,7807
thrombosis|7808,7818
in|7819,7821
either|7822,7828
<EOL>|7829,7830
extremity|7830,7839
.|7839,7840
<EOL>|7841,7842
2.|7842,7844
Right|7845,7850
_|7851,7852
_|7852,7853
_|7853,7854
cyst|7855,7859
measuring|7860,7869
up|7870,7872
to|7873,7875
1.8|7876,7879
cm|7880,7882
across|7883,7889
maximal|7890,7897
<EOL>|7898,7899
diameter|7899,7907
is|7908,7910
<EOL>|7911,7912
unchanged|7912,7921
in|7922,7924
size|7925,7929
compared|7930,7938
to|7939,7941
_|7942,7943
_|7943,7944
_|7944,7945
.|7945,7946
<EOL>|7947,7948
<EOL>|7950,7951
=|7951,7952
=|7952,7953
=|7953,7954
=|7954,7955
=|7955,7956
=|7956,7957
=|7957,7958
=|7958,7959
=|7959,7960
=|7960,7961
=|7961,7962
=|7962,7963
=|7963,7964
=|7964,7965
=|7965,7966
=|7966,7967
=|7967,7968
=|7968,7969
=|7969,7970
=|7970,7971
=|7971,7972
=|7972,7973
=|7973,7974
=|7974,7975
=|7975,7976
=|7976,7977
=|7977,7978
=|7978,7979
=|7979,7980
=|7980,7981
<EOL>|7981,7982
MICROBIOLOGY|7983,7995
<EOL>|7995,7996
=|7996,7997
=|7997,7998
=|7998,7999
=|7999,8000
=|8000,8001
=|8001,8002
=|8002,8003
=|8003,8004
=|8004,8005
=|8005,8006
=|8006,8007
=|8007,8008
=|8008,8009
=|8009,8010
=|8010,8011
=|8011,8012
=|8012,8013
=|8013,8014
=|8014,8015
=|8015,8016
=|8016,8017
=|8017,8018
=|8018,8019
=|8019,8020
=|8020,8021
=|8021,8022
=|8022,8023
=|8023,8024
=|8024,8025
=|8025,8026
<EOL>|8026,8027
URINE|8028,8033
CULTURE|8034,8041
_|8042,8043
_|8043,8044
_|8044,8045
:|8045,8046
ENTEROCOCCUS|8047,8059
SP|8060,8062
.|8062,8063
.|8063,8064
>|8068,8069
100,000|8069,8076
CFU|8077,8080
/|8080,8081
mL|8081,8083
.|8083,8084
<EOL>|8084,8085
BLOOD|8086,8091
CULTURE|8092,8099
_|8100,8101
_|8101,8102
_|8102,8103
:|8103,8104
Blood|8105,8110
Culture|8111,8118
:|8118,8119
PENDING|8120,8127
<EOL>|8128,8129
BLOOD|8130,8135
CULTURE|8136,8143
_|8144,8145
_|8145,8146
_|8146,8147
:|8147,8148
Blood|8149,8154
Culture|8155,8162
:|8162,8163
PENDING|8164,8171
<EOL>|8172,8173
<EOL>|8173,8174
=|8174,8175
=|8175,8176
=|8176,8177
=|8177,8178
=|8178,8179
=|8179,8180
=|8180,8181
=|8181,8182
=|8182,8183
=|8183,8184
=|8184,8185
=|8185,8186
=|8186,8187
=|8187,8188
=|8188,8189
=|8189,8190
=|8190,8191
=|8191,8192
=|8192,8193
=|8193,8194
=|8194,8195
=|8195,8196
=|8196,8197
=|8197,8198
=|8198,8199
=|8199,8200
=|8200,8201
=|8201,8202
=|8202,8203
=|8203,8204
<EOL>|8204,8205
DISCHARGE|8206,8215
LABS|8216,8220
<EOL>|8220,8221
=|8221,8222
=|8222,8223
=|8223,8224
=|8224,8225
=|8225,8226
=|8226,8227
=|8227,8228
=|8228,8229
=|8229,8230
=|8230,8231
=|8231,8232
=|8232,8233
=|8233,8234
=|8234,8235
=|8235,8236
=|8236,8237
=|8237,8238
=|8238,8239
=|8239,8240
=|8240,8241
=|8241,8242
=|8242,8243
=|8243,8244
=|8244,8245
=|8245,8246
=|8246,8247
=|8247,8248
=|8248,8249
=|8249,8250
=|8250,8251
<EOL>|8251,8252
_|8252,8253
_|8253,8254
_|8254,8255
05|8256,8258
:|8258,8259
45AM|8259,8263
BLOOD|8264,8269
WBC|8270,8273
-|8273,8274
5.1|8274,8277
RBC|8278,8281
-|8281,8282
2|8282,8283
.|8283,8284
57|8284,8286
*|8286,8287
Hgb|8288,8291
-|8291,8292
7|8292,8293
.|8293,8294
9|8294,8295
*|8295,8296
Hct|8297,8300
-|8300,8301
24|8301,8303
.|8303,8304
5|8304,8305
*|8305,8306
<EOL>|8307,8308
MCV|8308,8311
-|8311,8312
95|8312,8314
MCH|8315,8318
-|8318,8319
30.7|8319,8323
MCHC|8324,8328
-|8328,8329
32.2|8329,8333
RDW|8334,8337
-|8337,8338
15.0|8338,8342
RDWSD|8343,8348
-|8348,8349
51|8349,8351
.|8351,8352
8|8352,8353
*|8353,8354
Plt|8355,8358
_|8359,8360
_|8360,8361
_|8361,8362
<EOL>|8362,8363
_|8363,8364
_|8364,8365
_|8365,8366
05|8367,8369
:|8369,8370
45AM|8370,8374
BLOOD|8375,8380
Glucose|8381,8388
-|8388,8389
144|8389,8392
*|8392,8393
UreaN|8394,8399
-|8399,8400
49|8400,8402
*|8402,8403
Creat|8404,8409
-|8409,8410
2|8410,8411
.|8411,8412
6|8412,8413
*|8413,8414
Na|8415,8417
-|8417,8418
147|8418,8421
<EOL>|8422,8423
K|8423,8424
-|8424,8425
4.0|8425,8428
Cl|8429,8431
-|8431,8432
105|8432,8435
HCO3|8436,8440
-|8440,8441
24|8441,8443
AnGap|8444,8449
-|8449,8450
_|8450,8451
_|8451,8452
_|8452,8453
yo|8454,8456
F|8457,8458
PMH|8460,8463
CAD|8464,8467
c|8468,8469
/|8469,8470
b|8470,8471
ischemic|8472,8480
MR|8481,8483
_|8484,8485
_|8485,8486
_|8486,8487
DES|8488,8491
to|8492,8494
_|8495,8496
_|8496,8497
_|8497,8498
_|8499,8500
_|8500,8501
_|8501,8502
,|8502,8503
TTE|8504,8507
_|8508,8509
_|8509,8510
_|8510,8511
<EOL>|8512,8513
with|8513,8517
mild|8518,8522
regional|8523,8531
LV|8532,8534
systolic|8535,8543
dysfunction|8544,8555
)|8555,8556
,|8556,8557
HFpEF|8558,8563
(|8564,8565
LVEF|8565,8569
50|8570,8572
%|8572,8573
<EOL>|8574,8575
_|8575,8576
_|8576,8577
_|8577,8578
,|8578,8579
PAD|8580,8583
,|8583,8584
CKD|8585,8588
(|8589,8590
stage|8590,8595
IV|8596,8598
)|8598,8599
,|8599,8600
prior|8601,8606
DVT|8607,8610
c|8611,8612
/|8612,8613
b|8613,8614
severe|8615,8621
UGIV|8622,8626
on|8627,8629
AC|8630,8632
,|8632,8633
<EOL>|8634,8635
T2DM|8635,8639
presents|8640,8648
with|8649,8653
subacute|8654,8662
SOB|8663,8666
,|8666,8667
weight|8668,8674
gain|8675,8679
,|8679,8680
c|8681,8682
/|8682,8683
f|8683,8684
acute|8685,8690
heart|8691,8696
<EOL>|8697,8698
failure|8698,8705
exacerbation|8706,8718
.|8718,8719
She|8721,8724
underwent|8725,8734
diuresis|8735,8743
with|8744,8748
IV|8749,8751
Lasix|8752,8757
80|8758,8760
<EOL>|8761,8762
mg|8762,8764
,|8764,8765
120mg|8766,8771
IV|8772,8774
x2|8775,8777
with|8778,8782
rapid|8783,8788
improvement|8789,8800
in|8801,8803
subjective|8804,8814
dyspnea|8815,8822
.|8822,8823
<EOL>|8825,8826
_|8826,8827
_|8827,8828
_|8828,8829
showed|8830,8836
no|8837,8839
acute|8840,8845
DVT|8846,8849
,|8849,8850
CXR|8851,8854
without|8855,8862
sign|8863,8867
of|8868,8870
consolidation|8871,8884
.|8884,8885
<EOL>|8887,8888
Given|8888,8893
her|8894,8897
improvement|8898,8909
in|8910,8912
dyspnea|8913,8920
,|8920,8921
no|8922,8924
supplemental|8925,8937
O2|8938,8940
<EOL>|8941,8942
requirement|8942,8953
,|8953,8954
the|8955,8958
patient|8959,8966
was|8967,8970
discharged|8971,8981
w|8982,8983
/|8983,8984
o|8984,8985
medication|8986,8996
changes|8997,9004
.|9004,9005
<EOL>|9005,9006
<EOL>|9006,9007
#|9007,9008
Shortness|9009,9018
of|9019,9021
breath|9022,9028
<EOL>|9028,9029
#|9029,9030
Hypoxia|9031,9038
<EOL>|9038,9039
#|9039,9040
acute|9041,9046
exacerbation|9047,9059
of|9060,9062
chronic|9063,9070
diastolic|9071,9080
heart|9081,9086
failure|9087,9094
with|9095,9099
<EOL>|9100,9101
preserved|9101,9110
LVEF|9111,9115
(|9116,9117
50|9117,9119
%|9119,9120
)|9120,9121
<EOL>|9121,9122
Dry|9122,9125
weight|9126,9132
per|9133,9136
pt|9137,9139
154|9140,9143
lbs|9144,9147
.|9147,9148
Admission|9150,9159
weight|9160,9166
above|9167,9172
baseline|9173,9181
,|9181,9182
BNP|9183,9186
<EOL>|9187,9188
elevated|9188,9196
.|9196,9197
Regarding|9199,9208
trigger|9209,9216
,|9216,9217
suspect|9218,9225
dietary|9226,9233
vs|9234,9236
uncontrolled|9237,9249
<EOL>|9250,9251
BP|9251,9253
.|9253,9254
No|9255,9257
EKG|9258,9261
changes|9262,9269
for|9270,9273
ACS|9274,9277
,|9277,9278
trop|9279,9283
negative|9284,9292
,|9292,9293
repeat|9294,9300
TTE|9301,9304
showed|9305,9311
<EOL>|9312,9313
mild|9313,9317
regional|9318,9326
LV|9327,9329
systolic|9330,9338
dysfunction|9339,9350
c|9351,9352
/|9352,9353
w|9353,9354
prior|9355,9360
myocardial|9361,9371
<EOL>|9372,9373
infarction|9373,9383
in|9384,9386
the|9387,9390
RCA|9391,9394
territory|9395,9404
,|9404,9405
as|9406,9408
well|9409,9413
as|9414,9416
Grade|9417,9422
II|9423,9425
LV|9426,9428
<EOL>|9429,9430
diastolic|9430,9439
dysfunction|9440,9451
and|9452,9455
similar|9456,9463
to|9464,9466
prior|9467,9472
_|9473,9474
_|9474,9475
_|9475,9476
TTE|9477,9480
.|9480,9481
Doubt|9482,9487
PNA|9488,9491
<EOL>|9492,9493
given|9493,9498
CXR|9499,9502
and|9503,9506
lack|9507,9511
of|9512,9514
cough|9515,9520
/|9520,9521
fever|9521,9526
,|9526,9527
doubt|9528,9533
PE|9534,9536
given|9537,9542
low|9543,9546
Wells|9547,9552
'|9552,9553
<EOL>|9554,9555
score|9555,9560
1.5|9561,9564
,|9564,9565
and|9566,9569
stable|9570,9576
repeat|9577,9583
_|9584,9585
_|9585,9586
_|9586,9587
.|9587,9588
Underwent|9589,9598
diuresis|9599,9607
with|9608,9612
IV|9613,9615
<EOL>|9616,9617
Lasix|9617,9622
80|9623,9625
mg|9626,9628
,|9628,9629
120mg|9630,9635
IV|9636,9638
x2|9639,9641
with|9642,9646
rapid|9647,9652
improvement|9653,9664
in|9665,9667
subjective|9668,9678
<EOL>|9679,9680
dyspnea|9680,9687
.|9687,9688
Resumed|9690,9697
home|9698,9702
torsemide|9703,9712
40mg|9713,9717
,|9717,9718
nifedipine|9719,9729
60mg|9730,9734
BID|9735,9738
and|9739,9742
<EOL>|9743,9744
carvedilol|9744,9754
25mg|9755,9759
BID|9760,9763
.|9763,9764
Was|9766,9769
stable|9770,9776
on|9777,9779
RA|9780,9782
prior|9783,9788
to|9789,9791
discharge|9792,9801
.|9801,9802
<EOL>|9802,9803
<EOL>|9803,9804
#|9804,9805
Hypertension|9806,9818
-|9819,9820
Patient|9821,9828
missed|9829,9835
her|9836,9839
antiHTN|9840,9847
medications|9848,9859
earlier|9860,9867
<EOL>|9868,9869
day|9869,9872
of|9873,9875
admission|9876,9885
.|9885,9886
Continued|9887,9896
home|9897,9901
carvedilol|9902,9912
25mg|9913,9917
BID|9918,9921
and|9922,9925
<EOL>|9926,9927
nifedipine|9927,9937
60mg|9938,9942
BID|9943,9946
with|9947,9951
holding|9952,9959
parameters|9960,9970
.|9970,9971
Appears|9972,9979
that|9980,9984
a|9985,9986
<EOL>|9987,9988
trial|9988,9993
of|9994,9996
_|9997,9998
_|9998,9999
_|9999,10000
or|10001,10003
spironolactone|10004,10018
would|10019,10024
be|10025,10027
limited|10028,10035
by|10036,10038
<EOL>|10039,10040
hyperkalemia|10040,10052
,|10052,10053
so|10054,10056
this|10057,10061
was|10062,10065
deferred|10066,10074
.|10074,10075
<EOL>|10075,10076
<EOL>|10081,10082
#|10082,10083
Urinary|10084,10091
frequency|10092,10101
/|10101,10102
urge|10102,10106
incontinence|10107,10119
:|10119,10120
occurred|10121,10129
in|10130,10132
setting|10133,10140
of|10141,10143
<EOL>|10144,10145
diuresis|10145,10153
,|10153,10154
however|10155,10162
UCx|10163,10166
ordered|10167,10174
in|10175,10177
ED|10178,10180
did|10181,10184
grow|10185,10189
enterococci|10190,10201
,|10201,10202
likely|10203,10209
<EOL>|10210,10211
colonization|10211,10223
.|10223,10224
If|10225,10227
symptoms|10228,10236
persists|10237,10245
would|10246,10251
revaluate|10252,10261
/|10261,10262
treat|10262,10267
.|10267,10268
<EOL>|10268,10269
<EOL>|10278,10279
CHRONIC|10279,10286
STABLE|10287,10293
ISSUES|10294,10300
<EOL>|10300,10301
<EOL>|10301,10302
#|10302,10303
Normocytic|10304,10314
anemia|10315,10321
(|10322,10323
recent|10323,10329
baseline|10330,10338
Hb|10339,10341
9.4|10342,10345
_|10346,10347
_|10347,10348
_|10348,10349
-|10350,10351
Hb|10352,10354
was|10355,10358
at|10359,10361
<EOL>|10362,10363
baseline|10363,10371
,|10371,10372
no|10373,10375
signs|10376,10381
of|10382,10384
active|10385,10391
bleeding|10392,10400
.|10400,10401
Likely|10403,10409
multifactorial|10410,10424
,|10424,10425
<EOL>|10426,10427
anemia|10427,10433
of|10434,10436
chronic|10437,10444
disease|10445,10452
as|10453,10455
well|10456,10460
as|10461,10463
decreased|10464,10473
erythropoiten|10474,10487
<EOL>|10488,10489
production|10489,10499
iso|10500,10503
CKD|10504,10507
.|10507,10508
<EOL>|10508,10509
<EOL>|10510,10511
#|10511,10512
Non|10513,10516
anion|10517,10522
gap|10523,10526
metabolic|10527,10536
acidosis|10537,10545
-|10546,10547
Patient|10548,10555
has|10556,10559
intermittently|10560,10574
<EOL>|10575,10576
had|10576,10579
a|10580,10581
NAGMA|10582,10587
in|10588,10590
the|10591,10594
past|10595,10599
.|10599,10600
No|10602,10604
recent|10605,10611
diarrhea|10612,10620
.|10620,10621
_|10623,10624
_|10624,10625
_|10625,10626
suspect|10627,10634
Type|10635,10639
<EOL>|10640,10641
IV|10641,10643
RTA|10644,10647
given|10648,10653
advanced|10654,10662
age|10663,10666
and|10667,10670
history|10671,10678
of|10679,10681
T2DM|10682,10686
(|10687,10688
both|10688,10692
of|10693,10695
which|10696,10701
can|10702,10705
<EOL>|10706,10707
cause|10707,10712
hyporeninemia|10713,10726
)|10726,10727
.|10727,10728
<EOL>|10728,10729
<EOL>|10729,10730
#|10730,10731
Stage|10732,10737
IV|10738,10740
Chronic|10741,10748
Kidney|10749,10755
Disease|10756,10763
(|10764,10765
baseline|10765,10773
Cr|10774,10776
2.3|10777,10780
-|10780,10781
2.8|10781,10784
)|10784,10785
-|10786,10787
CKD|10788,10791
<EOL>|10792,10793
iso|10793,10796
HTN|10797,10800
and|10801,10804
T2DM|10805,10809
,|10809,10810
Cr|10811,10813
is|10814,10816
currently|10817,10826
at|10827,10829
baseline|10830,10838
.|10838,10839
Low|10840,10843
K|10844,10845
/|10845,10846
Phos|10846,10850
/|10850,10851
Na|10851,10853
<EOL>|10854,10855
diet|10855,10859
.|10859,10860
Continued|10861,10870
home|10871,10875
calcitriol|10876,10886
,|10886,10887
avoided|10888,10895
nephrotoxins|10896,10908
and|10909,10912
<EOL>|10913,10914
renally|10914,10921
dosed|10922,10927
all|10928,10931
medications|10932,10943
.|10943,10944
<EOL>|10944,10945
<EOL>|10945,10946
#|10946,10947
Coronary|10948,10956
artery|10957,10963
disease|10964,10971
_|10972,10973
_|10973,10974
_|10974,10975
DES|10976,10979
to|10980,10982
LCX|10983,10986
_|10987,10988
_|10988,10989
_|10989,10990
:|10990,10991
troponins|10992,11001
were|11002,11006
<EOL>|11007,11008
trended|11008,11015
from|11016,11020
<|11021,11022
0.01|11023,11027
to|11028,11030
0.05|11031,11035
to|11036,11038
0.04|11039,11043
then|11044,11048
stopped|11049,11056
.|11056,11057
CK|11058,11060
-|11060,11061
MB|11061,11063
was|11064,11067
<EOL>|11068,11069
flat|11069,11073
.|11073,11074
Patient|11076,11083
deneied|11084,11091
any|11092,11095
chest|11096,11101
pain|11102,11106
.|11106,11107
A|11108,11109
TTE|11110,11113
showed|11114,11120
mild|11121,11125
<EOL>|11126,11127
regional|11127,11135
LV|11136,11138
systolic|11139,11147
dysfunction|11148,11159
c|11160,11161
/|11161,11162
w|11162,11163
prior|11164,11169
myocardial|11170,11180
infarction|11181,11191
<EOL>|11192,11193
in|11193,11195
the|11196,11199
RCA|11200,11203
territory|11204,11213
and|11214,11217
similar|11218,11225
to|11226,11228
prior|11229,11234
_|11235,11236
_|11236,11237
_|11237,11238
TTE|11239,11242
.|11242,11243
Continued|11244,11253
<EOL>|11254,11255
home|11255,11259
aspirin|11260,11267
81mg|11268,11272
qd|11273,11275
,|11275,11276
home|11277,11281
carvedilol|11282,11292
25mg|11293,11297
BID|11298,11301
with|11302,11306
holding|11307,11314
<EOL>|11315,11316
parameters|11316,11326
,|11326,11327
home|11328,11332
atorvastatin|11333,11345
80mg|11346,11350
qHS|11351,11354
.|11354,11355
<EOL>|11355,11356
<EOL>|11357,11358
#|11358,11359
Type|11360,11364
II|11365,11367
Diabetes|11368,11376
Mellitus|11377,11385
(|11386,11387
last|11387,11391
HbA1C|11392,11397
6.4|11398,11401
%|11401,11402
_|11403,11404
_|11404,11405
_|11405,11406
-|11407,11408
Under|11409,11414
<EOL>|11415,11416
excellent|11416,11425
control|11426,11433
,|11433,11434
most|11435,11439
recently|11440,11448
in|11449,11451
the|11452,11455
pre-diabetic|11456,11468
range|11469,11474
.|11474,11475
<EOL>|11475,11476
-|11476,11477
Continue|11478,11486
home|11487,11491
70|11492,11494
/|11494,11495
30|11495,11497
sliding|11498,11505
scale|11506,11511
(|11512,11513
_|11513,11514
_|11514,11515
_|11515,11516
t|11516,11517
dinner|11518,11524
if|11525,11527
<EOL>|11528,11529
blood|11529,11534
sugar|11535,11540
over|11541,11545
130|11546,11549
,|11549,11550
10|11551,11553
units|11554,11559
90|11560,11562
-|11562,11563
130|11563,11566
,|11566,11567
none|11568,11572
if|11573,11575
blood|11576,11581
sugar|11582,11587
under|11588,11593
<EOL>|11594,11595
90|11595,11597
)|11597,11598
<EOL>|11599,11600
<EOL>|11600,11601
#|11601,11602
Dyslipidemia|11603,11615
:|11615,11616
continued|11617,11626
home|11627,11631
atorvastatin|11632,11644
<EOL>|11644,11645
<EOL>|11645,11646
#|11646,11647
Insomnia|11648,11656
:|11656,11657
continued|11658,11667
home|11668,11672
gabapentin|11673,11683
<EOL>|11683,11684
<EOL>|11684,11685
#|11685,11686
Gout|11687,11691
:|11691,11692
continued|11693,11702
home|11703,11707
allopurinol|11708,11719
<EOL>|11719,11720
<EOL>|11721,11722
=|11722,11723
=|11723,11724
=|11724,11725
=|11725,11726
=|11726,11727
=|11727,11728
=|11728,11729
=|11729,11730
=|11730,11731
=|11731,11732
=|11732,11733
=|11733,11734
=|11734,11735
=|11735,11736
=|11736,11737
=|11737,11738
=|11738,11739
=|11739,11740
=|11740,11741
=|11741,11742
=|11742,11743
=|11743,11744
=|11744,11745
=|11745,11746
=|11746,11747
=|11747,11748
=|11748,11749
=|11749,11750
=|11750,11751
=|11751,11752
<EOL>|11752,11753
TRANSITIONAL|11754,11766
ISSUES|11767,11773
<EOL>|11773,11774
=|11774,11775
=|11775,11776
=|11776,11777
=|11777,11778
=|11778,11779
=|11779,11780
=|11780,11781
=|11781,11782
=|11782,11783
=|11783,11784
=|11784,11785
=|11785,11786
=|11786,11787
=|11787,11788
=|11788,11789
=|11789,11790
=|11790,11791
=|11791,11792
=|11792,11793
=|11793,11794
=|11794,11795
=|11795,11796
=|11796,11797
=|11797,11798
=|11798,11799
=|11799,11800
=|11800,11801
=|11801,11802
=|11802,11803
=|11803,11804
<EOL>|11804,11805
-|11805,11806
Discharge|11807,11816
weight|11817,11823
:|11823,11824
69.2|11825,11829
kg|11829,11831
<EOL>|11831,11832
-|11832,11833
Discharge|11834,11843
creatinine|11844,11854
:|11854,11855
2.6|11856,11859
<EOL>|11859,11860
-|11860,11861
Discharge|11862,11871
oral|11872,11876
diuretic|11877,11885
:|11885,11886
torsemide|11887,11896
40mg|11897,11901
daily|11902,11907
<EOL>|11907,11908
-|11908,11909
Transitional|11910,11922
issue|11923,11928
:|11928,11929
consider|11930,11938
outpatient|11939,11949
epo|11950,11953
with|11954,11958
renal|11959,11964
<EOL>|11965,11966
-|11966,11967
Transitional|11968,11980
issue|11981,11986
:|11986,11987
BP|11988,11990
goal|11991,11995
of|11996,11998
140|11999,12002
/|12002,12003
90|12003,12005
per|12006,12009
accord|12010,12016
or|12017,12019
even|12020,12024
<EOL>|12025,12026
130|12026,12029
/|12029,12030
80|12030,12032
per|12033,12036
ACC|12037,12040
/|12040,12041
AHA|12041,12044
_|12045,12046
_|12046,12047
_|12047,12048
guidelines|12049,12059
however|12060,12067
anticipate|12068,12078
difficulty|12079,12089
<EOL>|12090,12091
in|12091,12093
adding|12094,12100
additional|12101,12111
agents|12112,12118
iso|12119,12122
CKD|12123,12126
(|12127,12128
limits|12128,12134
use|12135,12138
of|12139,12141
clonidine|12142,12151
)|12151,12152
<EOL>|12153,12154
and|12154,12157
baseline|12158,12166
potassium|12167,12176
(|12177,12178
would|12178,12183
likely|12184,12190
limit|12191,12196
_|12197,12198
_|12198,12199
_|12199,12200
or|12201,12203
<EOL>|12204,12205
spironolactone|12205,12219
)|12219,12220
<EOL>|12221,12222
-|12222,12223
TTE|12224,12227
showed|12228,12234
prior|12235,12240
LV|12241,12243
hypokinesis|12244,12255
,|12255,12256
could|12257,12262
consider|12263,12271
MIBI|12272,12276
or|12277,12279
<EOL>|12280,12281
outpatient|12281,12291
pharmacological|12292,12307
stress|12308,12314
test|12315,12319
<EOL>|12319,12320
-|12320,12321
had|12322,12325
some|12326,12330
urinary|12331,12338
retention|12339,12348
/|12348,12349
incontinence|12349,12361
while|12362,12367
undergoing|12368,12378
IV|12379,12381
<EOL>|12382,12383
diuresis|12383,12391
would|12392,12397
assess|12398,12404
for|12405,12408
recurrent|12409,12418
symptoms|12419,12427
at|12428,12430
routine|12431,12438
<EOL>|12439,12440
outpatient|12440,12450
visits|12451,12457
<EOL>|12457,12458
<EOL>|12458,12459
#|12459,12460
CODE|12460,12464
:|12464,12465
Full|12466,12470
(|12471,12472
confirmed|12472,12481
)|12481,12482
<EOL>|12484,12485
#|12485,12486
CONTACT|12486,12493
:|12493,12494
_|12495,12496
_|12496,12497
_|12497,12498
(|12499,12500
husband|12500,12507
)|12507,12508
_|12509,12510
_|12510,12511
_|12511,12512
<EOL>|12512,12513
<EOL>|12514,12515
Medications|12515,12526
on|12527,12529
Admission|12530,12539
:|12539,12540
<EOL>|12540,12541
The|12541,12544
Preadmission|12545,12557
Medication|12558,12568
list|12569,12573
is|12574,12576
accurate|12577,12585
and|12586,12589
complete|12590,12598
.|12598,12599
<EOL>|12599,12600
1.|12600,12602
Allopurinol|12603,12614
_|12615,12616
_|12616,12617
_|12617,12618
mg|12619,12621
PO|12622,12624
EVERY|12625,12630
OTHER|12631,12636
DAY|12637,12640
<EOL>|12641,12642
2.|12642,12644
Atorvastatin|12645,12657
80|12658,12660
mg|12661,12663
PO|12664,12666
QPM|12667,12670
<EOL>|12671,12672
3.|12672,12674
Calcitriol|12675,12685
0.5|12686,12689
mcg|12690,12693
PO|12694,12696
DAILY|12697,12702
<EOL>|12703,12704
4.|12704,12706
Carvedilol|12707,12717
25|12718,12720
mg|12721,12723
PO|12724,12726
BID|12727,12730
<EOL>|12731,12732
5.|12732,12734
Gabapentin|12735,12745
100|12746,12749
mg|12750,12752
PO|12753,12755
QHS|12756,12759
<EOL>|12760,12761
6.|12761,12763
NIFEdipine|12764,12774
(|12775,12776
Extended|12776,12784
Release|12785,12792
)|12792,12793
60|12794,12796
mg|12797,12799
PO|12800,12802
BID|12803,12806
<EOL>|12807,12808
7.|12808,12810
Torsemide|12811,12820
40|12821,12823
mg|12824,12826
PO|12827,12829
DAILY|12830,12835
<EOL>|12836,12837
8.|12837,12839
Nitroglycerin|12840,12853
SL|12854,12856
0.3|12857,12860
mg|12861,12863
SL|12864,12866
Q5MIN|12867,12872
:|12872,12873
PRN|12873,12876
chest|12877,12882
pain|12883,12887
<EOL>|12888,12889
9.|12889,12891
Acetaminophen|12892,12905
325|12906,12909
-|12909,12910
650|12910,12913
mg|12914,12916
PO|12917,12919
Q6H|12920,12923
:|12923,12924
PRN|12924,12927
Pain|12928,12932
-|12933,12934
Mild|12935,12939
<EOL>|12940,12941
10.|12941,12944
Aspirin|12945,12952
81|12953,12955
mg|12956,12958
PO|12959,12961
DAILY|12962,12967
<EOL>|12968,12969
11.|12969,12972
Insulin|12973,12980
SC|12981,12983
<EOL>|12984,12985
Sliding|12991,12998
Scale|12999,13004
<EOL>|13004,13005
Insulin|13005,13012
SC|13013,13015
Sliding|13016,13023
Scale|13024,13029
using|13030,13035
70|13036,13038
/|13038,13039
30|13039,13041
Insulin|13042,13049
<EOL>|13049,13050
<EOL>|13050,13051
<EOL>|13052,13053
Discharge|13053,13062
Medications|13063,13074
:|13074,13075
<EOL>|13075,13076
1.|13076,13078
Acetaminophen|13080,13093
325|13094,13097
-|13097,13098
650|13098,13101
mg|13102,13104
PO|13105,13107
Q6H|13108,13111
:|13111,13112
PRN|13112,13115
Pain|13116,13120
-|13121,13122
Mild|13123,13127
<EOL>|13129,13130
2.|13130,13132
Allopurinol|13134,13145
_|13146,13147
_|13147,13148
_|13148,13149
mg|13150,13152
PO|13153,13155
EVERY|13156,13161
OTHER|13162,13167
DAY|13168,13171
<EOL>|13173,13174
3.|13174,13176
Aspirin|13178,13185
81|13186,13188
mg|13189,13191
PO|13192,13194
DAILY|13195,13200
<EOL>|13202,13203
4.|13203,13205
Atorvastatin|13207,13219
80|13220,13222
mg|13223,13225
PO|13226,13228
QPM|13229,13232
<EOL>|13234,13235
5.|13235,13237
Calcitriol|13239,13249
0.5|13250,13253
mcg|13254,13257
PO|13258,13260
DAILY|13261,13266
<EOL>|13268,13269
6.|13269,13271
Carvedilol|13273,13283
25|13284,13286
mg|13287,13289
PO|13290,13292
BID|13293,13296
<EOL>|13298,13299
7.|13299,13301
Gabapentin|13303,13313
100|13314,13317
mg|13318,13320
PO|13321,13323
QHS|13324,13327
<EOL>|13329,13330
8.|13330,13332
Insulin|13334,13341
SC|13342,13344
<EOL>|13345,13346
Sliding|13352,13359
Scale|13360,13365
<EOL>|13365,13366
Insulin|13366,13373
SC|13374,13376
Sliding|13377,13384
Scale|13385,13390
using|13391,13396
70|13397,13399
/|13399,13400
30|13400,13402
Insulin|13403,13410
<EOL>|13411,13412
9.|13412,13414
NIFEdipine|13416,13426
(|13427,13428
Extended|13428,13436
Release|13437,13444
)|13444,13445
60|13446,13448
mg|13449,13451
PO|13452,13454
BID|13455,13458
<EOL>|13460,13461
10.|13461,13464
Nitroglycerin|13466,13479
SL|13480,13482
0.3|13483,13486
mg|13487,13489
SL|13490,13492
Q5MIN|13493,13498
:|13498,13499
PRN|13499,13502
chest|13503,13508
pain|13509,13513
<EOL>|13515,13516
11|13516,13518
.|13518,13519
Torsemide|13521,13530
40|13531,13533
mg|13534,13536
PO|13537,13539
DAILY|13540,13545
<EOL>|13547,13548
<EOL>|13548,13549
<EOL>|13550,13551
Discharge|13551,13560
Disposition|13561,13572
:|13572,13573
<EOL>|13573,13574
Home|13574,13578
With|13579,13583
Service|13584,13591
<EOL>|13591,13592
<EOL>|13593,13594
Facility|13594,13602
:|13602,13603
<EOL>|13603,13604
_|13604,13605
_|13605,13606
_|13606,13607
<EOL>|13607,13608
<EOL>|13609,13610
Discharge|13610,13619
Diagnosis|13620,13629
:|13629,13630
<EOL>|13630,13631
PRIMARY|13631,13638
DIAGNOSIS|13639,13648
<EOL>|13648,13649
-|13649,13650
Acute|13651,13656
on|13657,13659
chronic|13660,13667
diastolic|13668,13677
congestive|13678,13688
heart|13689,13694
failure|13695,13702
<EOL>|13702,13703
<EOL>|13703,13704
SECONDARY|13704,13713
DIAGNOSES|13714,13723
<EOL>|13723,13724
-|13724,13725
Hypertension|13726,13738
<EOL>|13738,13739
-|13739,13740
History|13741,13748
of|13749,13751
prior|13752,13757
DVT|13758,13761
<EOL>|13761,13762
-|13762,13763
Anemia|13764,13770
,|13770,13771
NOS|13772,13775
<EOL>|13775,13776
-|13776,13777
Chronic|13778,13785
Kidney|13786,13792
Disease|13793,13800
stage|13801,13806
IV|13807,13809
<EOL>|13809,13810
-|13810,13811
Coronary|13812,13820
Artery|13821,13827
Disease|13828,13835
_|13836,13837
_|13837,13838
_|13838,13839
drug|13840,13844
eluting|13845,13852
stent|13853,13858
<EOL>|13858,13859
-|13859,13860
Diabetes|13861,13869
Mellitus|13870,13878
Type|13879,13883
2|13884,13885
controlled|13886,13896
<EOL>|13896,13897
<EOL>|13897,13898
<EOL>|13899,13900
Discharge|13900,13909
Condition|13910,13919
:|13919,13920
<EOL>|13920,13921
Mental|13921,13927
Status|13928,13934
:|13934,13935
Clear|13936,13941
and|13942,13945
coherent|13946,13954
.|13954,13955
<EOL>|13955,13956
Level|13956,13961
of|13962,13964
Consciousness|13965,13978
:|13978,13979
Alert|13980,13985
and|13986,13989
interactive|13990,14001
.|14001,14002
<EOL>|14002,14003
Activity|14003,14011
Status|14012,14018
:|14018,14019
Ambulatory|14020,14030
-|14031,14032
Independent|14033,14044
.|14044,14045
<EOL>|14045,14046
<EOL>|14046,14047
<EOL>|14048,14049
Discharge|14049,14058
Instructions|14059,14071
:|14071,14072
<EOL>|14072,14073
Dear|14073,14077
_|14078,14079
_|14079,14080
_|14080,14081
,|14081,14082
<EOL>|14082,14083
<EOL>|14083,14084
You|14084,14087
were|14088,14092
admitted|14093,14101
to|14102,14104
the|14105,14108
hospital|14109,14117
with|14118,14122
shortness|14123,14132
of|14133,14135
breath|14136,14142
and|14143,14146
<EOL>|14147,14148
weight|14148,14154
gain|14155,14159
.|14159,14160
This|14162,14166
was|14167,14170
likely|14171,14177
caused|14178,14184
by|14185,14187
an|14188,14190
exacerbation|14191,14203
of|14204,14206
your|14207,14211
<EOL>|14212,14213
heart|14213,14218
failure|14219,14226
possibly|14227,14235
from|14236,14240
salty|14241,14246
foods|14247,14252
over|14253,14257
the|14258,14261
holiday|14262,14269
.|14269,14270
<EOL>|14271,14272
<EOL>|14272,14273
While|14273,14278
you|14279,14282
were|14283,14287
in|14288,14290
the|14291,14294
hospital|14295,14303
:|14303,14304
<EOL>|14304,14305
-|14305,14306
we|14307,14309
gave|14310,14314
you|14315,14318
IV|14319,14321
diuretics|14322,14331
to|14332,14334
help|14335,14339
remove|14340,14346
extra|14347,14352
fluid|14353,14358
<EOL>|14358,14359
-|14359,14360
we|14361,14363
checked|14364,14371
for|14372,14375
pneumonia|14376,14385
with|14386,14390
a|14391,14392
chest|14393,14398
x-ray|14399,14404
,|14404,14405
there|14406,14411
was|14412,14415
no|14416,14418
sign|14419,14423
<EOL>|14424,14425
of|14425,14427
a|14428,14429
pneumonia|14430,14439
<EOL>|14439,14440
-|14440,14441
we|14442,14444
checked|14445,14452
for|14453,14456
signs|14457,14462
on|14463,14465
new|14466,14469
clots|14470,14475
in|14476,14478
your|14479,14483
legs|14484,14488
,|14488,14489
there|14490,14495
was|14496,14499
no|14500,14502
<EOL>|14503,14504
new|14504,14507
clot|14508,14512
<EOL>|14512,14513
<EOL>|14513,14514
Now|14514,14517
that|14518,14522
you|14523,14526
are|14527,14530
going|14531,14536
home|14537,14541
:|14541,14542
<EOL>|14542,14543
-|14543,14544
continue|14545,14553
to|14554,14556
take|14557,14561
all|14562,14565
of|14566,14568
your|14569,14573
medications|14574,14585
as|14586,14588
prescribed|14589,14599
<EOL>|14599,14600
-|14600,14601
monitor|14602,14609
your|14610,14614
salt|14615,14619
intake|14620,14626
,|14626,14627
this|14628,14632
should|14633,14639
be|14640,14642
no|14643,14645
more|14646,14650
than|14651,14655
2|14656,14657
grams|14658,14663
<EOL>|14664,14665
every|14665,14670
day|14671,14674
,|14674,14675
ask|14676,14679
your|14680,14684
doctors|14685,14692
for|14693,14696
help|14697,14701
with|14702,14706
this|14707,14711
if|14712,14714
you|14715,14718
do|14719,14721
not|14722,14725
<EOL>|14726,14727
know|14727,14731
how|14732,14735
to|14736,14738
keep|14739,14743
track|14744,14749
of|14750,14752
your|14753,14757
salt|14758,14762
<EOL>|14762,14763
-|14763,14764
continue|14765,14773
to|14774,14776
weigh|14777,14782
yourself|14783,14791
every|14792,14797
morning|14798,14805
,|14805,14806
call|14807,14811
your|14812,14816
doctor|14817,14823
if|14824,14826
<EOL>|14827,14828
weight|14828,14834
goes|14835,14839
up|14840,14842
more|14843,14847
than|14848,14852
3|14853,14854
lbs|14855,14858
.|14858,14859
<EOL>|14859,14860
-|14860,14861
follow|14862,14868
-|14868,14869
up|14869,14871
with|14872,14876
your|14877,14881
primary|14882,14889
care|14890,14894
doctor|14895,14901
regarding|14902,14911
your|14912,14916
blood|14917,14922
<EOL>|14923,14924
pressure|14924,14932
and|14933,14936
blood|14937,14942
sugar|14943,14948
control|14949,14956
<EOL>|14956,14957
<EOL>|14957,14958
It|14958,14960
was|14961,14964
a|14965,14966
pleasure|14967,14975
taking|14976,14982
care|14983,14987
of|14988,14990
you|14991,14994
!|14994,14995
<EOL>|14995,14996
<EOL>|14996,14997
Your|14997,15001
_|15002,15003
_|15003,15004
_|15004,15005
Inpatient|15006,15015
Care|15016,15020
Team|15021,15025
<EOL>|15025,15026
<EOL>|15027,15028
Followup|15028,15036
Instructions|15037,15049
:|15049,15050
<EOL>|15050,15051
_|15051,15052
_|15052,15053
_|15053,15054
<EOL>|15054,15055

