 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|50,59|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|50,59|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|50,64|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|84,93|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|84,93|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|84,93|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|84,93|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|84,93|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|84,98|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|116,121|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|116,121|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|116,121|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|140,143|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|140,143|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|140,143|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|140,143|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|140,143|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|151,158|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|151,158|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|160,168|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Drug|Organic Chemical|Allergies|183,191|false|false|false|C0086787|Percocet|Percocet
Drug|Pharmacologic Substance|Allergies|183,191|false|false|false|C0086787|Percocet|Percocet
Drug|Organic Chemical|Allergies|194,201|false|false|false|C0483514|Vicodin|Vicodin
Drug|Pharmacologic Substance|Allergies|194,201|false|false|false|C0483514|Vicodin|Vicodin
Event|Event|Allergies|204,213|false|false|false|||Attending
Finding|Functional Concept|Allergies|204,213|false|false|false|C1999232|Attending (action)|Attending
Anatomy|Body Location or Region|Chief Complaint|239,248|false|false|false|C0000726|Abdomen|Abdominal
Finding|Sign or Symptom|Chief Complaint|239,253|false|false|false|C0000737|Abdominal Pain|Abdominal pain
Attribute|Clinical Attribute|Chief Complaint|249,253|false|false|false|C2598155||pain
Event|Event|Chief Complaint|249,253|false|false|false|||pain
Finding|Functional Concept|Chief Complaint|249,253|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Chief Complaint|249,253|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Classification|Chief Complaint|256,261|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|262,270|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|262,270|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|274,292|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|283,292|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|283,292|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|283,292|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|283,292|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|283,292|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|Chief Complaint|298,310|false|false|false|||Paracentesis
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|298,310|false|false|false|C0034115|Paracentesis|Paracentesis
Disorder|Disease or Syndrome|History of Present Illness|349,352|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Disorder|Virus|History of Present Illness|349,352|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Drug|Immunologic Factor|History of Present Illness|349,352|false|false|false|C0086413|HIV Vaccine|HIV
Drug|Pharmacologic Substance|History of Present Illness|349,352|false|false|false|C0086413|HIV Vaccine|HIV
Event|Event|History of Present Illness|349,352|false|false|false|||HIV
Event|Event|History of Present Illness|356,361|false|false|false|||HAART
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|356,361|false|false|false|C0887947|Antiretroviral Therapy, Highly Active|HAART
Disorder|Disease or Syndrome|History of Present Illness|363,367|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|History of Present Illness|363,367|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|History of Present Illness|363,367|false|false|false|||COPD
Finding|Gene or Genome|History of Present Illness|363,367|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|History of Present Illness|374,378|false|false|false|||home
Finding|Idea or Concept|History of Present Illness|374,378|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|History of Present Illness|374,378|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|History of Present Illness|374,378|false|false|false|C1553498|home health encounter|home
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|390,393|false|false|false|C2744672|SAT1 protein, human|sat
Drug|Enzyme|History of Present Illness|390,393|false|false|false|C2744672|SAT1 protein, human|sat
Finding|Gene or Genome|History of Present Illness|390,393|false|false|false|C0871290;C1705827;C1822614|College Entrance Examination Board Scholastic Aptitude Test;SAT1 gene;SAT1 wt Allele|sat
Finding|Intellectual Product|History of Present Illness|390,393|false|false|false|C0871290;C1705827;C1822614|College Entrance Examination Board Scholastic Aptitude Test;SAT1 gene;SAT1 wt Allele|sat
Event|Event|History of Present Illness|413,422|false|false|false|||admission
Procedure|Health Care Activity|History of Present Illness|413,422|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Disorder|Disease or Syndrome|History of Present Illness|425,428|false|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|HCV
Disorder|Virus|History of Present Illness|425,428|false|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|HCV
Event|Event|History of Present Illness|425,428|false|false|false|||HCV
Disorder|Disease or Syndrome|History of Present Illness|429,438|false|false|false|C0023890;C1623038|Cirrhosis;Liver Cirrhosis|cirrhosis
Event|Event|History of Present Illness|429,438|false|false|false|||cirrhosis
Disorder|Disease or Syndrome|History of Present Illness|443,450|false|false|false|C0003962|Ascites|ascites
Event|Event|History of Present Illness|443,450|false|false|false|||ascites
Finding|Pathologic Function|History of Present Illness|443,450|false|false|false|C5441966|Peritoneal Effusion|ascites
Event|Event|History of Present Illness|451,460|false|false|false|||requiring
Drug|Organic Chemical|History of Present Illness|471,482|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Drug|Pharmacologic Substance|History of Present Illness|471,482|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Event|Event|History of Present Illness|471,482|false|false|false|||therapeutic
Finding|Functional Concept|History of Present Illness|471,482|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Finding|Intellectual Product|History of Present Illness|471,482|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|471,482|false|false|false|C0087111|Therapeutic procedure|therapeutic
Event|Event|History of Present Illness|483,495|false|false|false|||paracenteses
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|483,495|false|false|false|C0034115|Paracentesis|paracenteses
Anatomy|Body Location or Region|History of Present Illness|497,504|false|false|false|C0205054|Hepatic|hepatic
Disorder|Disease or Syndrome|History of Present Illness|497,519|false|false|false|C0019151|Hepatic Encephalopathy|hepatic encephalopathy
Disorder|Disease or Syndrome|History of Present Illness|505,519|false|false|false|C0085584|Encephalopathies|encephalopathy
Event|Event|History of Present Illness|505,519|false|false|false|||encephalopathy
Anatomy|Tissue|History of Present Illness|529,539|false|false|false|C0332835|Transplanted tissue|transplant
Finding|Finding|History of Present Illness|529,539|false|false|false|C0478647;C3841811|Transplant;Transplanted organ and tissue status|transplant
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|529,539|false|false|false|C0040732|Transplantation|transplant
Event|Event|History of Present Illness|540,544|false|false|false|||list
Finding|Intellectual Product|History of Present Illness|540,544|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|History of Present Illness|549,562|false|false|false|||comorbidities
Finding|Finding|History of Present Illness|549,562|false|false|false|C0009488|Comorbidity|comorbidities
Event|Event|History of Present Illness|578,583|false|false|false|||girth
Anatomy|Body Location or Region|History of Present Illness|588,591|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|abd
Disorder|Cell or Molecular Dysfunction|History of Present Illness|588,591|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|abd
Attribute|Clinical Attribute|History of Present Illness|593,597|false|false|false|C2598155||pain
Event|Event|History of Present Illness|593,597|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|593,597|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|593,597|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|History of Present Illness|617,621|false|false|false|C2598155||pain
Event|Event|History of Present Illness|617,621|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|617,621|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|617,621|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Disorder|Disease or Syndrome|History of Present Illness|631,638|false|false|false|C0003962|Ascites|ascites
Event|Event|History of Present Illness|631,638|false|false|false|||ascites
Finding|Pathologic Function|History of Present Illness|631,638|false|false|false|C5441966|Peritoneal Effusion|ascites
Event|Event|History of Present Illness|644,648|false|false|false|||felt
Event|Event|History of Present Illness|649,656|false|false|false|||overdue
Event|Event|History of Present Illness|664,676|false|false|false|||paracentesis
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|664,676|false|false|false|C0034115|Paracentesis|paracentesis
Event|Event|History of Present Illness|691,703|false|false|false|||paracentesis
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|691,703|false|false|false|C0034115|Paracentesis|paracentesis
Event|Event|History of Present Illness|721,729|false|false|false|||reported
Event|Event|History of Present Illness|739,744|false|false|false|||began
Event|Event|History of Present Illness|745,752|false|false|false|||feeling
Finding|Idea or Concept|History of Present Illness|753,762|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Anatomy|Body Location or Region|History of Present Illness|763,772|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|History of Present Illness|763,777|false|true|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|History of Present Illness|773,777|false|false|false|C2598155||pain
Event|Event|History of Present Illness|773,777|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|773,777|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|773,777|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Intellectual Product|History of Present Illness|780,788|false|false|false|C1720529|Constant - dosing instruction fragment|constant
Anatomy|Body Location or Region|History of Present Illness|790,800|false|false|false|C0521440|Epigastric|epigastric
Event|Event|History of Present Illness|805,813|false|false|false|||radiates
Drug|Food|History of Present Illness|831,835|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Drug|Immunologic Factor|History of Present Illness|831,835|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Drug|Pharmacologic Substance|History of Present Illness|831,835|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Event|Event|History of Present Illness|852,861|false|false|false|||increased
Finding|Idea or Concept|History of Present Illness|904,907|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|History of Present Illness|904,907|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|History of Present Illness|917,924|false|false|false|||brought
Finding|Gene or Genome|History of Present Illness|942,945|false|false|false|C1420310|SON gene|son
Attribute|Clinical Attribute|History of Present Illness|962,966|false|false|false|C2598155||pain
Event|Event|History of Present Illness|962,966|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|962,966|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|962,966|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|980,989|false|false|false|C0009676|Confusion|confusion
Event|Event|History of Present Illness|980,989|false|false|false|||confusion
Finding|Finding|History of Present Illness|980,989|false|false|false|C0683369|Clouded consciousness|confusion
Attribute|Clinical Attribute|History of Present Illness|998,1003|false|false|false|C5890168||alert
Drug|Organic Chemical|History of Present Illness|998,1003|false|false|false|C0718338|Alert brand of caffeine|alert
Drug|Pharmacologic Substance|History of Present Illness|998,1003|false|false|false|C0718338|Alert brand of caffeine|alert
Event|Event|History of Present Illness|998,1003|false|false|false|||alert
Finding|Finding|History of Present Illness|998,1003|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Functional Concept|History of Present Illness|998,1003|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Intellectual Product|History of Present Illness|998,1003|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Event|Event|History of Present Illness|1008,1016|false|false|false|||oriented
Finding|Finding|History of Present Illness|1008,1016|false|false|false|C1961028|Oriented to place|oriented
Finding|Body Substance|History of Present Illness|1025,1032|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1025,1032|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1025,1032|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|1039,1047|false|false|false|||reported
Event|Event|History of Present Illness|1061,1064|false|false|false|||ran
Event|Event|History of Present Illness|1084,1088|false|false|false|||home
Finding|Idea or Concept|History of Present Illness|1084,1088|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|History of Present Illness|1084,1088|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|History of Present Illness|1084,1088|false|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|History of Present Illness|1090,1101|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|History of Present Illness|1090,1101|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|History of Present Illness|1090,1101|false|false|false|||medications
Finding|Intellectual Product|History of Present Illness|1090,1101|false|false|false|C4284232|Medications|medications
Event|Event|History of Present Illness|1107,1113|false|false|false|||denied
Event|Event|History of Present Illness|1118,1123|false|false|false|||fever
Finding|Finding|History of Present Illness|1118,1123|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|History of Present Illness|1118,1123|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|History of Present Illness|1125,1131|false|false|false|||chills
Finding|Sign or Symptom|History of Present Illness|1125,1131|true|false|false|C0085593|Chills|chills
Event|Event|History of Present Illness|1133,1142|false|false|false|||shortness
Attribute|Clinical Attribute|History of Present Illness|1133,1152|true|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|History of Present Illness|1133,1152|true|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|History of Present Illness|1146,1152|false|false|false|C0225386|Breath|breath
Drug|Organic Chemical|History of Present Illness|1155,1160|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|1155,1160|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|History of Present Illness|1155,1160|false|false|false|||cough
Finding|Sign or Symptom|History of Present Illness|1155,1160|false|false|false|C0010200|Coughing|cough
Event|Event|History of Present Illness|1162,1169|false|false|false|||dysuria
Finding|Sign or Symptom|History of Present Illness|1162,1169|false|false|false|C0013428|Dysuria|dysuria
Event|Event|History of Present Illness|1175,1183|false|false|false|||reported
Finding|Sign or Symptom|History of Present Illness|1184,1195|false|false|false|C2129214|Loose stool|loose stool
Event|Event|History of Present Illness|1190,1195|false|false|false|||stool
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1198,1201|false|false|false|C0045724;C0671702|2-(4-ethoxybenzyl)-1-diethylaminoethyl-5-isothiocyanatobenzimidazole;PTPNS1 protein, human|bit
Drug|Organic Chemical|History of Present Illness|1198,1201|false|false|false|C0045724;C0671702|2-(4-ethoxybenzyl)-1-diethylaminoethyl-5-isothiocyanatobenzimidazole;PTPNS1 protein, human|bit
Drug|Pharmacologic Substance|History of Present Illness|1198,1201|false|false|false|C0045724;C0671702|2-(4-ethoxybenzyl)-1-diethylaminoethyl-5-isothiocyanatobenzimidazole;PTPNS1 protein, human|bit
Event|Event|History of Present Illness|1198,1201|false|false|false|||bit
Finding|Gene or Genome|History of Present Illness|1198,1201|false|false|false|C0671702;C1705300;C1822726;C4321288|Breast-Impact of Treatment Scale;PTPNS1 protein, human;SIRPA gene;SIRPA wt Allele|bit
Finding|Intellectual Product|History of Present Illness|1198,1201|false|false|false|C0671702;C1705300;C1822726;C4321288|Breast-Impact of Treatment Scale;PTPNS1 protein, human;SIRPA gene;SIRPA wt Allele|bit
Finding|Receptor|History of Present Illness|1198,1201|false|false|false|C0671702;C1705300;C1822726;C4321288|Breast-Impact of Treatment Scale;PTPNS1 protein, human;SIRPA gene;SIRPA wt Allele|bit
Event|Event|History of Present Illness|1224,1234|false|false|false|||attributed
Drug|Organic Chemical|History of Present Illness|1241,1250|false|false|false|C0022957|lactulose|lactulose
Drug|Pharmacologic Substance|History of Present Illness|1241,1250|false|false|false|C0022957|lactulose|lactulose
Event|Event|History of Present Illness|1251,1254|false|false|false|||use
Finding|Functional Concept|History of Present Illness|1251,1254|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|History of Present Illness|1251,1254|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Event|Event|History of Present Illness|1267,1273|false|false|false|||vitals
Event|Event|History of Present Illness|1308,1312|false|false|false|||Labs
Lab|Laboratory or Test Result|History of Present Illness|1308,1312|false|false|false|C0587081|Laboratory test finding|Labs
Event|Event|History of Present Illness|1318,1329|false|false|false|||significant
Finding|Idea or Concept|History of Present Illness|1318,1329|false|false|false|C0750502|Significant|significant
Event|Event|History of Present Illness|1334,1336|false|false|false|||Na
Drug|Organic Chemical|History of Present Illness|1348,1355|false|false|false|C0022924;C0376261|Lactates;lactate|lactate
Drug|Pharmacologic Substance|History of Present Illness|1348,1355|false|false|false|C0022924;C0376261|Lactates;lactate|lactate
Event|Event|History of Present Illness|1348,1355|false|false|false|||lactate
Procedure|Laboratory Procedure|History of Present Illness|1348,1355|false|false|false|C0202115|Lactic acid measurement|lactate
Attribute|Clinical Attribute|History of Present Illness|1360,1363|false|false|false|C0368980|Coagulation tissue factor induced.INR|INR
Event|Event|History of Present Illness|1360,1363|false|false|false|||INR
Procedure|Laboratory Procedure|History of Present Illness|1360,1363|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1360,1363|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Disorder|Neoplastic Process|History of Present Illness|1369,1372|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1369,1372|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|History of Present Illness|1369,1372|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|History of Present Illness|1369,1372|false|false|false|||ALT
Finding|Gene or Genome|History of Present Illness|1369,1372|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|History of Present Illness|1369,1372|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|History of Present Illness|1369,1372|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1369,1372|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|History of Present Illness|1377,1380|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|History of Present Illness|1377,1380|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1377,1380|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|History of Present Illness|1377,1380|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|History of Present Illness|1377,1380|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|History of Present Illness|1377,1380|false|false|false|||AST
Finding|Gene or Genome|History of Present Illness|1377,1380|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Disorder|Disease or Syndrome|History of Present Illness|1396,1408|true|false|false|C0023518|Leukocytosis|leukocytosis
Event|Event|History of Present Illness|1396,1408|false|false|false|||leukocytosis
Finding|Finding|History of Present Illness|1396,1408|true|false|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Finding|Body Substance|History of Present Illness|1411,1424|false|false|false|C5441965|Ascitic Fluid|Ascitic fluid
Drug|Substance|History of Present Illness|1419,1424|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|History of Present Illness|1419,1424|false|false|false|||fluid
Finding|Intellectual Product|History of Present Illness|1419,1424|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|History of Present Illness|1425,1431|false|false|false|||showed
Anatomy|Cell|History of Present Illness|1436,1439|false|false|false|C0023516|Leukocytes|WBC
Event|Event|History of Present Illness|1436,1439|false|false|false|||WBC
Drug|Organic Chemical|History of Present Illness|1455,1463|false|false|false|C0026549|morphine|Morphine
Drug|Pharmacologic Substance|History of Present Illness|1455,1463|false|false|false|C0026549|morphine|Morphine
Event|Event|History of Present Illness|1455,1463|false|false|false|||Morphine
Drug|Organic Chemical|History of Present Illness|1455,1471|false|false|false|C0066814|morphine sulfate|Morphine Sulfate
Drug|Pharmacologic Substance|History of Present Illness|1455,1471|false|false|false|C0066814|morphine sulfate|Morphine Sulfate
Drug|Element, Ion, or Isotope|History of Present Illness|1464,1471|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Inorganic Chemical|History of Present Illness|1464,1471|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Pharmacologic Substance|History of Present Illness|1464,1471|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Event|Event|History of Present Illness|1472,1473|false|false|false|||5
Finding|Intellectual Product|History of Present Illness|1481,1485|false|false|false|C1720092|Once - dosing instruction fragment|ONCE
Event|Event|History of Present Illness|1486,1489|false|false|false|||MR1
Finding|Gene or Genome|History of Present Illness|1486,1489|false|false|false|C1415592;C1418706|MR1 gene;PNKD gene|MR1
Drug|Food|History of Present Illness|1500,1508|false|false|false|C0678420|Cocktail|cocktail
Event|Event|History of Present Illness|1500,1508|false|false|false|||cocktail
Disorder|Disease or Syndrome|Past Medical History|1536,1539|false|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|HCV
Disorder|Virus|Past Medical History|1536,1539|false|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|HCV
Event|Event|Past Medical History|1536,1539|false|false|false|||HCV
Disorder|Disease or Syndrome|Past Medical History|1540,1549|false|false|false|C0023890;C1623038|Cirrhosis;Liver Cirrhosis|Cirrhosis
Event|Event|Past Medical History|1540,1549|false|false|false|||Cirrhosis
Event|Event|Past Medical History|1551,1559|false|false|false|||genotype
Procedure|Laboratory Procedure|Past Medical History|1551,1559|false|false|false|C1285573|Genotype determination|genotype
Disorder|Disease or Syndrome|Past Medical History|1567,1570|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Disorder|Virus|Past Medical History|1567,1570|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Drug|Immunologic Factor|Past Medical History|1567,1570|false|false|false|C0086413|HIV Vaccine|HIV
Drug|Pharmacologic Substance|Past Medical History|1567,1570|false|false|false|C0086413|HIV Vaccine|HIV
Event|Event|Past Medical History|1567,1570|false|false|false|||HIV
Event|Event|Past Medical History|1575,1580|false|false|false|||HAART
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1575,1580|false|false|false|C0887947|Antiretroviral Therapy, Highly Active|HAART
Drug|Amino Acid, Peptide, or Protein|Past Medical History|1586,1589|false|false|false|C0003323;C4048280|CD4 Antigens;T-Cell Surface Glycoprotein CD4, human|CD4
Drug|Biologically Active Substance|Past Medical History|1586,1589|false|false|false|C0003323;C4048280|CD4 Antigens;T-Cell Surface Glycoprotein CD4, human|CD4
Drug|Immunologic Factor|Past Medical History|1586,1589|false|false|false|C0003323;C4048280|CD4 Antigens;T-Cell Surface Glycoprotein CD4, human|CD4
Finding|Gene or Genome|Past Medical History|1586,1589|false|false|false|C0003323;C1332714|CD4 Antigens;CD4 gene|CD4
Finding|Receptor|Past Medical History|1586,1589|false|false|false|C0003323;C1332714|CD4 Antigens;CD4 gene|CD4
Procedure|Laboratory Procedure|Past Medical History|1586,1595|false|false|false|C0243009;C3541261|CD4 Count determination procedure;CD4 Expressing Cell Count|CD4 count
Event|Event|Past Medical History|1590,1595|false|false|false|||count
Disorder|Disease or Syndrome|Past Medical History|1605,1608|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Disorder|Virus|Past Medical History|1605,1608|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Drug|Immunologic Factor|Past Medical History|1605,1608|false|false|false|C0086413|HIV Vaccine|HIV
Drug|Pharmacologic Substance|Past Medical History|1605,1608|false|false|false|C0086413|HIV Vaccine|HIV
Event|Event|Past Medical History|1605,1608|false|false|false|||HIV
Procedure|Laboratory Procedure|Past Medical History|1605,1619|false|false|false|C1168369|HIV viral load|HIV viral load
Finding|Functional Concept|Past Medical History|1609,1614|false|false|false|C0521026|Viral|viral
Finding|Finding|Past Medical History|1609,1619|false|false|false|C0376705|Viral Load result|viral load
Procedure|Laboratory Procedure|Past Medical History|1609,1619|false|false|false|C1261478|Viral load (procedure)|viral load
Event|Activity|Past Medical History|1615,1619|false|false|false|C1708715|Loading Technique|load
Event|Event|Past Medical History|1615,1619|false|false|false|||load
Finding|Idea or Concept|Past Medical History|1615,1619|false|false|false|C1550025|Load - Remote control command|load
Attribute|Clinical Attribute|Past Medical History|1621,1633|false|false|false|C3827727|Undetectable|undetectable
Disorder|Disease or Syndrome|Past Medical History|1638,1642|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Past Medical History|1638,1642|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Past Medical History|1638,1642|false|false|false|||COPD
Finding|Gene or Genome|Past Medical History|1638,1642|false|false|false|C1412502|ARCN1 gene|COPD
Anatomy|Body Location or Region|Past Medical History|1648,1651|false|false|false|C5239891|area PFt|PFT
Drug|Indicator, Reagent, or Diagnostic Aid|Past Medical History|1648,1651|false|false|false|C0053122|bentiromide|PFT
Drug|Pharmacologic Substance|Past Medical History|1648,1651|false|false|false|C0053122|bentiromide|PFT
Event|Event|Past Medical History|1648,1651|false|false|false|||PFT
Procedure|Diagnostic Procedure|Past Medical History|1648,1651|false|false|false|C0024119;C0279232|Pulmonary function tests;fluorouracil/melphalan/tamoxifen|PFT
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1648,1651|false|false|false|C0024119;C0279232|Pulmonary function tests;fluorouracil/melphalan/tamoxifen|PFT
Event|Event|Past Medical History|1652,1658|false|false|false|||showed
Event|Event|Past Medical History|1659,1662|false|false|false|||FVC
Lab|Laboratory or Test Result|Past Medical History|1659,1662|false|false|false|C3714541|Forced Vital Capacity|FVC
Attribute|Clinical Attribute|Past Medical History|1675,1679|false|false|false|C0802965||FEV1
Event|Event|Past Medical History|1675,1679|false|false|false|||FEV1
Procedure|Diagnostic Procedure|Past Medical History|1675,1679|false|false|false|C0849974|Pulmonary Function Test/Forced Expiratory Volume 1|FEV1
Disorder|Mental or Behavioral Dysfunction|Past Medical History|1715,1741|false|false|false|C0005586;C1839839;C1852197;C1970943;C1970945;C2700438;C2700439;C2700440|Bipolar Disorder;MAJOR AFFECTIVE DISORDER 1;MAJOR AFFECTIVE DISORDER 2;MAJOR AFFECTIVE DISORDER 4;MAJOR AFFECTIVE DISORDER 6;MAJOR AFFECTIVE DISORDER 7;MAJOR AFFECTIVE DISORDER 8;MAJOR AFFECTIVE DISORDER 9|Bipolar Affective Disorder
Disorder|Mental or Behavioral Dysfunction|Past Medical History|1723,1741|false|false|false|C0525045|Mood Disorders|Affective Disorder
Disorder|Disease or Syndrome|Past Medical History|1733,1741|false|false|false|C0012634|Disease|Disorder
Event|Event|Past Medical History|1733,1741|false|false|false|||Disorder
Disorder|Disease or Syndrome|Past Medical History|1746,1750|false|false|false|C0038436;C0878676|6-pyruvoyl-tetrahydropterin synthase deficiency;Post-Traumatic Stress Disorder|PTSD
Disorder|Mental or Behavioral Dysfunction|Past Medical History|1746,1750|false|false|false|C0038436;C0878676|6-pyruvoyl-tetrahydropterin synthase deficiency;Post-Traumatic Stress Disorder|PTSD
Event|Event|Past Medical History|1746,1750|false|false|false|||PTSD
Disorder|Injury or Poisoning|Past Medical History|1761,1768|false|false|false|C0274659|Poisoning by cocaine|cocaine
Drug|Biomedical or Dental Material|Past Medical History|1761,1768|false|false|false|C0009170|cocaine|cocaine
Drug|Hazardous or Poisonous Substance|Past Medical History|1761,1768|false|false|false|C0009170|cocaine|cocaine
Drug|Organic Chemical|Past Medical History|1761,1768|false|false|false|C0009170|cocaine|cocaine
Drug|Pharmacologic Substance|Past Medical History|1761,1768|false|false|false|C0009170|cocaine|cocaine
Event|Event|Past Medical History|1761,1768|false|false|false|||cocaine
Procedure|Laboratory Procedure|Past Medical History|1761,1768|false|false|false|C0202362|Cocaine measurement|cocaine
Disorder|Injury or Poisoning|Past Medical History|1773,1779|false|false|false|C0161541|Poisoning by heroin|heroin
Drug|Hazardous or Poisonous Substance|Past Medical History|1773,1779|false|false|false|C0011892|heroin|heroin
Drug|Organic Chemical|Past Medical History|1773,1779|false|false|false|C0011892|heroin|heroin
Drug|Pharmacologic Substance|Past Medical History|1773,1779|false|false|false|C0011892|heroin|heroin
Event|Event|Past Medical History|1773,1779|false|false|false|||heroin
Disorder|Mental or Behavioral Dysfunction|Past Medical History|1773,1785|false|false|false|C0600241|heroin abuse|heroin abuse
Disorder|Mental or Behavioral Dysfunction|Past Medical History|1780,1785|false|false|false|C0013146|Drug abuse|abuse
Event|Event|Past Medical History|1780,1785|false|false|false|||abuse
Event|Event|Past Medical History|1780,1785|false|false|false|C1546935|Abuse|abuse
Finding|Finding|Past Medical History|1780,1785|false|false|false|C0562381|Victim of abuse (finding)|abuse
Disorder|Neoplastic Process|Past Medical History|1793,1807|false|false|false|C0007114|Malignant neoplasm of skin|of skin cancer
Anatomy|Body System|Past Medical History|1796,1800|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|Past Medical History|1796,1800|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|Past Medical History|1796,1800|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Finding|Body Substance|Past Medical History|1796,1800|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|Past Medical History|1796,1800|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Disorder|Neoplastic Process|Past Medical History|1796,1807|false|false|false|C0007114|Malignant neoplasm of skin|skin cancer
Disorder|Neoplastic Process|Past Medical History|1801,1807|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Past Medical History|1801,1807|false|false|false|||cancer
Finding|Body Substance|Past Medical History|1812,1819|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Past Medical History|1812,1819|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Past Medical History|1812,1819|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Past Medical History|1812,1826|false|false|false|C0747307|Patient-Reported|patient report
Attribute|Clinical Attribute|Past Medical History|1820,1826|false|false|false|C4255046||report
Event|Event|Past Medical History|1820,1826|false|false|false|||report
Finding|Intellectual Product|Past Medical History|1820,1826|false|false|false|C0684224|Report (document)|report
Procedure|Health Care Activity|Past Medical History|1820,1826|false|false|false|C0700287|Reporting|report
Event|Event|Family Medical History|1913,1920|false|false|false|||talking
Finding|Conceptual Entity|Family Medical History|1956,1963|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|brother
Finding|Idea or Concept|Family Medical History|1956,1963|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|brother
Event|Event|Family Medical History|1979,1984|false|false|false|||touch
Finding|Mental Process|Family Medical History|1979,1984|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Finding|Organ or Tissue Function|Family Medical History|1979,1984|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Procedure|Therapeutic or Preventive Procedure|Family Medical History|1979,1984|false|false|false|C0152054|Therapeutic Touch|touch
Event|Event|Family Medical History|1995,2000|false|false|false|||lives
Event|Event|Family Medical History|2020,2025|false|false|false|||aware
Finding|Mental Process|Family Medical History|2020,2025|true|false|false|C0004448|Awareness|aware
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2045,2050|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Family Medical History|2045,2050|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Family Medical History|2045,2050|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Family Medical History|2045,2050|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Family Medical History|2045,2050|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Family Medical History|2045,2050|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|Family Medical History|2045,2050|false|false|false|||liver
Finding|Finding|Family Medical History|2045,2050|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Family Medical History|2045,2050|false|false|false|C0872387|Procedures on liver|liver
Disorder|Disease or Syndrome|Family Medical History|2052,2059|false|false|false|C0012634|Disease|disease
Event|Event|Family Medical History|2052,2059|false|false|false|||disease
Drug|Amino Acid, Peptide, or Protein|Family Medical History|2063,2073|false|false|false|C3812393|ErbB Receptors|her family
Drug|Enzyme|Family Medical History|2063,2073|false|false|false|C3812393|ErbB Receptors|her family
Finding|Receptor|Family Medical History|2063,2073|false|false|false|C3812393|ErbB Receptors|her family
Finding|Classification|Family Medical History|2067,2073|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Family Medical History|2067,2073|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Family Medical History|2067,2073|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Family Medical History|2067,2073|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Procedure|Health Care Activity|General Exam|2094,2103|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|General Exam|2104,2112|false|false|false|||PHYSICAL
Finding|Finding|General Exam|2104,2112|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|General Exam|2104,2112|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|General Exam|2104,2112|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|General Exam|2104,2117|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|General Exam|2104,2117|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Event|Event|General Exam|2113,2117|false|false|false|||EXAM
Finding|Functional Concept|General Exam|2113,2117|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|2113,2117|false|false|false|C0582103|Medical Examination|EXAM
Drug|Biologically Active Substance|General Exam|2191,2198|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|2191,2198|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|2191,2198|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|2191,2198|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|2191,2198|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|2191,2198|false|false|false|C0337438|Glucose measurement|Glucose
Event|Event|General Exam|2206,2213|false|false|false|||GENERAL
Finding|Classification|General Exam|2206,2213|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|General Exam|2206,2213|false|false|false|C3812897|General medical service|GENERAL
Disorder|Disease or Syndrome|General Exam|2215,2218|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|2215,2218|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|2215,2218|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|2215,2218|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|2215,2218|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|General Exam|2215,2218|false|false|false|||NAD
Finding|Finding|General Exam|2215,2218|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Event|Event|General Exam|2220,2225|false|false|false|||lying
Finding|Functional Concept|General Exam|2233,2238|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|General Exam|2245,2250|false|false|false|C1512338|HEENT|HEENT
Event|Event|General Exam|2259,2263|false|false|false|||EOMI
Event|Event|General Exam|2265,2270|false|false|false|||PERRL
Finding|Finding|General Exam|2265,2270|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Finding|Finding|General Exam|2272,2281|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|General Exam|2282,2288|false|false|false|C0036410|Sclera|sclera
Disorder|Disease or Syndrome|General Exam|2282,2288|false|false|false|C0036412|Scleral Diseases|sclera
Event|Event|General Exam|2282,2288|false|false|false|||sclera
Procedure|Health Care Activity|General Exam|2282,2288|false|false|false|C2228481|examination of sclera|sclera
Anatomy|Body Part, Organ, or Organ Component|General Exam|2295,2306|false|false|false|C0009758;C0229274|Structure of palpebral conjunctiva;conjunctiva|conjunctiva
Disorder|Disease or Syndrome|General Exam|2295,2306|false|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|conjunctiva
Disorder|Neoplastic Process|General Exam|2295,2306|false|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|conjunctiva
Event|Event|General Exam|2295,2306|false|false|false|||conjunctiva
Finding|Body Substance|General Exam|2295,2306|false|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|conjunctiva
Finding|Intellectual Product|General Exam|2295,2306|false|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|conjunctiva
Procedure|Health Care Activity|General Exam|2295,2306|false|false|false|C0872390;C2228431|Procedure on conjunctiva;examination of conjunctiva|conjunctiva
Anatomy|Body Part, Organ, or Organ Component|General Exam|2309,2312|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|General Exam|2309,2312|false|false|false|C0026987|Myelofibrosis|MMM
Event|Event|General Exam|2309,2312|false|false|false|||MMM
Finding|Idea or Concept|General Exam|2314,2318|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Anatomy|Body Part, Organ, or Organ Component|General Exam|2319,2328|false|false|false|C0011443;C0040426|Dentition;Tooth structure|dentition
Anatomy|Body Location or Region|General Exam|2331,2335|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|General Exam|2331,2335|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|General Exam|2331,2335|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Finding|Functional Concept|General Exam|2347,2353|false|false|false|C0332254|Supple|supple
Finding|Finding|General Exam|2347,2358|false|false|false|C2230237|Supple neck|supple neck
Anatomy|Body Location or Region|General Exam|2354,2358|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|General Exam|2354,2358|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|General Exam|2354,2358|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Anatomy|Body Part, Organ, or Organ Component|General Exam|2363,2366|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|General Exam|2363,2366|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|General Exam|2363,2366|false|false|false|||LAD
Finding|Gene or Genome|General Exam|2363,2366|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Event|General Exam|2371,2374|false|false|false|||JVD
Finding|Finding|General Exam|2371,2374|true|false|false|C0425687|Jugular venous engorgement|JVD
Anatomy|Body Part, Organ, or Organ Component|General Exam|2377,2384|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|General Exam|2377,2384|false|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Event|General Exam|2386,2389|false|false|false|||RRR
Event|Event|General Exam|2401,2408|false|false|false|||murmurs
Finding|Finding|General Exam|2401,2408|true|false|false|C0018808|Heart murmur|murmurs
Event|Event|General Exam|2410,2417|false|false|false|||gallops
Event|Event|General Exam|2422,2426|false|false|false|||rubs
Finding|Finding|General Exam|2422,2426|true|false|false|C0232267|Pericardial friction rub|rubs
Anatomy|Body Location or Region|General Exam|2429,2433|false|false|false|C0024109;C4037972|Chest>Lung;Lung|LUNG
Anatomy|Body Part, Organ, or Organ Component|General Exam|2429,2433|false|false|false|C0024109;C4037972|Chest>Lung;Lung|LUNG
Disorder|Disease or Syndrome|General Exam|2429,2433|false|false|false|C0024115|Lung diseases|LUNG
Event|Event|General Exam|2429,2433|false|false|false|||LUNG
Finding|Finding|General Exam|2429,2433|false|false|false|C0740941|Lung Problem|LUNG
Drug|Organic Chemical|General Exam|2435,2439|false|false|false|C0951233|cetrimonium bromide|CTAB
Event|Event|General Exam|2435,2439|false|false|false|||CTAB
Event|Event|General Exam|2444,2451|false|false|false|||wheezes
Finding|Sign or Symptom|General Exam|2444,2451|true|false|false|C0043144|Wheezing|wheezes
Event|Event|General Exam|2453,2458|false|false|false|||rales
Finding|Finding|General Exam|2453,2458|true|false|false|C0034642;C0240859|Basilar Rales;Rales|rales
Event|Event|General Exam|2460,2467|false|false|false|||rhonchi
Finding|Finding|General Exam|2460,2467|true|false|false|C0035508|Rhonchi|rhonchi
Event|Event|General Exam|2469,2478|false|false|false|||breathing
Event|Event|General Exam|2500,2503|false|false|false|||use
Finding|Functional Concept|General Exam|2500,2503|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|General Exam|2500,2503|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Functional Concept|General Exam|2500,2506|true|false|false|C1524063|Use of|use of
Finding|Finding|General Exam|2500,2524|true|false|false|C1821466|Use of accessory muscles|use of accessory muscles
Disorder|Congenital Abnormality|General Exam|2507,2524|false|false|false|C0158784|Accessory skeletal muscle|accessory muscles
Anatomy|Body Part, Organ, or Organ Component|General Exam|2517,2524|false|false|false|C0026845;C1995013;C4083049|Muscle (organ);Muscle Tissue;Set of muscles|muscles
Anatomy|Tissue|General Exam|2517,2524|false|false|false|C0026845;C1995013;C4083049|Muscle (organ);Muscle Tissue;Set of muscles|muscles
Anatomy|Body Location or Region|General Exam|2527,2534|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|General Exam|2527,2534|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|General Exam|2527,2534|false|false|false|||ABDOMEN
Finding|Finding|General Exam|2527,2534|false|false|false|C0941288|Abdomen problem|ABDOMEN
Event|Event|General Exam|2536,2545|false|false|false|||distended
Finding|Finding|General Exam|2536,2545|false|false|false|C0700124|Dilated|distended
Drug|Substance|General Exam|2549,2554|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|General Exam|2549,2554|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Finding|General Exam|2549,2559|false|false|false|C0426682|Fluid thrill in abdomen|fluid wave
Event|Event|General Exam|2555,2559|false|false|false|||wave
Finding|Gene or Genome|General Exam|2555,2559|false|false|false|C1421479|WASF1 gene|wave
Phenomenon|Natural Phenomenon or Process|General Exam|2555,2559|false|false|false|C0678544||wave
Disorder|Mental or Behavioral Dysfunction|General Exam|2565,2570|true|false|false|C0233494|Tension|tense
Event|Event|General Exam|2565,2570|false|false|false|||tense
Finding|Sign or Symptom|General Exam|2565,2570|true|false|false|C0235108|Feeling tense|tense
Event|Event|General Exam|2572,2576|false|false|false|||NABS
Event|Event|General Exam|2578,2587|false|false|false|||nontender
Anatomy|Body Part, Organ, or Organ Component|General Exam|2590,2601|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Event|Event|General Exam|2606,2614|false|false|false|||cyanosis
Finding|Sign or Symptom|General Exam|2606,2614|true|false|false|C0010520|Cyanosis|cyanosis
Disorder|Anatomical Abnormality|General Exam|2616,2624|true|false|false|C0149651|Clubbing|clubbing
Event|Event|General Exam|2616,2624|false|false|false|||clubbing
Attribute|Clinical Attribute|General Exam|2628,2633|true|false|false|C1717255||edema
Event|Event|General Exam|2628,2633|false|false|false|||edema
Finding|Pathologic Function|General Exam|2628,2633|true|false|false|C0013604|Edema|edema
Event|Event|General Exam|2635,2641|false|false|false|||moving
Anatomy|Body Part, Organ, or Organ Component|General Exam|2649,2660|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Event|Event|General Exam|2649,2660|false|false|false|||extremities
Drug|Organic Chemical|General Exam|2666,2673|false|false|false|C1995603|PURPOSE (pharmacologic preparation)|purpose
Drug|Pharmacologic Substance|General Exam|2666,2673|false|false|false|C1995603|PURPOSE (pharmacologic preparation)|purpose
Event|Event|General Exam|2666,2673|false|false|false|||purpose
Finding|Functional Concept|General Exam|2666,2673|false|false|false|C1285529|Purpose|purpose
Drug|Food|General Exam|2674,2680|false|false|false|C5890763||PULSES
Event|Event|General Exam|2674,2680|false|false|false|||PULSES
Finding|Physiologic Function|General Exam|2674,2680|false|false|false|C0391850|Physiologic pulse|PULSES
Procedure|Health Care Activity|General Exam|2674,2680|false|false|false|C0034107|Pulse taking|PULSES
Drug|Food|General Exam|2688,2694|false|false|false|C5890763||pulses
Event|Event|General Exam|2688,2694|false|false|false|||pulses
Finding|Physiologic Function|General Exam|2688,2694|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|2688,2694|false|false|false|C0034107|Pulse taking|pulses
Event|Event|General Exam|2726,2732|false|false|false|||intact
Finding|Finding|General Exam|2726,2732|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Molecular Function|General Exam|2734,2738|false|false|false|C1817552|abscisic aldehyde oxidase activity|AAO3
Event|Event|General Exam|2743,2751|false|false|false|||asterxis
Anatomy|Body System|General Exam|2754,2758|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|General Exam|2754,2758|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|General Exam|2754,2758|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|General Exam|2754,2758|false|false|false|||SKIN
Finding|Body Substance|General Exam|2754,2758|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|General Exam|2754,2758|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Event|Event|General Exam|2760,2764|false|false|false|||warm
Finding|Finding|General Exam|2760,2764|false|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|General Exam|2760,2764|false|false|false|C0687712|warming process|warm
Finding|Finding|General Exam|2769,2773|false|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|2774,2782|false|false|false|||perfused
Disorder|Injury or Poisoning|General Exam|2787,2799|true|false|false|C0015256|Excoriation|excoriations
Event|Event|General Exam|2787,2799|false|false|false|||excoriations
Event|Event|General Exam|2803,2810|false|false|false|||lesions
Finding|Finding|General Exam|2803,2810|true|false|false|C0221198|Lesion|lesions
Event|Event|General Exam|2816,2822|false|false|false|||rashes
Finding|Sign or Symptom|General Exam|2816,2822|false|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Finding|Body Substance|General Exam|2824,2833|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|2824,2833|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|2824,2833|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|2824,2833|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|General Exam|2834,2842|false|false|false|||PHYSICAL
Finding|Finding|General Exam|2834,2842|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|General Exam|2834,2842|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|General Exam|2834,2842|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|General Exam|2834,2847|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|General Exam|2834,2847|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Event|Event|General Exam|2843,2847|false|false|false|||EXAM
Finding|Functional Concept|General Exam|2843,2847|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|2843,2847|false|false|false|C0582103|Medical Examination|EXAM
Event|Event|General Exam|2899,2901|false|false|false|||BP
Event|Event|General Exam|2948,2955|false|false|false|||GENERAL
Finding|Classification|General Exam|2948,2955|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|General Exam|2948,2955|false|false|false|C3812897|General medical service|GENERAL
Disorder|Disease or Syndrome|General Exam|2957,2960|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|2957,2960|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|2957,2960|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|2957,2960|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|2957,2960|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|General Exam|2957,2960|false|false|false|||NAD
Finding|Finding|General Exam|2957,2960|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Event|Event|General Exam|2962,2967|false|false|false|||lying
Finding|Functional Concept|General Exam|2975,2980|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|General Exam|2987,2992|false|false|false|C1512338|HEENT|HEENT
Event|Event|General Exam|3001,3005|false|false|false|||EOMI
Event|Event|General Exam|3007,3012|false|false|false|||PERRL
Finding|Finding|General Exam|3007,3012|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Finding|Finding|General Exam|3014,3023|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|General Exam|3024,3030|false|false|false|C0036410|Sclera|sclera
Disorder|Disease or Syndrome|General Exam|3024,3030|false|false|false|C0036412|Scleral Diseases|sclera
Event|Event|General Exam|3024,3030|false|false|false|||sclera
Procedure|Health Care Activity|General Exam|3024,3030|false|false|false|C2228481|examination of sclera|sclera
Anatomy|Body Part, Organ, or Organ Component|General Exam|3037,3048|false|false|false|C0009758;C0229274|Structure of palpebral conjunctiva;conjunctiva|conjunctiva
Disorder|Disease or Syndrome|General Exam|3037,3048|false|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|conjunctiva
Disorder|Neoplastic Process|General Exam|3037,3048|false|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|conjunctiva
Event|Event|General Exam|3037,3048|false|false|false|||conjunctiva
Finding|Body Substance|General Exam|3037,3048|false|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|conjunctiva
Finding|Intellectual Product|General Exam|3037,3048|false|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|conjunctiva
Procedure|Health Care Activity|General Exam|3037,3048|false|false|false|C0872390;C2228431|Procedure on conjunctiva;examination of conjunctiva|conjunctiva
Anatomy|Body Part, Organ, or Organ Component|General Exam|3051,3054|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|General Exam|3051,3054|false|false|false|C0026987|Myelofibrosis|MMM
Event|Event|General Exam|3051,3054|false|false|false|||MMM
Finding|Idea or Concept|General Exam|3056,3060|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Anatomy|Body Part, Organ, or Organ Component|General Exam|3061,3070|false|false|false|C0011443;C0040426|Dentition;Tooth structure|dentition
Anatomy|Body Location or Region|General Exam|3073,3077|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|General Exam|3073,3077|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|General Exam|3073,3077|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Finding|Functional Concept|General Exam|3089,3095|false|false|false|C0332254|Supple|supple
Finding|Finding|General Exam|3089,3100|false|false|false|C2230237|Supple neck|supple neck
Anatomy|Body Location or Region|General Exam|3096,3100|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|General Exam|3096,3100|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|General Exam|3096,3100|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Anatomy|Body Part, Organ, or Organ Component|General Exam|3105,3108|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|General Exam|3105,3108|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|General Exam|3105,3108|false|false|false|||LAD
Finding|Gene or Genome|General Exam|3105,3108|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Event|General Exam|3113,3116|false|false|false|||JVD
Finding|Finding|General Exam|3113,3116|true|false|false|C0425687|Jugular venous engorgement|JVD
Anatomy|Body Part, Organ, or Organ Component|General Exam|3119,3126|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|General Exam|3119,3126|false|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Event|General Exam|3128,3131|false|false|false|||RRR
Event|Event|General Exam|3143,3150|false|false|false|||murmurs
Finding|Finding|General Exam|3143,3150|true|false|false|C0018808|Heart murmur|murmurs
Event|Event|General Exam|3152,3159|false|false|false|||gallops
Event|Event|General Exam|3164,3168|false|false|false|||rubs
Finding|Finding|General Exam|3164,3168|true|false|false|C0232267|Pericardial friction rub|rubs
Anatomy|Body Location or Region|General Exam|3171,3175|false|false|false|C0024109;C4037972|Chest>Lung;Lung|LUNG
Anatomy|Body Part, Organ, or Organ Component|General Exam|3171,3175|false|false|false|C0024109;C4037972|Chest>Lung;Lung|LUNG
Disorder|Disease or Syndrome|General Exam|3171,3175|false|false|false|C0024115|Lung diseases|LUNG
Event|Event|General Exam|3171,3175|false|false|false|||LUNG
Finding|Finding|General Exam|3171,3175|false|false|false|C0740941|Lung Problem|LUNG
Drug|Organic Chemical|General Exam|3177,3181|false|false|false|C0951233|cetrimonium bromide|CTAB
Event|Event|General Exam|3177,3181|false|false|false|||CTAB
Event|Event|General Exam|3186,3193|false|false|false|||wheezes
Finding|Sign or Symptom|General Exam|3186,3193|true|false|false|C0043144|Wheezing|wheezes
Event|Event|General Exam|3195,3200|false|false|false|||rales
Finding|Finding|General Exam|3195,3200|true|false|false|C0034642;C0240859|Basilar Rales;Rales|rales
Event|Event|General Exam|3202,3209|false|false|false|||rhonchi
Finding|Finding|General Exam|3202,3209|true|false|false|C0035508|Rhonchi|rhonchi
Event|Event|General Exam|3211,3220|false|false|false|||breathing
Event|Event|General Exam|3242,3245|false|false|false|||use
Finding|Functional Concept|General Exam|3242,3245|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|General Exam|3242,3245|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Functional Concept|General Exam|3242,3248|true|false|false|C1524063|Use of|use of
Finding|Finding|General Exam|3242,3266|true|false|false|C1821466|Use of accessory muscles|use of accessory muscles
Disorder|Congenital Abnormality|General Exam|3249,3266|false|false|false|C0158784|Accessory skeletal muscle|accessory muscles
Anatomy|Body Part, Organ, or Organ Component|General Exam|3259,3266|false|false|false|C0026845;C1995013;C4083049|Muscle (organ);Muscle Tissue;Set of muscles|muscles
Anatomy|Tissue|General Exam|3259,3266|false|false|false|C0026845;C1995013;C4083049|Muscle (organ);Muscle Tissue;Set of muscles|muscles
Anatomy|Body Location or Region|General Exam|3269,3276|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|General Exam|3269,3276|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|General Exam|3269,3276|false|false|false|||ABDOMEN
Finding|Finding|General Exam|3269,3276|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|General Exam|3278,3282|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|General Exam|3278,3282|false|false|false|||soft
Finding|Finding|General Exam|3284,3293|false|false|false|C0392756;C0442797|Decreasing;Reduced|decreased
Event|Event|General Exam|3294,3304|false|false|false|||distension
Finding|Finding|General Exam|3294,3304|true|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distension
Finding|Pathologic Function|General Exam|3294,3304|true|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distension
Disorder|Mental or Behavioral Dysfunction|General Exam|3310,3315|true|false|false|C0233494|Tension|tense
Event|Event|General Exam|3310,3315|false|false|false|||tense
Finding|Sign or Symptom|General Exam|3310,3315|true|false|false|C0235108|Feeling tense|tense
Event|Event|General Exam|3317,3321|false|false|false|||NABS
Event|Event|General Exam|3323,3332|false|false|false|||nontender
Anatomy|Body Part, Organ, or Organ Component|General Exam|3336,3347|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Event|Event|General Exam|3352,3360|false|false|false|||cyanosis
Finding|Sign or Symptom|General Exam|3352,3360|true|false|false|C0010520|Cyanosis|cyanosis
Disorder|Anatomical Abnormality|General Exam|3362,3370|true|false|false|C0149651|Clubbing|clubbing
Event|Event|General Exam|3362,3370|false|false|false|||clubbing
Attribute|Clinical Attribute|General Exam|3374,3379|true|false|false|C1717255||edema
Event|Event|General Exam|3374,3379|false|false|false|||edema
Finding|Pathologic Function|General Exam|3374,3379|true|false|false|C0013604|Edema|edema
Event|Event|General Exam|3381,3387|false|false|false|||moving
Anatomy|Body Part, Organ, or Organ Component|General Exam|3395,3406|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Event|Event|General Exam|3395,3406|false|false|false|||extremities
Drug|Organic Chemical|General Exam|3412,3419|false|false|false|C1995603|PURPOSE (pharmacologic preparation)|purpose
Drug|Pharmacologic Substance|General Exam|3412,3419|false|false|false|C1995603|PURPOSE (pharmacologic preparation)|purpose
Event|Event|General Exam|3412,3419|false|false|false|||purpose
Finding|Functional Concept|General Exam|3412,3419|false|false|false|C1285529|Purpose|purpose
Drug|Food|General Exam|3420,3426|false|false|false|C5890763||PULSES
Event|Event|General Exam|3420,3426|false|false|false|||PULSES
Finding|Physiologic Function|General Exam|3420,3426|false|false|false|C0391850|Physiologic pulse|PULSES
Procedure|Health Care Activity|General Exam|3420,3426|false|false|false|C0034107|Pulse taking|PULSES
Drug|Food|General Exam|3434,3440|false|false|false|C5890763||pulses
Event|Event|General Exam|3434,3440|false|false|false|||pulses
Finding|Physiologic Function|General Exam|3434,3440|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|3434,3440|false|false|false|C0034107|Pulse taking|pulses
Event|Event|General Exam|3472,3478|false|false|false|||intact
Finding|Finding|General Exam|3472,3478|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Molecular Function|General Exam|3480,3484|false|false|false|C1817552|abscisic aldehyde oxidase activity|AAO3
Event|Event|General Exam|3489,3497|false|false|false|||asterxis
Anatomy|Body System|General Exam|3500,3504|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|General Exam|3500,3504|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|General Exam|3500,3504|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|General Exam|3500,3504|false|false|false|||SKIN
Finding|Body Substance|General Exam|3500,3504|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|General Exam|3500,3504|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Event|Event|General Exam|3506,3510|false|false|false|||warm
Finding|Finding|General Exam|3506,3510|false|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|General Exam|3506,3510|false|false|false|C0687712|warming process|warm
Finding|Finding|General Exam|3515,3519|false|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|3520,3528|false|false|false|||perfused
Disorder|Injury or Poisoning|General Exam|3533,3545|true|false|false|C0015256|Excoriation|excoriations
Event|Event|General Exam|3533,3545|false|false|false|||excoriations
Event|Event|General Exam|3549,3556|false|false|false|||lesions
Finding|Finding|General Exam|3549,3556|true|false|false|C0221198|Lesion|lesions
Event|Event|General Exam|3562,3568|false|false|false|||rashes
Finding|Sign or Symptom|General Exam|3562,3568|false|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Procedure|Health Care Activity|General Exam|3590,3599|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|General Exam|3600,3604|false|false|false|||LABS
Lab|Laboratory or Test Result|General Exam|3600,3604|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|General Exam|3632,3637|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3632,3637|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3632,3637|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|3638,3641|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|3647,3650|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|3647,3650|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|3647,3650|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|3657,3660|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|3657,3660|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|3657,3660|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|3657,3660|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|3666,3669|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|3666,3669|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|3676,3679|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|3676,3679|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|3676,3679|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|3676,3679|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|3676,3679|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|3685,3688|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|3685,3688|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|3685,3688|false|false|false|||MCH
Finding|Gene or Genome|General Exam|3685,3688|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|3685,3688|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|3685,3688|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|3695,3699|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|3715,3718|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|3735,3740|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3735,3740|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3735,3740|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|3745,3748|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|General Exam|3745,3748|false|false|false|||PTT
Procedure|Laboratory Procedure|General Exam|3745,3748|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|General Exam|3770,3775|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3770,3775|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3770,3775|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|3770,3783|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|3770,3783|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|3770,3783|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|3776,3783|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|3776,3783|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|3776,3783|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|3776,3783|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|3776,3783|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|3776,3783|false|false|false|C0337438|Glucose measurement|Glucose
Event|Event|General Exam|3820,3821|false|false|false|||5
Drug|Inorganic Chemical|General Exam|3831,3835|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|3831,3835|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|3831,3835|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|3860,3865|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3860,3865|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|3866,3869|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|3866,3869|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|General Exam|3866,3869|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|General Exam|3866,3869|false|false|false|||ALT
Finding|Gene or Genome|General Exam|3866,3869|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|General Exam|3866,3869|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|General Exam|3866,3869|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|General Exam|3866,3869|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|General Exam|3875,3878|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|General Exam|3875,3878|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|3875,3878|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|General Exam|3875,3878|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|General Exam|3875,3878|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|General Exam|3875,3878|false|false|false|||AST
Finding|Gene or Genome|General Exam|3875,3878|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|3884,3891|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|General Exam|3884,3891|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|General Exam|3922,3927|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3922,3927|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3922,3927|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|3922,3935|false|false|false|C0853248|Blood albumin|BLOOD Albumin
Drug|Amino Acid, Peptide, or Protein|General Exam|3928,3935|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Biologically Active Substance|General Exam|3928,3935|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Pharmacologic Substance|General Exam|3928,3935|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Event|Event|General Exam|3928,3935|false|false|false|||Albumin
Finding|Gene or Genome|General Exam|3928,3935|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Finding|Physiologic Function|General Exam|3928,3935|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Procedure|Laboratory Procedure|General Exam|3928,3935|false|false|false|C0201838|Albumin measurement|Albumin
Drug|Biologically Active Substance|General Exam|3940,3947|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|3940,3947|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|3940,3947|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|3940,3947|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|3940,3947|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|General Exam|3940,3947|false|false|false|||Calcium
Finding|Physiologic Function|General Exam|3940,3947|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|3940,3947|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|General Exam|3981,3986|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3981,3986|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3981,3986|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|3981,3994|false|false|false|C3824990|lactate in blood (lab test)|BLOOD Lactate
Drug|Organic Chemical|General Exam|3987,3994|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Drug|Pharmacologic Substance|General Exam|3987,3994|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Procedure|Laboratory Procedure|General Exam|3987,3994|false|false|false|C0202115|Lactic acid measurement|Lactate
Lab|Laboratory or Test Result|General Exam|4009,4013|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|General Exam|4039,4046|false|false|false|C0003962|Ascites|ASCITES
Event|Event|General Exam|4039,4046|false|false|false|||ASCITES
Finding|Pathologic Function|General Exam|4039,4046|false|false|false|C5441966|Peritoneal Effusion|ASCITES
Anatomy|Cell|General Exam|4047,4050|false|false|false|C0023516|Leukocytes|WBC
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|4060,4065|false|false|false|C0032400;C0071360|5'-Inosinic acid, 2'-deoxy-2'-fluoro-, homopolymer;Poly A|Polys
Event|Event|General Exam|4071,4077|false|false|false|||Lymphs
Finding|Body Substance|General Exam|4071,4077|false|false|false|C0024202|Lymph|Lymphs
Drug|Antibiotic|General Exam|4082,4087|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|General Exam|4082,4087|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|General Exam|4082,4087|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|General Exam|4136,4143|false|false|false|C0003962|Ascites|ASCITES
Event|Event|General Exam|4136,4143|false|false|false|||ASCITES
Finding|Pathologic Function|General Exam|4136,4143|false|false|false|C5441966|Peritoneal Effusion|ASCITES
Drug|Biologically Active Substance|General Exam|4155,4162|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|4155,4162|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|4155,4162|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|4155,4162|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|4155,4162|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|4155,4162|false|false|false|C0337438|Glucose measurement|Glucose
Event|Event|General Exam|4168,4180|false|false|false|||MICROBIOLOGY
Finding|Functional Concept|General Exam|4168,4180|false|false|false|C0025953;C1571921;C4049106|Microbiological;Microbiology - Laboratory Class;Microbiology Diagnostic Service Section ID|MICROBIOLOGY
Finding|Intellectual Product|General Exam|4168,4180|false|false|false|C0025953;C1571921;C4049106|Microbiological;Microbiology - Laboratory Class;Microbiology Diagnostic Service Section ID|MICROBIOLOGY
Procedure|Laboratory Procedure|General Exam|4168,4180|false|false|false|C0085672|Microbiology procedure|MICROBIOLOGY
Anatomy|Body Location or Region|General Exam|4207,4217|false|false|false|C0031153;C0442034|Peritoneum;peritoneal|PERITONEAL
Anatomy|Tissue|General Exam|4207,4217|false|false|false|C0031153;C0442034|Peritoneum;peritoneal|PERITONEAL
Finding|Body Substance|General Exam|4207,4223|false|false|false|C0003964|Peritoneal fluid (substance)|PERITONEAL FLUID
Procedure|Laboratory Procedure|General Exam|4207,4223|false|false|false|C2053903|Peritoneal fluid analysis|PERITONEAL FLUID
Drug|Substance|General Exam|4218,4223|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|FLUID
Event|Event|General Exam|4218,4223|false|false|false|||FLUID
Finding|Intellectual Product|General Exam|4218,4223|false|false|false|C1546638|Fluid Specimen Code|FLUID
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|4228,4238|false|false|false|C0061856|Gram's stain|GRAM STAIN
Drug|Organic Chemical|General Exam|4228,4238|false|false|false|C0061856|Gram's stain|GRAM STAIN
Procedure|Laboratory Procedure|General Exam|4228,4238|false|false|false|C0200966|Bacterial stain, routine|GRAM STAIN
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|4233,4238|false|false|false|C0038128|Stains|STAIN
Event|Event|General Exam|4233,4238|false|false|false|||STAIN
Procedure|Laboratory Procedure|General Exam|4233,4238|false|false|false|C0487602|Staining method|STAIN
Finding|Idea or Concept|General Exam|4240,4245|false|false|false|C1546485|Diagnosis Type - Final|Final
Anatomy|Cell|General Exam|4261,4289|false|false|false|C0018183;C0027950|granulocyte;neutrophil|POLYMORPHONUCLEAR LEUKOCYTES
Anatomy|Cell|General Exam|4279,4289|false|false|false|C0023516|Leukocytes|LEUKOCYTES
Finding|Body Substance|General Exam|4279,4289|true|false|false|C1547962;C1550647|Specimen Type - Leukocytes|LEUKOCYTES
Finding|Intellectual Product|General Exam|4279,4289|true|false|false|C1547962;C1550647|Specimen Type - Leukocytes|LEUKOCYTES
Event|Event|General Exam|4290,4294|false|false|false|||SEEN
Finding|Finding|General Exam|4306,4325|false|false|false|C2924473|Microorganisms seen|MICROORGANISMS SEEN
Event|Event|General Exam|4321,4325|false|false|false|||SEEN
Drug|Substance|General Exam|4332,4337|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|FLUID
Event|Event|General Exam|4332,4337|false|false|false|||FLUID
Finding|Intellectual Product|General Exam|4332,4337|false|false|false|C1546638|Fluid Specimen Code|FLUID
Drug|Biomedical or Dental Material|General Exam|4338,4345|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|General Exam|4338,4345|false|false|false|||CULTURE
Finding|Functional Concept|General Exam|4338,4345|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|General Exam|4338,4345|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|General Exam|4338,4345|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|General Exam|4347,4352|false|false|false|||Final
Finding|Idea or Concept|General Exam|4347,4352|false|false|false|C1546485|Diagnosis Type - Final|Final
Event|Event|General Exam|4364,4370|false|false|false|||GROWTH
Finding|Finding|General Exam|4364,4370|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organ or Tissue Function|General Exam|4364,4370|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organism Function|General Exam|4364,4370|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Physiologic Function|General Exam|4364,4370|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Phenomenon|Phenomenon or Process|General Exam|4364,4370|true|false|false|C2911660|Growth action|GROWTH
Procedure|Laboratory Procedure|General Exam|4377,4394|false|false|false|C1273935|Anaerobic microbial culture|ANAEROBIC CULTURE
Drug|Biomedical or Dental Material|General Exam|4387,4394|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|General Exam|4387,4394|false|false|false|||CULTURE
Finding|Functional Concept|General Exam|4387,4394|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|General Exam|4387,4394|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|General Exam|4387,4394|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|General Exam|4416,4422|false|false|false|||GROWTH
Finding|Finding|General Exam|4416,4422|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organ or Tissue Function|General Exam|4416,4422|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organism Function|General Exam|4416,4422|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Physiologic Function|General Exam|4416,4422|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Phenomenon|Phenomenon or Process|General Exam|4416,4422|true|false|false|C2911660|Growth action|GROWTH
Event|Event|General Exam|4433,4439|false|false|false|||screen
Procedure|Diagnostic Procedure|General Exam|4433,4439|false|false|false|C0199230;C0220908;C0430054;C1710031|Disease Screening;Screening for cancer;Screening procedure;Toxicology screen, general (procedure)|screen
Procedure|Laboratory Procedure|General Exam|4433,4439|false|false|false|C0199230;C0220908;C0430054;C1710031|Disease Screening;Screening for cancer;Screening procedure;Toxicology screen, general (procedure)|screen
Event|Event|General Exam|4444,4447|false|false|false|||VRE
Event|Event|General Exam|4448,4456|false|false|false|||isolated
Event|Event|General Exam|4459,4466|false|false|false|||IMAGING
Finding|Finding|General Exam|4459,4466|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|General Exam|4459,4466|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Event|Event|General Exam|4467,4474|false|false|false|||STUDIES
Procedure|Research Activity|General Exam|4467,4474|false|false|false|C0947630|Scientific Study|STUDIES
Event|Event|General Exam|4491,4494|false|false|false|||CXR
Procedure|Diagnostic Procedure|General Exam|4491,4494|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Intellectual Product|General Exam|4502,4507|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Location or Region|General Exam|4508,4523|false|false|false|C0553534|Cardiopulmonary|cardiopulmonary
Disorder|Disease or Syndrome|General Exam|4508,4523|false|false|false|C4072686|Cardiovascular disease+Pulmonary disease|cardiopulmonary
Anatomy|Body Part, Organ, or Organ Component|General Exam|4524,4531|false|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|General Exam|4524,4531|true|false|false|C1951340|Process Pharmacologic Substance|process
Event|Event|General Exam|4524,4531|false|false|false|||process
Finding|Functional Concept|General Exam|4524,4531|true|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|General Exam|4524,4531|true|false|false|C1522240|Process|process
Finding|Intellectual Product|General Exam|4555,4559|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Finding|General Exam|4555,4572|false|false|false|C1865190|Mild splenomegaly|mild splenomegaly
Event|Event|General Exam|4560,4572|false|false|false|||splenomegaly
Finding|Finding|General Exam|4560,4572|false|false|false|C0038002|Splenomegaly|splenomegaly
Disorder|Disease or Syndrome|General Exam|4577,4584|false|false|false|C0003962|Ascites|ascites
Event|Event|General Exam|4577,4584|false|false|false|||ascites
Finding|Pathologic Function|General Exam|4577,4584|false|false|false|C5441966|Peritoneal Effusion|ascites
Drug|Biomedical or Dental Material|General Exam|4589,4594|false|false|false|C0302909;C1378566|Solid Dose Form;solid substance|solid
Drug|Substance|General Exam|4589,4594|false|false|false|C0302909;C1378566|Solid Dose Form;solid substance|solid
Finding|Functional Concept|General Exam|4614,4618|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|General Exam|4614,4636|false|false|false|C0227486|Left lobe of liver|left lobe of the liver
Anatomy|Body Part, Organ, or Organ Component|General Exam|4619,4623|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|General Exam|4619,4623|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Anatomy|Body Part, Organ, or Organ Component|General Exam|4631,4636|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|General Exam|4631,4636|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|General Exam|4631,4636|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|General Exam|4631,4636|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|General Exam|4631,4636|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|General Exam|4631,4636|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|General Exam|4631,4636|false|false|false|||liver
Finding|Finding|General Exam|4631,4636|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|General Exam|4631,4636|false|false|false|C0872387|Procedures on liver|liver
Event|Event|General Exam|4640,4646|false|false|false|||stable
Finding|Intellectual Product|General Exam|4640,4646|false|false|false|C1547311|Patient Condition Code - Stable|stable
Attribute|Clinical Attribute|General Exam|4659,4669|false|false|false|C0550215||appearance
Event|Event|General Exam|4659,4669|false|false|false|||appearance
Procedure|Health Care Activity|General Exam|4659,4669|false|false|false|C2051406|patient appearance regarding mental status exam|appearance
Finding|Body Substance|General Exam|4673,4682|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|4673,4682|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|4673,4682|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|4673,4682|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|General Exam|4683,4687|false|false|false|||LABS
Lab|Laboratory or Test Result|General Exam|4683,4687|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|General Exam|4715,4720|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4715,4720|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4715,4720|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|4721,4724|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|4729,4732|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|4729,4732|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|4729,4732|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|4739,4742|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|4739,4742|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|4739,4742|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|4739,4742|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|4749,4752|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|4749,4752|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|4760,4763|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|4760,4763|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|4760,4763|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|4760,4763|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|4760,4763|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|4769,4772|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|4769,4772|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|4769,4772|false|false|false|||MCH
Finding|Gene or Genome|General Exam|4769,4772|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|4769,4772|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|4769,4772|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|4779,4783|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|4799,4802|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|4819,4824|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4819,4824|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4819,4824|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|4829,4832|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|General Exam|4829,4832|false|false|false|||PTT
Procedure|Laboratory Procedure|General Exam|4829,4832|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|General Exam|4854,4859|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4854,4859|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4854,4859|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|4854,4867|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|4854,4867|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|4854,4867|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|4860,4867|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|4860,4867|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|4860,4867|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|4860,4867|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|4860,4867|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|4860,4867|false|false|false|C0337438|Glucose measurement|Glucose
Event|Event|General Exam|4902,4903|false|false|false|||5
Drug|Inorganic Chemical|General Exam|4914,4918|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|4914,4918|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|4914,4918|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|4943,4948|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4943,4948|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4943,4948|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|4949,4952|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|4949,4952|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|General Exam|4949,4952|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|General Exam|4949,4952|false|false|false|||ALT
Finding|Gene or Genome|General Exam|4949,4952|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|General Exam|4949,4952|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|General Exam|4949,4952|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|General Exam|4949,4952|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|General Exam|4958,4961|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|General Exam|4958,4961|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|4958,4961|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|General Exam|4958,4961|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|General Exam|4958,4961|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Finding|Gene or Genome|General Exam|4958,4961|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|4967,4974|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|General Exam|4967,4974|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|General Exam|5005,5010|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|5005,5010|false|false|false|||BLOOD
Finding|Body Substance|General Exam|5005,5010|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|5005,5018|false|false|false|C0853248|Blood albumin|BLOOD Albumin
Drug|Amino Acid, Peptide, or Protein|General Exam|5011,5018|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Biologically Active Substance|General Exam|5011,5018|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Pharmacologic Substance|General Exam|5011,5018|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Event|Event|General Exam|5011,5018|false|false|false|||Albumin
Finding|Gene or Genome|General Exam|5011,5018|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Finding|Physiologic Function|General Exam|5011,5018|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Procedure|Laboratory Procedure|General Exam|5011,5018|false|false|false|C0201838|Albumin measurement|Albumin
Drug|Biologically Active Substance|General Exam|5023,5030|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|5023,5030|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|5023,5030|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|5023,5030|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|5023,5030|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|General Exam|5023,5030|false|false|false|||Calcium
Finding|Physiologic Function|General Exam|5023,5030|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|5023,5030|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|General Exam|5056,5059|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Disorder|Virus|General Exam|5056,5059|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Drug|Immunologic Factor|General Exam|5056,5059|false|false|false|C0086413|HIV Vaccine|HIV
Drug|Pharmacologic Substance|General Exam|5056,5059|false|false|false|C0086413|HIV Vaccine|HIV
Event|Event|General Exam|5056,5059|false|false|false|||HIV
Event|Event|General Exam|5063,5068|false|false|false|||HAART
Procedure|Therapeutic or Preventive Procedure|General Exam|5063,5068|false|false|false|C0887947|Antiretroviral Therapy, Highly Active|HAART
Disorder|Disease or Syndrome|General Exam|5070,5074|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|General Exam|5070,5074|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|General Exam|5070,5074|false|false|false|||COPD
Finding|Gene or Genome|General Exam|5070,5074|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|General Exam|5081,5085|false|false|false|||home
Finding|Idea or Concept|General Exam|5081,5085|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|General Exam|5081,5085|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|General Exam|5081,5085|false|false|false|C1553498|home health encounter|home
Disorder|Disease or Syndrome|General Exam|5090,5093|false|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|HCV
Disorder|Virus|General Exam|5090,5093|false|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|HCV
Disorder|Disease or Syndrome|General Exam|5094,5103|false|false|false|C0023890;C1623038|Cirrhosis;Liver Cirrhosis|cirrhosis
Event|Event|General Exam|5094,5103|false|false|false|||cirrhosis
Disorder|Disease or Syndrome|General Exam|5120,5127|false|false|false|C0003962|Ascites|ascites
Event|Event|General Exam|5120,5127|false|false|false|||ascites
Finding|Pathologic Function|General Exam|5120,5127|false|false|false|C5441966|Peritoneal Effusion|ascites
Event|Event|General Exam|5128,5137|false|false|false|||requiring
Drug|Organic Chemical|General Exam|5147,5158|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Drug|Pharmacologic Substance|General Exam|5147,5158|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Event|Event|General Exam|5147,5158|false|false|false|||therapeutic
Finding|Functional Concept|General Exam|5147,5158|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Finding|Intellectual Product|General Exam|5147,5158|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Procedure|Therapeutic or Preventive Procedure|General Exam|5147,5158|false|false|false|C0087111|Therapeutic procedure|therapeutic
Event|Event|General Exam|5160,5172|false|false|false|||paracenteses
Procedure|Therapeutic or Preventive Procedure|General Exam|5160,5172|false|false|false|C0034115|Paracentesis|paracenteses
Anatomy|Body Location or Region|General Exam|5174,5181|false|false|false|C0205054|Hepatic|hepatic
Disorder|Disease or Syndrome|General Exam|5174,5196|false|false|false|C0019151|Hepatic Encephalopathy|hepatic encephalopathy
Disorder|Disease or Syndrome|General Exam|5182,5196|false|false|false|C0085584|Encephalopathies|encephalopathy
Event|Event|General Exam|5182,5196|false|false|false|||encephalopathy
Anatomy|Tissue|General Exam|5205,5215|false|false|false|C0332835|Transplanted tissue|transplant
Finding|Finding|General Exam|5205,5215|false|false|false|C0478647;C3841811|Transplant;Transplanted organ and tissue status|transplant
Procedure|Therapeutic or Preventive Procedure|General Exam|5205,5215|false|false|false|C0040732|Transplantation|transplant
Event|Event|General Exam|5216,5220|false|false|false|||list
Finding|Intellectual Product|General Exam|5216,5220|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|General Exam|5228,5241|false|false|false|||comorbidities
Finding|Finding|General Exam|5228,5241|false|false|false|C0009488|Comorbidity|comorbidities
Anatomy|Body Location or Region|General Exam|5257,5260|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|abd
Disorder|Cell or Molecular Dysfunction|General Exam|5257,5260|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|abd
Attribute|Clinical Attribute|General Exam|5271,5275|false|false|false|C2598155||pain
Event|Event|General Exam|5271,5275|false|false|false|||pain
Finding|Functional Concept|General Exam|5271,5275|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|General Exam|5271,5275|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|General Exam|5280,5285|false|false|false|C2979882||Goals
Event|Event|General Exam|5280,5285|false|false|false|||Goals
Finding|Idea or Concept|General Exam|5280,5285|false|false|false|C0018017;C0679840;C1546459|What subject filter - Goals;objective (goal);treatment goals|Goals
Finding|Intellectual Product|General Exam|5280,5285|false|false|false|C0018017;C0679840;C1546459|What subject filter - Goals;objective (goal);treatment goals|Goals
Procedure|Health Care Activity|General Exam|5280,5293|false|false|false|C2930505|Goals of Care|Goals of care
Event|Activity|General Exam|5289,5293|false|false|false|C1947933|care activity|care
Event|Event|General Exam|5289,5293|false|false|false|||care
Finding|Finding|General Exam|5289,5293|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|General Exam|5289,5293|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Body Substance|General Exam|5300,5307|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|General Exam|5300,5307|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|General Exam|5300,5307|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|General Exam|5308,5317|false|false|false|||expressed
Finding|Mental Process|General Exam|5327,5333|false|false|false|C0871633|desire|desire
Event|Event|General Exam|5343,5345|false|false|false|||go
Finding|Idea or Concept|General Exam|5357,5362|false|false|false|C0680443|peace|peace
Event|Event|General Exam|5371,5376|false|false|false|||tired
Finding|Finding|General Exam|5371,5376|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Finding|Intellectual Product|General Exam|5371,5376|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Finding|Sign or Symptom|General Exam|5371,5376|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Event|Event|General Exam|5381,5389|false|false|false|||fighting
Finding|Social Behavior|General Exam|5381,5389|false|false|false|C0424324|Fighting|fighting
Drug|Amino Acid, Peptide, or Protein|General Exam|5395,5398|false|false|false|C0082420|Endoglin, human|end
Drug|Immunologic Factor|General Exam|5395,5398|false|false|false|C0082420|Endoglin, human|end
Finding|Functional Concept|General Exam|5395,5398|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Finding|Gene or Genome|General Exam|5395,5398|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Attribute|Clinical Attribute|General Exam|5399,5404|false|false|false|C1300072|Tumor stage|stage
Event|Event|General Exam|5399,5404|false|false|false|||stage
Anatomy|Body Part, Organ, or Organ Component|General Exam|5406,5411|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|General Exam|5406,5411|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|General Exam|5406,5411|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|General Exam|5406,5411|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|General Exam|5406,5411|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|General Exam|5406,5411|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|General Exam|5406,5411|false|false|false|||liver
Finding|Finding|General Exam|5406,5411|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|General Exam|5406,5411|false|false|false|C0872387|Procedures on liver|liver
Disorder|Disease or Syndrome|General Exam|5406,5419|false|false|false|C0023895;C0267792|Hepatobiliary Disorder;Liver diseases|liver disease
Disorder|Disease or Syndrome|General Exam|5412,5419|false|false|false|C0012634|Disease|disease
Event|Event|General Exam|5412,5419|false|false|false|||disease
Event|Event|General Exam|5433,5437|false|false|false|||feel
Finding|Idea or Concept|General Exam|5453,5457|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Event|Event|General Exam|5458,5465|false|false|false|||quality
Event|Event|General Exam|5470,5474|false|false|false|||life
Finding|Idea or Concept|General Exam|5470,5474|false|false|false|C0376558|Life|life
Procedure|Diagnostic Procedure|General Exam|5470,5474|false|false|false|C1522684|Laser-Induced Fluorescence Endoscopy|life
Event|Event|General Exam|5480,5486|false|false|false|||wished
Event|Event|General Exam|5490,5494|false|false|false|||meet
Event|Activity|General Exam|5502,5516|false|false|false|C1882932|Representation (action)|representative
Event|Event|General Exam|5522,5529|false|false|false|||hospice
Procedure|Health Care Activity|General Exam|5522,5529|false|false|false|C0085555|Hospice Care|hospice
Event|Event|General Exam|5546,5550|false|false|false|||able
Finding|Finding|General Exam|5546,5550|false|false|false|C1299581|Able (qualifier value)|able
Event|Event|General Exam|5554,5561|false|false|false|||arrange
Event|Event|General Exam|5571,5578|false|false|false|||decided
Event|Event|General Exam|5606,5610|false|false|false|||home
Finding|Idea or Concept|General Exam|5606,5610|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|General Exam|5606,5610|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|General Exam|5606,5610|false|false|false|C1553498|home health encounter|home
Event|Event|General Exam|5616,5623|false|false|false|||hospice
Procedure|Health Care Activity|General Exam|5616,5623|false|false|false|C0085555|Hospice Care|hospice
Event|Event|General Exam|5627,5639|false|false|false|||conversation
Finding|Social Behavior|General Exam|5627,5639|false|false|false|C0871703|conversation|conversation
Event|Event|General Exam|5644,5648|false|false|false|||held
Finding|Body Substance|General Exam|5659,5666|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|General Exam|5659,5666|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|General Exam|5659,5666|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Occupational Activity|General Exam|5677,5681|false|false|false|C0009219|Coding|code
Finding|Intellectual Product|General Exam|5677,5681|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|code
Procedure|Health Care Activity|General Exam|5677,5688|false|false|false|C0742531|CODE STATUS|code status
Attribute|Clinical Attribute|General Exam|5682,5688|false|false|false|C5889824||status
Event|Event|General Exam|5682,5688|false|false|false|||status
Finding|Idea or Concept|General Exam|5682,5688|false|false|false|C1546481|What subject filter - Status|status
Event|Event|General Exam|5694,5699|false|false|false|||noted
Finding|Finding|General Exam|5715,5723|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|probably
Finding|Idea or Concept|General Exam|5715,5723|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|probably
Attribute|Clinical Attribute|General Exam|5728,5731|false|false|false|C4285234||DNR
Drug|Antibiotic|General Exam|5728,5731|false|false|false|C0011015|daunorubicin|DNR
Drug|Organic Chemical|General Exam|5728,5731|false|false|false|C0011015|daunorubicin|DNR
Event|Event|General Exam|5728,5731|false|false|false|||DNR
Finding|Finding|General Exam|5728,5731|false|false|false|C0079252;C0582114|Do not resuscitate status;Do-Not-Resuscitate Orders|DNR
Finding|Intellectual Product|General Exam|5728,5731|false|false|false|C0079252;C0582114|Do not resuscitate status;Do-Not-Resuscitate Orders|DNR
Event|Event|General Exam|5732,5735|false|false|false|||DNI
Event|Event|General Exam|5755,5762|false|false|false|||discuss
Finding|Gene or Genome|General Exam|5775,5778|false|false|true|C1420310|SON gene|son
Disorder|Disease or Syndrome|General Exam|5780,5783|false|false|true|C0162531|Hereditary Coproporphyria|HCP
Event|Event|General Exam|5780,5783|false|false|false|||HCP
Finding|Gene or Genome|General Exam|5780,5783|false|false|true|C1335283;C1412376;C1413681;C1705637;C5780748|AMBP gene;AMBP wt Allele;CPOX gene;PTPN6 gene;PTPN6 wt Allele|HCP
Finding|Finding|General Exam|5806,5810|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|General Exam|5806,5810|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|General Exam|5806,5810|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|General Exam|5816,5823|false|false|false|||remains
Event|Event|General Exam|5829,5833|false|false|false|||code
Event|Occupational Activity|General Exam|5829,5833|false|false|false|C0009219|Coding|code
Finding|Intellectual Product|General Exam|5829,5833|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|code
Event|Event|General Exam|5844,5853|false|false|false|||discussed
Event|Event|General Exam|5858,5869|false|false|false|||possibility
Event|Event|General Exam|5895,5903|false|false|false|||catheter
Finding|Intellectual Product|General Exam|5895,5903|false|false|true|C1546572||catheter
Event|Event|General Exam|5905,5911|false|false|false|||placed
Event|Event|General Exam|5936,5948|false|false|false|||paracenteses
Procedure|Therapeutic or Preventive Procedure|General Exam|5936,5948|false|false|false|C0034115|Paracentesis|paracenteses
Event|Event|General Exam|5958,5968|false|false|false|||discharged
Event|Event|General Exam|5973,5977|false|false|false|||home
Finding|Idea or Concept|General Exam|5973,5977|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|General Exam|5973,5977|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|General Exam|5973,5977|false|false|false|C1553498|home health encounter|home
Event|Event|General Exam|5983,5990|false|false|false|||hospice
Procedure|Health Care Activity|General Exam|5983,5990|false|false|false|C0085555|Hospice Care|hospice
Disorder|Disease or Syndrome|General Exam|6016,6019|false|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|HCV
Disorder|Virus|General Exam|6016,6019|false|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|HCV
Event|Event|General Exam|6016,6019|false|false|false|||HCV
Disorder|Disease or Syndrome|General Exam|6020,6029|false|false|false|C0023890;C1623038|Cirrhosis;Liver Cirrhosis|cirrhosis
Event|Event|General Exam|6020,6029|false|false|false|||cirrhosis
Disorder|Disease or Syndrome|General Exam|6035,6042|false|false|false|C0003962|Ascites|ascites
Event|Event|General Exam|6035,6042|false|false|false|||ascites
Finding|Pathologic Function|General Exam|6035,6042|false|false|false|C5441966|Peritoneal Effusion|ascites
Finding|Body Substance|General Exam|6048,6055|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|General Exam|6048,6055|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|General Exam|6048,6055|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|General Exam|6057,6066|false|false|false|||presented
Finding|Idea or Concept|General Exam|6057,6066|false|false|false|C0449450|Presentation|presented
Finding|Idea or Concept|General Exam|6072,6081|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Disorder|Disease or Syndrome|General Exam|6082,6089|false|false|false|C0003962|Ascites|ascites
Event|Event|General Exam|6082,6089|false|false|false|||ascites
Finding|Pathologic Function|General Exam|6082,6089|false|false|false|C5441966|Peritoneal Effusion|ascites
Attribute|Clinical Attribute|General Exam|6095,6099|false|false|false|C2598155||pain
Event|Event|General Exam|6095,6099|false|false|false|||pain
Finding|Functional Concept|General Exam|6095,6099|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|General Exam|6095,6099|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|General Exam|6114,6121|false|false|false|||managed
Drug|Organic Chemical|General Exam|6128,6136|false|false|false|C0040610|tramadol|tramadol
Drug|Pharmacologic Substance|General Exam|6128,6136|false|false|false|C0040610|tramadol|tramadol
Event|Event|General Exam|6128,6136|false|false|false|||tramadol
Procedure|Laboratory Procedure|General Exam|6128,6136|false|false|false|C1266765|Tramadol measurement (procedure)|tramadol
Drug|Organic Chemical|General Exam|6141,6149|false|false|false|C0026549|morphine|morphine
Drug|Pharmacologic Substance|General Exam|6141,6149|false|false|false|C0026549|morphine|morphine
Event|Event|General Exam|6141,6149|false|false|false|||morphine
Event|Event|General Exam|6169,6181|false|false|false|||paracentesis
Procedure|Therapeutic or Preventive Procedure|General Exam|6169,6181|false|false|false|C0034115|Paracentesis|paracentesis
Event|Activity|General Exam|6195,6202|false|false|false|C1883720|Removing (action)|removal
Event|Event|General Exam|6195,6202|false|false|false|||removal
Procedure|Therapeutic or Preventive Procedure|General Exam|6195,6202|false|false|false|C0015252;C0185115;C0728940|Excision;Extraction;removal technique|removal
Drug|Amino Acid, Peptide, or Protein|General Exam|6228,6235|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Drug|Biologically Active Substance|General Exam|6228,6235|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Drug|Pharmacologic Substance|General Exam|6228,6235|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Event|Event|General Exam|6228,6235|false|false|false|||albumin
Finding|Gene or Genome|General Exam|6228,6235|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|albumin
Finding|Physiologic Function|General Exam|6228,6235|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|albumin
Procedure|Laboratory Procedure|General Exam|6228,6235|false|false|false|C0201838|Albumin measurement|albumin
Event|Event|General Exam|6237,6244|false|false|false|||Studies
Procedure|Research Activity|General Exam|6237,6244|false|false|false|C0947630|Scientific Study|Studies
Drug|Substance|General Exam|6253,6258|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|General Exam|6253,6258|false|false|false|||fluid
Finding|Intellectual Product|General Exam|6253,6258|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|General Exam|6264,6272|false|false|false|||negative
Finding|Classification|General Exam|6264,6272|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|General Exam|6264,6272|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|General Exam|6264,6272|false|false|false|C5237010|Expression Negative|negative
Event|Event|General Exam|6282,6290|false|false|false|||reported
Event|Event|General Exam|6293,6304|false|false|false|||significant
Finding|Idea or Concept|General Exam|6293,6304|false|false|false|C0750502|Significant|significant
Event|Event|General Exam|6306,6317|false|false|false|||improvement
Finding|Conceptual Entity|General Exam|6306,6317|false|false|false|C2986411|Improvement|improvement
Attribute|Clinical Attribute|General Exam|6325,6329|false|false|false|C2598155||pain
Event|Event|General Exam|6325,6329|false|false|false|||pain
Finding|Functional Concept|General Exam|6325,6329|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|General Exam|6325,6329|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|General Exam|6335,6347|false|false|false|||Hyperkalemia
Finding|Finding|General Exam|6335,6347|false|false|false|C0020461;C5700154|Hyperkalemia;Serum potassium level above reference range|Hyperkalemia
Event|Event|General Exam|6360,6375|false|false|false|||hospitalization
Procedure|Health Care Activity|General Exam|6360,6375|false|false|false|C0019993|Hospitalization|hospitalization
Event|Event|General Exam|6384,6389|false|false|false|||noted
Event|Event|General Exam|6404,6416|false|false|false|||hyperkalemia
Finding|Finding|General Exam|6404,6416|false|false|false|C0020461;C5700154|Hyperkalemia;Serum potassium level above reference range|hyperkalemia
Event|Event|General Exam|6443,6446|false|false|false|||EKG
Finding|Intellectual Product|General Exam|6443,6446|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|General Exam|6443,6446|false|false|false|C1623258|Electrocardiography|EKG
Event|Event|General Exam|6447,6454|false|false|false|||changes
Finding|Functional Concept|General Exam|6447,6454|true|false|false|C0392747|Changing|changes
Procedure|Health Care Activity|General Exam|6457,6472|false|false|false|C0001758|Aftercare|After treatment
Event|Event|General Exam|6463,6472|false|false|false|||treatment
Finding|Conceptual Entity|General Exam|6463,6472|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|General Exam|6463,6472|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|General Exam|6463,6472|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|General Exam|6463,6472|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Drug|Biologically Active Substance|General Exam|6478,6485|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Element, Ion, or Isotope|General Exam|6478,6485|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Inorganic Chemical|General Exam|6478,6485|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Pharmacologic Substance|General Exam|6478,6485|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Vitamin|General Exam|6478,6485|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Event|Event|General Exam|6478,6485|false|false|false|||calcium
Finding|Physiologic Function|General Exam|6478,6485|false|false|false|C4553026|Calcium metabolic function|calcium
Procedure|Laboratory Procedure|General Exam|6478,6485|false|false|false|C0201925|Calcium measurement|calcium
Drug|Organic Chemical|General Exam|6478,6495|false|false|false|C0006699|calcium gluconate|calcium gluconate
Drug|Pharmacologic Substance|General Exam|6478,6495|false|false|false|C0006699|calcium gluconate|calcium gluconate
Drug|Biologically Active Substance|General Exam|6486,6495|false|false|false|C0017714;C0220836|Gluconates;gluconate|gluconate
Drug|Organic Chemical|General Exam|6486,6495|false|false|false|C0017714;C0220836|Gluconates;gluconate|gluconate
Drug|Pharmacologic Substance|General Exam|6486,6495|false|false|false|C0017714;C0220836|Gluconates;gluconate|gluconate
Event|Event|General Exam|6496,6499|false|false|false|||2gm
Drug|Amino Acid, Peptide, or Protein|General Exam|6504,6511|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|General Exam|6504,6511|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|General Exam|6504,6511|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|General Exam|6504,6511|false|false|false|||insulin
Finding|Gene or Genome|General Exam|6504,6511|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|General Exam|6504,6511|false|false|false|C0202098|Insulin measurement|insulin
Event|Event|General Exam|6530,6540|false|false|false|||kayexelate
Event|Event|General Exam|6548,6559|false|false|false|||downtrended
Finding|Idea or Concept|General Exam|6584,6596|false|false|false|C0750508|persistently|persistently
Event|Event|General Exam|6597,6605|false|false|false|||elevated
Event|Event|General Exam|6629,6637|false|false|false|||continue
Event|Event|General Exam|6645,6654|false|false|false|||monitored
Anatomy|Body Location or Region|General Exam|6659,6666|false|false|false|C0205054|Hepatic|Hepatic
Disorder|Disease or Syndrome|General Exam|6659,6681|false|false|false|C0019151|Hepatic Encephalopathy|Hepatic encephalopathy
Disorder|Disease or Syndrome|General Exam|6667,6681|false|false|false|C0085584|Encephalopathies|encephalopathy
Event|Event|General Exam|6667,6681|false|false|false|||encephalopathy
Finding|Body Substance|General Exam|6687,6694|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|General Exam|6687,6694|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|General Exam|6687,6694|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Mental Process|General Exam|6697,6703|false|false|false|C0229992|Psyche structure|mental
Attribute|Clinical Attribute|General Exam|6697,6710|false|false|false|C0488568;C0488569||mental status
Finding|Finding|General Exam|6697,6710|false|false|false|C0278060|Mental state|mental status
Attribute|Clinical Attribute|General Exam|6704,6710|false|false|false|C5889824||status
Event|Event|General Exam|6704,6710|false|false|false|||status
Finding|Idea or Concept|General Exam|6704,6710|false|false|false|C1546481|What subject filter - Status|status
Event|Event|General Exam|6725,6734|false|false|false|||admission
Procedure|Health Care Activity|General Exam|6725,6734|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|General Exam|6744,6753|false|false|false|||continued
Drug|Organic Chemical|General Exam|6757,6766|false|false|false|C0073374|rifaximin|rifaximin
Drug|Pharmacologic Substance|General Exam|6757,6766|false|false|false|C0073374|rifaximin|rifaximin
Event|Event|General Exam|6757,6766|false|false|false|||rifaximin
Drug|Organic Chemical|General Exam|6771,6780|false|false|false|C0022957|lactulose|lactulose
Drug|Pharmacologic Substance|General Exam|6771,6780|false|false|false|C0022957|lactulose|lactulose
Event|Event|General Exam|6771,6780|false|false|false|||lactulose
Finding|Idea or Concept|General Exam|6782,6790|false|false|false|C4288901|In-House|in-house
Event|Event|General Exam|6798,6807|false|false|false|||discharge
Finding|Body Substance|General Exam|6798,6807|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|General Exam|6798,6807|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|General Exam|6798,6807|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|General Exam|6798,6807|false|false|false|C0030685|Patient Discharge|discharge
Finding|Intellectual Product|General Exam|6810,6817|false|false|false|C1547296|Chronic - Admission Level of Care Code|CHRONIC
Procedure|Health Care Activity|General Exam|6810,6817|false|false|false|C1555457|Provision of recurring care for chronic illness|CHRONIC
Disorder|Disease or Syndrome|General Exam|6843,6855|false|false|false|C0020625|Hyponatremia|Hyponatremia
Finding|Body Substance|General Exam|6862,6869|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|General Exam|6862,6869|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|General Exam|6862,6869|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|General Exam|6862,6873|false|false|false|C0332310|Has patient|patient has
Event|Event|General Exam|6876,6883|false|false|false|||history
Finding|Conceptual Entity|General Exam|6876,6883|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|General Exam|6876,6883|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|General Exam|6876,6883|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|General Exam|6876,6886|false|false|false|C0262926|Medical History|history of
Event|Event|General Exam|6887,6899|false|false|false|||asymptomatic
Finding|Finding|General Exam|6887,6899|false|false|false|C0231221;C0332151|Asymptomatic (finding);Asymptomatic diagnosis of|asymptomatic
Disorder|Disease or Syndrome|General Exam|6901,6913|false|false|false|C0020625|Hyponatremia|hyponatremia
Event|Event|General Exam|6901,6913|false|false|false|||hyponatremia
Finding|Idea or Concept|General Exam|6921,6932|false|false|false|C0750501|most likely|most likely
Finding|Finding|General Exam|6926,6932|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|General Exam|6926,6932|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Disorder|Disease or Syndrome|General Exam|6946,6958|false|true|false|C0020625|Hyponatremia|hyponatremia
Event|Event|General Exam|6946,6958|false|false|false|||hyponatremia
Drug|Organic Chemical|General Exam|6960,6967|false|false|false|C0163712|Relate - vinyl resin|related
Event|Event|General Exam|6960,6967|false|false|false|||related
Finding|Finding|General Exam|6960,6967|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|General Exam|6960,6967|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Event|Event|General Exam|6971,6981|false|false|false|||underlying
Anatomy|Body Part, Organ, or Organ Component|General Exam|6982,6987|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|General Exam|6982,6987|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|General Exam|6982,6987|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|General Exam|6982,6987|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|General Exam|6982,6987|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|General Exam|6982,6987|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Finding|Finding|General Exam|6982,6987|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|General Exam|6982,6987|false|false|false|C0872387|Procedures on liver|liver
Disorder|Disease or Syndrome|General Exam|6982,6995|false|false|false|C0023895;C0267792|Hepatobiliary Disorder;Liver diseases|liver disease
Disorder|Disease or Syndrome|General Exam|6988,6995|false|false|false|C0012634|Disease|disease
Event|Event|General Exam|6988,6995|false|false|false|||disease
Finding|Finding|General Exam|6999,7003|false|false|false|C5575035|Well (answer to question)|well
Drug|Hormone|General Exam|7007,7018|false|false|false|C0002006|aldosterone|aldosterone
Drug|Organic Chemical|General Exam|7007,7018|false|false|false|C0002006|aldosterone|aldosterone
Drug|Pharmacologic Substance|General Exam|7007,7018|false|false|false|C0002006|aldosterone|aldosterone
Event|Event|General Exam|7007,7018|false|false|false|||aldosterone
Procedure|Laboratory Procedure|General Exam|7007,7018|false|false|false|C0373535|Aldosterone measurement|aldosterone
Anatomy|Body Part, Organ, or Organ Component|General Exam|7019,7023|false|false|false|C0004457|Axis vertebra|axis
Disorder|Injury or Poisoning|General Exam|7019,7023|false|false|false|C0349013|Fracture of second cervical vertebra|axis
Disorder|Disease or Syndrome|General Exam|7025,7036|false|true|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Event|Event|General Exam|7025,7036|false|false|false|||dysfunction
Finding|Conceptual Entity|General Exam|7025,7036|false|true|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|General Exam|7025,7036|false|true|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|General Exam|7025,7036|false|true|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Drug|Organic Chemical|General Exam|7037,7044|false|false|false|C0163712|Relate - vinyl resin|related
Event|Event|General Exam|7037,7044|false|false|false|||related
Finding|Finding|General Exam|7037,7044|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|General Exam|7037,7044|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Anatomy|Body Part, Organ, or Organ Component|General Exam|7048,7053|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|General Exam|7048,7053|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|General Exam|7048,7053|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|General Exam|7048,7053|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|General Exam|7048,7053|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|General Exam|7048,7053|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|General Exam|7048,7053|false|false|false|||liver
Finding|Finding|General Exam|7048,7053|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|General Exam|7048,7053|false|false|false|C0872387|Procedures on liver|liver
Disorder|Disease or Syndrome|General Exam|7048,7061|false|false|false|C0023895;C0267792|Hepatobiliary Disorder;Liver diseases|liver disease
Disorder|Disease or Syndrome|General Exam|7054,7061|false|false|false|C0012634|Disease|disease
Event|Event|General Exam|7054,7061|false|false|false|||disease
Event|Event|General Exam|7067,7075|false|false|false|||remained
Event|Event|General Exam|7076,7088|false|false|false|||asymptomatic
Finding|Finding|General Exam|7076,7088|false|false|false|C0231221;C0332151|Asymptomatic (finding);Asymptomatic diagnosis of|asymptomatic
Event|Event|General Exam|7102,7117|false|false|false|||hospitalization
Procedure|Health Care Activity|General Exam|7102,7117|false|false|false|C0019993|Hospitalization|hospitalization
Event|Event|General Exam|7140,7147|false|false|false|||started
Drug|Organic Chemical|General Exam|7160,7170|false|false|false|C0016860|furosemide|furosemide
Drug|Pharmacologic Substance|General Exam|7160,7170|false|false|false|C0016860|furosemide|furosemide
Event|Event|General Exam|7160,7170|false|false|false|||furosemide
Event|Event|General Exam|7174,7178|false|false|false|||help
Event|Event|General Exam|7179,7186|false|false|false|||prevent
Drug|Substance|General Exam|7187,7192|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|General Exam|7187,7192|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|General Exam|7193,7208|false|false|false|||re-accumulation
Event|Event|General Exam|7220,7227|false|false|false|||require
Finding|Classification|General Exam|7253,7263|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|General Exam|7253,7263|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|General Exam|7264,7271|false|false|false|||setting
Finding|Mental Process|General Exam|7264,7271|false|false|false|C0542559|contextual factors|setting
Disorder|Disease or Syndrome|General Exam|7276,7279|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Disorder|Virus|General Exam|7276,7279|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Drug|Immunologic Factor|General Exam|7276,7279|false|false|false|C0086413|HIV Vaccine|HIV
Drug|Pharmacologic Substance|General Exam|7276,7279|false|false|false|C0086413|HIV Vaccine|HIV
Event|Event|General Exam|7276,7279|false|false|false|||HIV
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|7281,7294|false|false|false|C0909839|emtricitabine|Emtricitabine
Drug|Pharmacologic Substance|General Exam|7281,7294|false|false|false|C0909839|emtricitabine|Emtricitabine
Drug|Organic Chemical|General Exam|7281,7304|false|false|false|C1532298|Emtricitabine- and tenofovir-containing product|Emtricitabine-Tenofovir
Drug|Pharmacologic Substance|General Exam|7281,7304|false|false|false|C1532298|Emtricitabine- and tenofovir-containing product|Emtricitabine-Tenofovir
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|7295,7304|false|false|false|C0384228|tenofovir|Tenofovir
Drug|Pharmacologic Substance|General Exam|7295,7304|false|false|false|C0384228|tenofovir|Tenofovir
Event|Event|General Exam|7295,7304|false|false|false|||Tenofovir
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|7306,7313|false|false|false|C1528494|Truvada|Truvada
Drug|Pharmacologic Substance|General Exam|7306,7313|false|false|false|C1528494|Truvada|Truvada
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|7319,7330|false|false|false|C1871526|raltegravir|Raltegravir
Drug|Pharmacologic Substance|General Exam|7319,7330|false|false|false|C1871526|raltegravir|Raltegravir
Event|Event|General Exam|7319,7330|false|false|false|||Raltegravir
Event|Event|General Exam|7337,7346|false|false|false|||continued
Finding|Idea or Concept|General Exam|7347,7355|false|false|false|C4288901|In-House|in-house
Event|Event|General Exam|7350,7355|false|false|false|||house
Event|Event|General Exam|7363,7372|false|false|false|||discharge
Finding|Body Substance|General Exam|7363,7372|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|General Exam|7363,7372|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|General Exam|7363,7372|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|General Exam|7363,7372|false|false|false|C0030685|Patient Discharge|discharge
Disorder|Disease or Syndrome|General Exam|7379,7383|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|General Exam|7379,7383|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|General Exam|7379,7383|false|false|false|||COPD
Finding|Gene or Genome|General Exam|7379,7383|false|false|false|C1412502|ARCN1 gene|COPD
Drug|Organic Chemical|General Exam|7385,7396|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|General Exam|7385,7396|false|false|false|C0082607|fluticasone|fluticasone
Event|Event|General Exam|7385,7396|false|false|false|||fluticasone
Drug|Organic Chemical|General Exam|7398,7408|false|false|false|C0213771|tiotropium|tiotropium
Drug|Pharmacologic Substance|General Exam|7398,7408|false|false|false|C0213771|tiotropium|tiotropium
Event|Event|General Exam|7398,7408|false|false|false|||tiotropium
Drug|Organic Chemical|General Exam|7413,7422|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|General Exam|7413,7422|false|false|false|C0001927|albuterol|albuterol
Event|Event|General Exam|7413,7422|false|false|false|||albuterol
Event|Event|General Exam|7428,7437|false|false|false|||continued
Finding|Idea or Concept|General Exam|7439,7447|false|false|false|C4288901|In-House|in-house
Event|Event|General Exam|7455,7464|false|false|false|||discharge
Finding|Body Substance|General Exam|7455,7464|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|General Exam|7455,7464|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|General Exam|7455,7464|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|General Exam|7455,7464|false|false|false|C0030685|Patient Discharge|discharge
Finding|Idea or Concept|General Exam|7467,7479|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Event|Event|General Exam|7511,7517|false|false|false|||Follow
Anatomy|Body Location or Region|General Exam|7521,7531|false|false|false|C0031153;C0442034|Peritoneum;peritoneal|peritoneal
Anatomy|Tissue|General Exam|7521,7531|false|false|false|C0031153;C0442034|Peritoneum;peritoneal|peritoneal
Finding|Body Substance|General Exam|7521,7537|false|false|false|C0003964|Peritoneal fluid (substance)|peritoneal fluid
Procedure|Laboratory Procedure|General Exam|7521,7537|false|false|false|C2053903|Peritoneal fluid analysis|peritoneal fluid
Procedure|Laboratory Procedure|General Exam|7521,7545|false|false|false|C1254423|Peritoneal Fluid Culture|peritoneal fluid culture
Drug|Substance|General Exam|7532,7537|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|General Exam|7532,7537|false|false|false|C1546638|Fluid Specimen Code|fluid
Drug|Biomedical or Dental Material|General Exam|7538,7545|false|false|false|C1706355|Culture Dose Form|culture
Event|Event|General Exam|7538,7545|false|false|false|||culture
Finding|Functional Concept|General Exam|7538,7545|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Finding|Idea or Concept|General Exam|7538,7545|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Procedure|Laboratory Procedure|General Exam|7538,7545|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|culture
Finding|Finding|General Exam|7550,7553|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Finding|Idea or Concept|General Exam|7550,7553|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Attribute|Clinical Attribute|General Exam|7562,7573|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|General Exam|7562,7573|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|General Exam|7562,7573|false|false|false|||medications
Finding|Intellectual Product|General Exam|7562,7573|false|false|false|C4284232|Medications|medications
Drug|Organic Chemical|General Exam|7575,7585|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|General Exam|7575,7585|false|false|false|C0016860|furosemide|Furosemide
Finding|Finding|General Exam|7598,7601|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|General Exam|7598,7601|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Event|Event|General Exam|7611,7623|false|false|false|||hyperkalemia
Finding|Finding|General Exam|7611,7623|false|false|false|C0020461;C5700154|Hyperkalemia;Serum potassium level above reference range|hyperkalemia
Disorder|Disease or Syndrome|General Exam|7628,7640|false|false|false|C0020625|Hyponatremia|hyponatremia
Event|Event|General Exam|7628,7640|false|false|false|||hyponatremia
Finding|Body Substance|General Exam|7646,7653|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|General Exam|7646,7653|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|General Exam|7646,7653|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|General Exam|7682,7688|false|false|false|C0871893|Script|script
Event|Event|General Exam|7689,7696|false|false|false|||written
Event|Event|General Exam|7725,7730|false|false|false|||given
Finding|Intellectual Product|General Exam|7743,7747|false|false|false|C1720092|Once - dosing instruction fragment|once
Finding|Gene or Genome|General Exam|7756,7759|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|Lab
Finding|Intellectual Product|General Exam|7756,7759|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|Lab
Finding|Intellectual Product|General Exam|7756,7767|false|false|false|C3244125|lab results|Lab results
Event|Event|General Exam|7760,7767|false|false|false|||results
Event|Event|General Exam|7776,7781|false|false|false|||faxed
Finding|Functional Concept|General Exam|7782,7786|false|false|false|C1519246|Send (transmission)|sent
Event|Event|General Exam|7804,7812|false|false|false|||Continue
Event|Event|General Exam|7813,7825|false|false|false|||conversation
Finding|Social Behavior|General Exam|7813,7825|false|false|false|C0871703|conversation|conversation
Finding|Intellectual Product|General Exam|7844,7852|false|false|false|C1546572||catheter
Procedure|Therapeutic or Preventive Procedure|General Exam|7844,7862|false|false|false|C0883301|Catheter placement|catheter placement
Event|Event|General Exam|7853,7862|false|false|false|||placement
Procedure|Health Care Activity|General Exam|7853,7862|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|General Exam|7853,7862|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Event|Occupational Activity|General Exam|7868,7872|false|false|false|C0009219|Coding|code
Finding|Intellectual Product|General Exam|7868,7872|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|code
Procedure|Health Care Activity|General Exam|7868,7879|false|false|false|C0742531|CODE STATUS|code status
Attribute|Clinical Attribute|General Exam|7873,7879|false|false|false|C5889824||status
Event|Event|General Exam|7873,7879|false|false|false|||status
Finding|Idea or Concept|General Exam|7873,7879|false|false|false|C1546481|What subject filter - Status|status
Event|Event|General Exam|7894,7902|false|false|false|||continue
Event|Event|General Exam|7924,7936|false|false|false|||paracenteses
Procedure|Therapeutic or Preventive Procedure|General Exam|7924,7936|false|false|false|C0034115|Paracentesis|paracenteses
Event|Event|General Exam|7940,7944|false|false|false|||Code
Event|Occupational Activity|General Exam|7940,7944|false|false|false|C0009219|Coding|Code
Finding|Intellectual Product|General Exam|7940,7944|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|Code
Event|Event|General Exam|7955,7964|false|false|false|||Emergency
Finding|Finding|General Exam|7955,7964|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Idea or Concept|General Exam|7955,7964|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Intellectual Product|General Exam|7955,7964|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Pathologic Function|General Exam|7955,7964|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Phenomenon|Phenomenon or Process|General Exam|7955,7964|false|false|false|C0013956|Emergency Situation|Emergency
Procedure|Health Care Activity|General Exam|7955,7964|false|false|false|C1553500|emergency encounter|Emergency
Finding|Functional Concept|General Exam|7955,7972|false|false|false|C1552023|emergency contact|Emergency Contact
Event|Activity|General Exam|7965,7972|false|false|false|C3812666|Personal Contact|Contact
Finding|Functional Concept|General Exam|7965,7972|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|Contact
Finding|Idea or Concept|General Exam|7965,7972|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|Contact
Finding|Intellectual Product|General Exam|7965,7972|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|Contact
Phenomenon|Phenomenon or Process|General Exam|7965,7972|false|false|false|C0392367|Physical contact|Contact
Procedure|Health Care Activity|General Exam|7992,8001|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|General Exam|8020,8030|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|General Exam|8020,8030|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|General Exam|8020,8035|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|General Exam|8031,8035|false|false|false|||list
Finding|Intellectual Product|General Exam|8031,8035|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|General Exam|8039,8047|false|false|false|||accurate
Drug|Organic Chemical|General Exam|8052,8060|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|General Exam|8052,8060|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|General Exam|8052,8060|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|General Exam|8052,8060|false|false|false|||complete
Finding|Functional Concept|General Exam|8052,8060|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|General Exam|8052,8060|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Biologically Active Substance|General Exam|8065,8072|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|8065,8072|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|8065,8072|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|8065,8072|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|8065,8072|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|General Exam|8065,8072|false|false|false|||Calcium
Finding|Physiologic Function|General Exam|8065,8072|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|8065,8072|false|false|false|C0201925|Calcium measurement|Calcium
Drug|Inorganic Chemical|General Exam|8065,8082|false|false|false|C0006681|calcium carbonate|Calcium Carbonate
Drug|Pharmacologic Substance|General Exam|8065,8082|false|false|false|C0006681|calcium carbonate|Calcium Carbonate
Drug|Element, Ion, or Isotope|General Exam|8073,8082|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|Carbonate
Drug|Organic Chemical|General Exam|8073,8082|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|Carbonate
Drug|Pharmacologic Substance|General Exam|8073,8082|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|Carbonate
Disorder|Mental or Behavioral Dysfunction|General Exam|8093,8096|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|General Exam|8093,8096|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|General Exam|8093,8096|false|false|false|C1530795|BID protein, human|BID
Event|Event|General Exam|8093,8096|false|false|false|||BID
Finding|Gene or Genome|General Exam|8093,8096|false|false|false|C1332410|BID gene|BID
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|8101,8114|false|false|false|C0909839|emtricitabine|Emtricitabine
Drug|Pharmacologic Substance|General Exam|8101,8114|false|false|false|C0909839|emtricitabine|Emtricitabine
Drug|Organic Chemical|General Exam|8101,8124|false|false|false|C1532298|Emtricitabine- and tenofovir-containing product|Emtricitabine-Tenofovir
Drug|Pharmacologic Substance|General Exam|8101,8124|false|false|false|C1532298|Emtricitabine- and tenofovir-containing product|Emtricitabine-Tenofovir
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|8115,8124|false|false|false|C0384228|tenofovir|Tenofovir
Drug|Pharmacologic Substance|General Exam|8115,8124|false|false|false|C0384228|tenofovir|Tenofovir
Event|Event|General Exam|8115,8124|false|false|false|||Tenofovir
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|8126,8133|false|false|false|C1528494|Truvada|Truvada
Drug|Pharmacologic Substance|General Exam|8126,8133|false|false|false|C1528494|Truvada|Truvada
Drug|Biomedical or Dental Material|General Exam|8137,8140|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|General Exam|8137,8140|false|false|false|||TAB
Drug|Organic Chemical|General Exam|8154,8165|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|General Exam|8154,8165|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|General Exam|8154,8165|false|false|false|||Fluticasone
Drug|Organic Chemical|General Exam|8154,8176|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|General Exam|8154,8176|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|General Exam|8166,8176|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Event|Event|General Exam|8186,8190|false|false|false|||PUFF
Disorder|Mental or Behavioral Dysfunction|General Exam|8194,8197|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|General Exam|8194,8197|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|General Exam|8194,8197|false|false|false|C1530795|BID protein, human|BID
Event|Event|General Exam|8194,8197|false|false|false|||BID
Finding|Gene or Genome|General Exam|8194,8197|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|General Exam|8202,8211|false|false|false|C0022957|lactulose|Lactulose
Drug|Pharmacologic Substance|General Exam|8202,8211|false|false|false|C0022957|lactulose|Lactulose
Event|Event|General Exam|8202,8211|false|false|false|||Lactulose
Event|Event|General Exam|8221,8224|false|false|false|||TID
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|8229,8240|false|false|false|C1871526|raltegravir|Raltegravir
Drug|Pharmacologic Substance|General Exam|8229,8240|false|false|false|C1871526|raltegravir|Raltegravir
Disorder|Mental or Behavioral Dysfunction|General Exam|8251,8254|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|General Exam|8251,8254|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|General Exam|8251,8254|false|false|false|C1530795|BID protein, human|BID
Event|Event|General Exam|8251,8254|false|false|false|||BID
Finding|Gene or Genome|General Exam|8251,8254|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|General Exam|8259,8268|false|false|false|C0073374|rifaximin|Rifaximin
Drug|Pharmacologic Substance|General Exam|8259,8268|false|false|false|C0073374|rifaximin|Rifaximin
Disorder|Mental or Behavioral Dysfunction|General Exam|8279,8282|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|General Exam|8279,8282|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|General Exam|8279,8282|false|false|false|C1530795|BID protein, human|BID
Event|Event|General Exam|8279,8282|false|false|false|||BID
Finding|Gene or Genome|General Exam|8279,8282|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|General Exam|8287,8295|false|false|false|C0040610|tramadol|TraMADOL
Drug|Pharmacologic Substance|General Exam|8287,8295|false|false|false|C0040610|tramadol|TraMADOL
Event|Event|General Exam|8287,8295|false|false|false|||TraMADOL
Procedure|Laboratory Procedure|General Exam|8287,8295|false|false|false|C1266765|Tramadol measurement (procedure)|TraMADOL
Drug|Organic Chemical|General Exam|8297,8303|false|false|false|C0724054|Ultram|Ultram
Drug|Pharmacologic Substance|General Exam|8297,8303|false|false|false|C0724054|Ultram|Ultram
Finding|Gene or Genome|General Exam|8319,8322|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|General Exam|8323,8327|false|false|false|C2598155||pain
Event|Event|General Exam|8323,8327|false|false|false|||pain
Finding|Functional Concept|General Exam|8323,8327|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|General Exam|8323,8327|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|General Exam|8332,8341|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|General Exam|8332,8341|false|false|false|C0001927|albuterol|albuterol
Event|Event|General Exam|8332,8341|false|false|false|||albuterol
Drug|Organic Chemical|General Exam|8332,8349|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|General Exam|8332,8349|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|General Exam|8342,8349|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|General Exam|8342,8349|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|General Exam|8342,8349|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Event|Event|General Exam|8342,8349|false|false|false|||sulfate
Finding|Functional Concept|General Exam|8367,8377|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Organism Function|General Exam|8367,8377|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Event|Event|General Exam|8378,8381|false|false|false|||Q6H
Finding|Gene or Genome|General Exam|8382,8385|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Sign or Symptom|General Exam|8387,8395|false|false|false|C0043144|Wheezing|Wheezing
Drug|Organic Chemical|General Exam|8400,8410|false|false|false|C0213771|tiotropium|Tiotropium
Drug|Pharmacologic Substance|General Exam|8400,8410|false|false|false|C0213771|tiotropium|Tiotropium
Event|Event|General Exam|8400,8410|false|false|false|||Tiotropium
Drug|Organic Chemical|General Exam|8400,8418|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Pharmacologic Substance|General Exam|8400,8418|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Inorganic Chemical|General Exam|8411,8418|false|false|false|C0006222|Bromides|Bromide
Event|Event|General Exam|8411,8418|false|false|false|||Bromide
Procedure|Laboratory Procedure|General Exam|8411,8418|false|false|false|C0202341|Bromides measurement|Bromide
Disorder|Congenital Abnormality|General Exam|8421,8424|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|CAP
Drug|Biomedical or Dental Material|General Exam|8421,8424|false|false|false|C0006935|capsule (pharmacologic)|CAP
Event|Event|General Exam|8421,8424|false|false|false|||CAP
Finding|Gene or Genome|General Exam|8421,8424|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|CAP
Procedure|Therapeutic or Preventive Procedure|General Exam|8421,8424|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|CAP
Event|Event|General Exam|8438,8447|false|false|false|||Discharge
Finding|Body Substance|General Exam|8438,8447|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|General Exam|8438,8447|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|General Exam|8438,8447|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|General Exam|8438,8447|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|General Exam|8438,8459|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|General Exam|8448,8459|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|General Exam|8448,8459|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|General Exam|8448,8459|false|false|false|||Medications
Finding|Intellectual Product|General Exam|8448,8459|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|General Exam|8464,8473|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|General Exam|8464,8473|false|false|false|C0001927|albuterol|albuterol
Event|Event|General Exam|8464,8473|false|false|false|||albuterol
Drug|Organic Chemical|General Exam|8464,8481|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|General Exam|8464,8481|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|General Exam|8474,8481|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|General Exam|8474,8481|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|General Exam|8474,8481|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Event|Event|General Exam|8474,8481|false|false|false|||sulfate
Finding|Functional Concept|General Exam|8499,8509|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Organism Function|General Exam|8499,8509|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Event|Event|General Exam|8510,8513|false|false|false|||Q6H
Finding|Gene or Genome|General Exam|8514,8517|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Sign or Symptom|General Exam|8519,8527|false|false|false|C0043144|Wheezing|Wheezing
Drug|Biologically Active Substance|General Exam|8532,8539|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|8532,8539|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|8532,8539|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|8532,8539|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|8532,8539|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|General Exam|8532,8539|false|false|false|||Calcium
Finding|Physiologic Function|General Exam|8532,8539|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|8532,8539|false|false|false|C0201925|Calcium measurement|Calcium
Drug|Inorganic Chemical|General Exam|8532,8549|false|false|false|C0006681|calcium carbonate|Calcium Carbonate
Drug|Pharmacologic Substance|General Exam|8532,8549|false|false|false|C0006681|calcium carbonate|Calcium Carbonate
Drug|Element, Ion, or Isotope|General Exam|8540,8549|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|Carbonate
Drug|Organic Chemical|General Exam|8540,8549|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|Carbonate
Drug|Pharmacologic Substance|General Exam|8540,8549|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|Carbonate
Disorder|Mental or Behavioral Dysfunction|General Exam|8560,8563|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|General Exam|8560,8563|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|General Exam|8560,8563|false|false|false|C1530795|BID protein, human|BID
Event|Event|General Exam|8560,8563|false|false|false|||BID
Finding|Gene or Genome|General Exam|8560,8563|false|false|false|C1332410|BID gene|BID
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|8568,8581|false|false|false|C0909839|emtricitabine|Emtricitabine
Drug|Pharmacologic Substance|General Exam|8568,8581|false|false|false|C0909839|emtricitabine|Emtricitabine
Drug|Organic Chemical|General Exam|8568,8591|false|false|false|C1532298|Emtricitabine- and tenofovir-containing product|Emtricitabine-Tenofovir
Drug|Pharmacologic Substance|General Exam|8568,8591|false|false|false|C1532298|Emtricitabine- and tenofovir-containing product|Emtricitabine-Tenofovir
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|8582,8591|false|false|false|C0384228|tenofovir|Tenofovir
Drug|Pharmacologic Substance|General Exam|8582,8591|false|false|false|C0384228|tenofovir|Tenofovir
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|8593,8600|false|false|false|C1528494|Truvada|Truvada
Drug|Pharmacologic Substance|General Exam|8593,8600|false|false|false|C1528494|Truvada|Truvada
Drug|Biomedical or Dental Material|General Exam|8604,8607|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|General Exam|8604,8607|false|false|false|||TAB
Drug|Organic Chemical|General Exam|8621,8632|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|General Exam|8621,8632|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|General Exam|8621,8632|false|false|false|||Fluticasone
Drug|Organic Chemical|General Exam|8621,8643|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|General Exam|8621,8643|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|General Exam|8633,8643|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Event|Event|General Exam|8644,8650|false|false|false|||110mcg
Event|Event|General Exam|8653,8657|false|false|false|||PUFF
Disorder|Mental or Behavioral Dysfunction|General Exam|8661,8664|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|General Exam|8661,8664|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|General Exam|8661,8664|false|false|false|C1530795|BID protein, human|BID
Event|Event|General Exam|8661,8664|false|false|false|||BID
Finding|Gene or Genome|General Exam|8661,8664|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|General Exam|8669,8678|false|false|false|C0022957|lactulose|Lactulose
Drug|Pharmacologic Substance|General Exam|8669,8678|false|false|false|C0022957|lactulose|Lactulose
Event|Event|General Exam|8688,8691|false|false|false|||TID
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|8696,8707|false|false|false|C1871526|raltegravir|Raltegravir
Drug|Pharmacologic Substance|General Exam|8696,8707|false|false|false|C1871526|raltegravir|Raltegravir
Event|Event|General Exam|8696,8707|false|false|false|||Raltegravir
Disorder|Mental or Behavioral Dysfunction|General Exam|8718,8721|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|General Exam|8718,8721|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|General Exam|8718,8721|false|false|false|C1530795|BID protein, human|BID
Event|Event|General Exam|8718,8721|false|false|false|||BID
Finding|Gene or Genome|General Exam|8718,8721|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|General Exam|8726,8735|false|false|false|C0073374|rifaximin|Rifaximin
Drug|Pharmacologic Substance|General Exam|8726,8735|false|false|false|C0073374|rifaximin|Rifaximin
Disorder|Mental or Behavioral Dysfunction|General Exam|8746,8749|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|General Exam|8746,8749|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|General Exam|8746,8749|false|false|false|C1530795|BID protein, human|BID
Event|Event|General Exam|8746,8749|false|false|false|||BID
Finding|Gene or Genome|General Exam|8746,8749|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|General Exam|8754,8764|false|false|false|C0213771|tiotropium|Tiotropium
Drug|Pharmacologic Substance|General Exam|8754,8764|false|false|false|C0213771|tiotropium|Tiotropium
Event|Event|General Exam|8754,8764|false|false|false|||Tiotropium
Drug|Organic Chemical|General Exam|8754,8772|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Pharmacologic Substance|General Exam|8754,8772|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Inorganic Chemical|General Exam|8765,8772|false|false|false|C0006222|Bromides|Bromide
Event|Event|General Exam|8765,8772|false|false|false|||Bromide
Procedure|Laboratory Procedure|General Exam|8765,8772|false|false|false|C0202341|Bromides measurement|Bromide
Disorder|Congenital Abnormality|General Exam|8775,8778|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|CAP
Drug|Biomedical or Dental Material|General Exam|8775,8778|false|false|false|C0006935|capsule (pharmacologic)|CAP
Event|Event|General Exam|8775,8778|false|false|false|||CAP
Finding|Gene or Genome|General Exam|8775,8778|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|CAP
Procedure|Therapeutic or Preventive Procedure|General Exam|8775,8778|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|CAP
Drug|Organic Chemical|General Exam|8792,8800|false|false|false|C0040610|tramadol|TraMADOL
Drug|Pharmacologic Substance|General Exam|8792,8800|false|false|false|C0040610|tramadol|TraMADOL
Event|Event|General Exam|8792,8800|false|false|false|||TraMADOL
Procedure|Laboratory Procedure|General Exam|8792,8800|false|false|false|C1266765|Tramadol measurement (procedure)|TraMADOL
Drug|Organic Chemical|General Exam|8802,8808|false|false|false|C0724054|Ultram|Ultram
Drug|Pharmacologic Substance|General Exam|8802,8808|false|false|false|C0724054|Ultram|Ultram
Finding|Gene or Genome|General Exam|8824,8827|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|General Exam|8828,8832|false|false|false|C2598155||pain
Event|Event|General Exam|8828,8832|false|false|false|||pain
Finding|Functional Concept|General Exam|8828,8832|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|General Exam|8828,8832|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|General Exam|8838,8848|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|General Exam|8838,8848|false|false|false|C0016860|furosemide|Furosemide
Drug|Organic Chemical|General Exam|8869,8879|false|false|false|C0016860|furosemide|furosemide
Drug|Pharmacologic Substance|General Exam|8869,8879|false|false|false|C0016860|furosemide|furosemide
Event|Event|General Exam|8869,8879|false|false|false|||furosemide
Drug|Biomedical or Dental Material|General Exam|8901,8907|false|false|false|C0039225|Tablet Dosage Form|tablet
Event|Event|General Exam|8901,8907|false|false|false|||tablet
Finding|Functional Concept|General Exam|8911,8919|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|General Exam|8914,8919|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|General Exam|8914,8919|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Event|General Exam|8928,8932|false|false|false|||take
Drug|Biomedical or Dental Material|General Exam|8935,8941|false|false|false|C0039225|Tablet Dosage Form|tablet
Event|Event|General Exam|8935,8941|false|false|false|||tablet
Drug|Biomedical or Dental Material|General Exam|8959,8965|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|General Exam|8966,8973|false|false|false|||Refills
Finding|Idea or Concept|General Exam|8966,8973|false|false|false|C0807726|refill|Refills
Finding|Classification|General Exam|8981,8991|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|Outpatient
Finding|Idea or Concept|General Exam|8981,8991|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|Outpatient
Finding|Gene or Genome|General Exam|8992,8995|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|Lab
Finding|Intellectual Product|General Exam|8992,8995|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|Lab
Event|Event|General Exam|8996,9000|false|false|false|||Work
Event|Occupational Activity|General Exam|8996,9000|false|false|false|C0043227|Work|Work
Drug|Amino Acid, Peptide, or Protein|General Exam|9024,9027|false|false|false|C0053932|Bone Morphogenetic Proteins|BMP
Drug|Biologically Active Substance|General Exam|9024,9027|false|false|false|C0053932|Bone Morphogenetic Proteins|BMP
Event|Event|General Exam|9024,9027|false|false|false|||BMP
Procedure|Therapeutic or Preventive Procedure|General Exam|9024,9027|false|false|false|C0279266|carmustine/methotrexate/procarbazine protocol|BMP
Event|Event|General Exam|9031,9038|false|false|false|||monitor
Event|Event|General Exam|9045,9047|false|false|false|||Na
Event|Event|General Exam|9056,9059|false|false|false|||fax
Event|Event|General Exam|9061,9068|false|false|false|||results
Event|Event|General Exam|9102,9111|false|false|false|||Discharge
Finding|Body Substance|General Exam|9102,9111|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|General Exam|9102,9111|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|General Exam|9102,9111|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|General Exam|9102,9111|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|General Exam|9102,9123|false|false|false|C4019243||Discharge Disposition
Finding|Finding|General Exam|9102,9123|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|General Exam|9112,9123|false|false|false|C2926604||Disposition
Event|Event|General Exam|9112,9123|false|false|false|||Disposition
Procedure|Health Care Activity|General Exam|9112,9123|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|General Exam|9125,9129|false|false|false|||Home
Finding|Idea or Concept|General Exam|9125,9129|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|General Exam|9125,9129|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|General Exam|9125,9129|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|General Exam|9135,9142|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|General Exam|9135,9142|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|General Exam|9145,9153|false|false|false|||Facility
Finding|Intellectual Product|General Exam|9145,9153|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|General Exam|9161,9170|false|false|false|||Discharge
Finding|Body Substance|General Exam|9161,9170|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|General Exam|9161,9170|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|General Exam|9161,9170|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|General Exam|9161,9170|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|General Exam|9161,9180|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|General Exam|9171,9180|false|false|false|C0945731||Diagnosis
Event|Event|General Exam|9171,9180|false|false|false|||Diagnosis
Finding|Classification|General Exam|9171,9180|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|General Exam|9171,9180|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|General Exam|9171,9180|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Disease or Syndrome|Principle Diagnosis|9233,9236|false|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|HCV
Disorder|Virus|Principle Diagnosis|9233,9236|false|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|HCV
Event|Event|Principle Diagnosis|9233,9236|false|false|false|||HCV
Disorder|Disease or Syndrome|Principle Diagnosis|9237,9246|false|false|false|C0023890;C1623038|Cirrhosis;Liver Cirrhosis|cirrhosis
Event|Event|Principle Diagnosis|9237,9246|false|false|false|||cirrhosis
Event|Event|Principle Diagnosis|9248,9260|false|false|false|||Hyperkalemia
Finding|Finding|Principle Diagnosis|9248,9260|false|false|false|C0020461;C5700154|Hyperkalemia;Serum potassium level above reference range|Hyperkalemia
Disorder|Neoplastic Process|Principle Diagnosis|9262,9271|false|false|false|C0027627|Neoplasm Metastasis|SECONDARY
Finding|Functional Concept|Principle Diagnosis|9262,9271|false|false|false|C1522484|metastatic qualifier|SECONDARY
Procedure|Diagnostic Procedure|Principle Diagnosis|9272,9281|false|false|false|C0011900|Diagnosis|DIAGNOSES
Disorder|Disease or Syndrome|Principle Diagnosis|9303,9306|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Disorder|Virus|Principle Diagnosis|9303,9306|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Drug|Immunologic Factor|Principle Diagnosis|9303,9306|false|false|false|C0086413|HIV Vaccine|HIV
Drug|Pharmacologic Substance|Principle Diagnosis|9303,9306|false|false|false|C0086413|HIV Vaccine|HIV
Event|Event|Principle Diagnosis|9303,9306|false|false|false|||HIV
Disorder|Disease or Syndrome|Principle Diagnosis|9308,9312|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Principle Diagnosis|9308,9312|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Principle Diagnosis|9308,9312|false|false|false|||COPD
Finding|Gene or Genome|Principle Diagnosis|9308,9312|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|Principle Diagnosis|9314,9326|false|false|false|C0020625|Hyponatremia|Hyponatremia
Event|Event|Principle Diagnosis|9314,9326|false|false|false|||Hyponatremia
Finding|Mental Process|Discharge Condition|9351,9357|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|9351,9364|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|9351,9364|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|9358,9364|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|9358,9364|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|9366,9371|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|9366,9371|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|9376,9384|false|false|false|||coherent
Finding|Finding|Discharge Condition|9376,9384|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|9386,9391|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|9386,9408|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|9386,9408|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|9395,9408|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|9395,9408|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|9395,9408|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|9410,9415|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|9410,9415|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|9410,9415|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|9410,9415|false|false|false|||Alert
Finding|Finding|Discharge Condition|9410,9415|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|9410,9415|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|9410,9415|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|9420,9431|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|9420,9431|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|9433,9441|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|9433,9441|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|9433,9441|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|9442,9448|false|false|false|C5889824||Status
Event|Event|Discharge Condition|9442,9448|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|9442,9448|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|9450,9460|false|false|false|||Ambulatory
Finding|Functional Concept|Discharge Condition|9450,9460|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|9450,9460|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|9450,9460|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|9450,9460|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|9463,9474|false|false|false|||Independent
Finding|Finding|Discharge Condition|9463,9474|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Condition|9463,9474|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Gene or Genome|Discharge Instructions|9503,9507|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|Discharge Instructions|9527,9535|false|false|false|||pleasure
Finding|Intellectual Product|Discharge Instructions|9527,9535|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|Discharge Instructions|9527,9535|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Event|Discharge Instructions|9536,9542|false|false|false|||caring
Event|Event|Discharge Instructions|9586,9594|false|false|false|||admitted
Anatomy|Body Location or Region|Discharge Instructions|9616,9625|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|Discharge Instructions|9616,9630|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|Discharge Instructions|9626,9630|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|9626,9630|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|9626,9630|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|9626,9630|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Discharge Instructions|9638,9644|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Discharge Instructions|9638,9644|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Attribute|Clinical Attribute|Discharge Instructions|9656,9660|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|9656,9660|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|9656,9660|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|9656,9660|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Substance|Discharge Instructions|9683,9688|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|Discharge Instructions|9683,9688|false|false|false|||fluid
Finding|Intellectual Product|Discharge Instructions|9683,9688|false|false|false|C1546638|Fluid Specimen Code|fluid
Anatomy|Body Location or Region|Discharge Instructions|9696,9703|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|Discharge Instructions|9696,9703|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Finding|Finding|Discharge Instructions|9696,9703|false|false|false|C0941288|Abdomen problem|abdomen
Disorder|Disease or Syndrome|Discharge Instructions|9715,9724|false|false|false|C0023890;C1623038|Cirrhosis;Liver Cirrhosis|cirrhosis
Event|Event|Discharge Instructions|9715,9724|false|false|false|||cirrhosis
Event|Event|Discharge Instructions|9734,9746|false|false|false|||paracentesis
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|9734,9746|false|false|false|C0034115|Paracentesis|paracentesis
Finding|Finding|Discharge Instructions|9756,9760|false|false|false|C4281574|Much|much
Drug|Substance|Discharge Instructions|9769,9774|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|Discharge Instructions|9769,9774|false|false|false|||fluid
Finding|Intellectual Product|Discharge Instructions|9769,9774|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|Discharge Instructions|9780,9787|false|false|false|||removed
Attribute|Clinical Attribute|Discharge Instructions|9794,9798|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|9794,9798|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|9794,9798|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|9794,9798|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Discharge Instructions|9799,9807|false|false|false|||improved
Event|Event|Discharge Instructions|9832,9837|false|false|false|||noted
Finding|Finding|Discharge Instructions|9849,9853|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|Discharge Instructions|9849,9853|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|Discharge Instructions|9849,9853|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Finding|Discharge Instructions|9849,9863|false|false|false|C0856882|Potassium increased|high potassium
Drug|Biologically Active Substance|Discharge Instructions|9854,9863|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Element, Ion, or Isotope|Discharge Instructions|9854,9863|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Food|Discharge Instructions|9854,9863|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Inorganic Chemical|Discharge Instructions|9854,9863|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Pharmacologic Substance|Discharge Instructions|9854,9863|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Event|Event|Discharge Instructions|9854,9863|false|false|false|||potassium
Finding|Physiologic Function|Discharge Instructions|9854,9863|false|false|false|C4553027|Potassium metabolic function|potassium
Procedure|Laboratory Procedure|Discharge Instructions|9854,9863|false|false|false|C0202194|Potassium measurement|potassium
Event|Event|Discharge Instructions|9876,9891|false|false|false|||hospitalization
Procedure|Health Care Activity|Discharge Instructions|9876,9891|false|false|false|C0019993|Hospitalization|hospitalization
Drug|Organic Chemical|Discharge Instructions|9899,9903|false|false|false|C0960273|CAME|came
Event|Event|Discharge Instructions|9899,9903|false|false|false|||came
Event|Event|Discharge Instructions|9915,9924|false|false|false|||treatment
Finding|Conceptual Entity|Discharge Instructions|9915,9924|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Discharge Instructions|9915,9924|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Discharge Instructions|9915,9924|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|9915,9924|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Event|Event|Discharge Instructions|9929,9933|false|false|false|||this
Event|Event|Discharge Instructions|9941,9949|false|false|false|||continue
Event|Event|Discharge Instructions|9956,9964|false|false|false|||followed
Event|Event|Discharge Instructions|9972,9982|false|false|false|||outpatient
Finding|Classification|Discharge Instructions|9972,9982|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Discharge Instructions|9972,9982|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|Discharge Instructions|9993,10003|false|false|false|||emphasized
Event|Event|Discharge Instructions|10009,10015|false|false|false|||desire
Finding|Mental Process|Discharge Instructions|10009,10015|false|false|false|C0871633|desire|desire
Event|Event|Discharge Instructions|10019,10024|false|false|false|||speak
Event|Activity|Discharge Instructions|10033,10047|false|false|false|C1882932|Representation (action)|representative
Event|Event|Discharge Instructions|10033,10047|false|false|false|||representative
Event|Event|Discharge Instructions|10053,10060|false|false|false|||hospice
Procedure|Health Care Activity|Discharge Instructions|10053,10060|false|false|false|C0085555|Hospice Care|hospice
Event|Event|Discharge Instructions|10078,10086|false|false|false|||repeated
Event|Event|Discharge Instructions|10088,10100|false|false|false|||paracenteses
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10088,10100|false|false|false|C0034115|Paracentesis|paracenteses
Event|Event|Discharge Instructions|10110,10119|false|false|false|||discussed
Event|Event|Discharge Instructions|10141,10148|false|false|false|||pleurex
Event|Event|Discharge Instructions|10150,10158|false|false|false|||catheter
Finding|Intellectual Product|Discharge Instructions|10150,10158|false|false|false|C1546572||catheter
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10150,10168|false|false|false|C0883301|Catheter placement|catheter placement
Event|Event|Discharge Instructions|10159,10168|false|false|false|||placement
Procedure|Health Care Activity|Discharge Instructions|10159,10168|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10159,10168|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Event|Event|Discharge Instructions|10173,10181|false|false|false|||arranged
Event|Event|Discharge Instructions|10193,10197|false|false|false|||meet
Event|Event|Discharge Instructions|10203,10210|false|false|false|||hospice
Procedure|Health Care Activity|Discharge Instructions|10203,10210|false|false|false|C0085555|Hospice Care|hospice
Event|Event|Discharge Instructions|10212,10224|false|false|false|||coordinators
Event|Event|Discharge Instructions|10253,10257|false|false|false|||home
Finding|Idea or Concept|Discharge Instructions|10253,10257|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Discharge Instructions|10253,10257|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Discharge Instructions|10253,10257|false|false|false|C1553498|home health encounter|home
Event|Event|Discharge Instructions|10263,10270|false|false|false|||hospice
Procedure|Health Care Activity|Discharge Instructions|10263,10270|false|false|false|C0085555|Hospice Care|hospice
Disorder|Disease or Syndrome|Discharge Instructions|10293,10297|false|false|false|C0339510|Vitelliform Macular Dystrophy|best
Event|Event|Discharge Instructions|10293,10297|false|false|false|||best
Finding|Gene or Genome|Discharge Instructions|10293,10297|false|false|false|C1826421;C5781213|BEST1 gene;BEST1 wt Allele|best
Event|Activity|Discharge Instructions|10309,10313|false|false|false|C1947933|care activity|care
Finding|Finding|Discharge Instructions|10309,10313|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|10309,10313|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Attribute|Clinical Attribute|Discharge Instructions|10309,10318|false|false|false|C4321316||care team
Finding|Finding|Discharge Instructions|10309,10318|false|false|false|C4321315|Care team|care team
Procedure|Health Care Activity|Discharge Instructions|10321,10329|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|10330,10342|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|10330,10342|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|10330,10342|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

