 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|26,30
No|31,33
:|33,34
_|37,38
_|38,39
_|39,40
<EOL>|40,41
<EOL>|42,43
Admission|43,52
Date|53,57
:|57,58
_|60,61
_|61,62
_|62,63
Discharge|77,86
Date|87,91
:|91,92
_|95,96
_|96,97
_|97,98
<EOL>|98,99
<EOL>|100,101
Date|101,105
of|106,108
Birth|109,114
:|114,115
_|117,118
_|118,119
_|119,120
Sex|133,136
:|136,137
F|140,141
<EOL>|141,142
<EOL>|143,144
Service|144,151
:|151,152
MEDICINE|153,161
<EOL>|161,162
<EOL>|163,164
No|176,178
Known|179,184
Allergies|185,194
/|195,196
Adverse|197,204
Drug|205,209
Reactions|210,219
<EOL>|219,220
<EOL>|221,222
Attending|222,231
:|231,232
_|233,234
_|234,235
_|235,236
.|236,237
<EOL>|237,238
<EOL>|239,240
subjective|257,267
fevers|268,274
,|274,275
lethargy|276,284
,|284,285
and|286,289
bloody|290,296
drain|297,302
output|303,309
<EOL>|310,311
<EOL>|312,313
Major|313,318
Surgical|319,327
or|328,330
Invasive|331,339
Procedure|340,349
:|349,350
<EOL>|350,351
_|351,352
_|352,353
_|353,354
:|354,355
For|356,359
the|360,363
large|364,369
pelvic|370,376
fluid|377,382
collections|383,394
,|394,395
CT|396,398
-|398,399
guided|399,405
<EOL>|406,407
repositioning|407,420
of|421,423
existing|424,432
drain|433,438
and|439,442
placement|443,452
of|453,455
an|456,458
additional|459,469
<EOL>|470,471
drain|471,476
.|476,477
<EOL>|477,478
<EOL>|478,479
_|479,480
_|480,481
_|481,482
:|482,483
Removal|484,491
of|492,494
more|495,499
recently|500,508
placed|509,515
drain|516,521
<EOL>|523,524
<EOL>|524,525
<EOL>|526,527
Ms.|555,558
_|559,560
_|560,561
_|561,562
is|563,565
an|566,568
_|569,570
_|570,571
_|571,572
with|573,577
PMH|578,581
of|582,584
hypertension|585,597
and|598,601
bladder|602,609
<EOL>|610,611
cancer|611,617
(|618,619
high|619,623
grade|624,629
invasive|630,638
urothelial|639,649
carcinoma|650,659
pT2b|660,664
)|664,665
s|666,667
/|667,668
p|668,669
<EOL>|670,671
TAH|671,674
/|674,675
BSO|675,678
,|678,679
radical|680,687
cystectomy|688,698
w|699,700
/|700,701
ileal|701,706
conduit|707,714
c|715,716
/|716,717
b|717,718
intra-abdominal|719,734
<EOL>|735,736
infection|736,745
and|746,749
pelvic|750,756
fluid|757,762
collection|763,773
s|774,775
/|775,776
p|776,777
_|778,779
_|779,780
_|780,781
guided|782,788
drain|789,794
<EOL>|795,796
placement|796,805
_|806,807
_|807,808
_|808,809
who|810,813
presents|814,822
with|823,827
2|828,829
days|830,834
of|835,837
generalized|838,849
<EOL>|850,851
malaise|851,858
and|859,862
1|863,864
day|865,868
of|869,871
fevers|872,878
.|878,879
<EOL>|881,882
Patient|883,890
underwent|891,900
_|901,902
_|902,903
_|903,904
guided|905,911
JP|912,914
drain|915,920
placement|921,930
for|931,934
<EOL>|935,936
intra-abdominal|936,951
fluid|952,957
collection|958,968
and|969,972
infection|973,982
,|982,983
thought|984,991
to|992,994
be|995,997
<EOL>|998,999
complicated|999,1010
of|1011,1013
recent|1014,1020
TAH|1021,1024
/|1024,1025
BSO|1025,1028
,|1028,1029
radical|1030,1037
cystectomy|1038,1048
and|1049,1052
pelvic|1053,1059
<EOL>|1060,1061
lymph|1061,1066
node|1067,1071
biopsy|1072,1078
.|1078,1079
This|1080,1084
procedure|1085,1094
was|1095,1098
done|1099,1103
on|1104,1106
_|1107,1108
_|1108,1109
_|1109,1110
.|1110,1111
Over|1112,1116
the|1117,1120
<EOL>|1121,1122
past|1122,1126
2|1127,1128
days|1129,1133
she|1134,1137
had|1138,1141
noticed|1142,1149
generalized|1150,1161
malaise|1162,1169
and|1170,1173
1|1174,1175
day|1176,1179
of|1180,1182
<EOL>|1183,1184
fever|1184,1189
w|1190,1191
/|1191,1192
rigors|1192,1198
to|1199,1201
Tmax|1202,1206
101.5|1207,1212
at|1213,1215
home|1216,1220
.|1220,1221
She|1222,1225
notes|1226,1231
that|1232,1236
the|1237,1240
<EOL>|1241,1242
drainage|1242,1250
from|1251,1255
her|1256,1259
intra-abdominal|1260,1275
drain|1276,1281
is|1282,1284
darker|1285,1291
,|1291,1292
but|1293,1296
her|1297,1300
<EOL>|1301,1302
urostomy|1302,1310
output|1311,1317
has|1318,1321
been|1322,1326
unchanged|1327,1336
.|1336,1337
She|1338,1341
notes|1342,1347
some|1348,1352
associated|1353,1363
<EOL>|1364,1365
mild|1365,1369
LLQ|1370,1373
pain|1374,1378
.|1378,1379
She|1380,1383
denies|1384,1390
diarrhea|1391,1399
,|1399,1400
BRBPR|1401,1406
,|1406,1407
rash|1408,1412
,|1412,1413
cough|1414,1419
,|1419,1420
<EOL>|1421,1422
headache|1422,1430
,|1430,1431
neck|1432,1436
stiffness|1437,1446
.|1446,1447
She|1448,1451
presented|1452,1461
initially|1462,1471
to|1472,1474
OSH|1475,1478
,|1478,1479
where|1480,1485
<EOL>|1486,1487
she|1487,1490
was|1491,1494
evaluated|1495,1504
with|1505,1509
BCx|1510,1513
and|1514,1517
drain|1518,1523
culture|1524,1531
and|1532,1535
was|1536,1539
started|1540,1547
on|1548,1550
<EOL>|1551,1552
zosyn|1552,1557
and|1558,1561
vancomycin|1562,1572
and|1573,1576
given|1577,1582
650mg|1583,1588
acetaminophen|1589,1602
.|1602,1603
She|1604,1607
was|1608,1611
<EOL>|1612,1613
transferred|1613,1624
to|1625,1627
_|1628,1629
_|1629,1630
_|1630,1631
for|1632,1635
further|1636,1643
management|1644,1654
.|1654,1655
<EOL>|1657,1658
<EOL>|1658,1659
<EOL>|1660,1661
-|1683,1684
Hypertension|1685,1697
<EOL>|1699,1700
-|1701,1702
s|1703,1704
/|1704,1705
p|1705,1706
lap|1707,1710
chole|1711,1716
<EOL>|1718,1719
-|1720,1721
s|1722,1723
/|1723,1724
p|1724,1725
left|1726,1730
knee|1731,1735
replacement|1736,1747
<EOL>|1749,1750
-|1751,1752
s|1753,1754
/|1754,1755
p|1755,1756
laminectomy|1757,1768
of|1769,1771
L5|1772,1774
-|1774,1775
S1|1775,1777
at|1778,1780
age|1781,1784
_|1785,1786
_|1786,1787
_|1787,1788
<EOL>|1790,1791
-|1792,1793
Bladder|1794,1801
Cancer|1802,1808
high|1809,1813
grade|1814,1819
TCC|1820,1823
,|1823,1824
T1|1825,1827
diagnosed|1828,1837
in|1838,1840
_|1841,1842
_|1842,1843
_|1843,1844
,|1844,1845
then|1846,1850
<EOL>|1851,1852
_|1852,1853
_|1853,1854
_|1854,1855
pelvic|1856,1862
MRI|1863,1866
w|1867,1868
/|1868,1869
invasion|1869,1877
into|1878,1882
bladder|1883,1890
wall|1891,1895
,|1895,1896
perivesical|1897,1908
<EOL>|1909,1910
soft|1910,1914
tissue|1915,1921
and|1922,1925
anterior|1926,1934
vaginal|1935,1942
wall|1943,1947
c|1948,1949
/|1949,1950
w|1950,1951
T4|1952,1954
staging|1955,1962
<EOL>|1964,1965
-|1966,1967
s|1968,1969
/|1969,1970
p|1970,1971
hysterectomy|1972,1984
and|1985,1988
bilateral|1989,1998
oophorectomy|1999,2011
for|2012,2015
large|2016,2021
uterus|2022,2028
<EOL>|2029,2030
w|2030,2031
/|2031,2032
fibroid|2032,2039
,|2039,2040
s|2041,2042
/|2042,2043
p|2043,2044
laparascopic|2045,2057
b|2058,2059
/|2059,2060
l|2060,2061
pelvic|2062,2068
lymph|2069,2074
node|2075,2079
resection|2080,2089
,|2089,2090
s|2091,2092
/|2092,2093
p|2093,2094
<EOL>|2095,2096
radical|2096,2103
cystectomy|2104,2114
and|2115,2118
anterior|2119,2127
vaginectomy|2128,2139
with|2140,2144
vaginal|2145,2152
<EOL>|2153,2154
reconstruction|2154,2168
with|2169,2173
ileal|2174,2179
conduit|2180,2187
creation|2188,2196
_|2197,2198
_|2198,2199
_|2199,2200
,|2200,2201
course|2202,2208
<EOL>|2209,2210
complicated|2210,2221
by|2222,2224
bacteremia|2225,2235
and|2236,2239
development|2240,2251
of|2252,2254
intra-abdominal|2255,2270
<EOL>|2271,2272
fluid|2272,2277
collection|2278,2288
,|2288,2289
no|2290,2292
s|2293,2294
/|2294,2295
p|2295,2296
drain|2297,2302
placement|2303,2312
by|2313,2315
_|2316,2317
_|2317,2318
_|2318,2319
_|2320,2321
_|2321,2322
_|2322,2323
<EOL>|2325,2326
-|2327,2328
h|2329,2330
/|2330,2331
o|2331,2332
LLE|2333,2336
DVT|2337,2340
and|2341,2344
PE|2345,2347
on|2348,2350
lovenox|2351,2358
<EOL>|2360,2361
<EOL>|2361,2362
<EOL>|2363,2364
:|2378,2379
<EOL>|2379,2380
_|2380,2381
_|2381,2382
_|2382,2383
<EOL>|2383,2384
:|2398,2399
<EOL>|2399,2400
Negative|2400,2408
for|2409,2412
bladder|2413,2420
CA|2421,2423
.|2423,2424
<EOL>|2424,2425
<EOL>|2425,2426
<EOL>|2427,2428
ADMISSION|2443,2452
EXAM|2453,2457
:|2457,2458
<EOL>|2458,2459
=|2459,2460
=|2460,2461
=|2461,2462
=|2462,2463
=|2463,2464
=|2464,2465
=|2465,2466
=|2466,2467
=|2467,2468
=|2468,2469
=|2469,2470
=|2470,2471
=|2471,2472
=|2472,2473
=|2473,2474
<EOL>|2474,2475
Vital|2476,2481
Signs|2482,2487
:|2487,2488
100.9|2489,2494
PO|2495,2497
130|2498,2501
/|2502,2503
54|2504,2506
L|2507,2508
Lying|2509,2514
80|2515,2517
24|2518,2520
95|2521,2523
RA|2524,2526
<EOL>|2528,2529
General|2530,2537
:|2537,2538
Alert|2539,2544
,|2544,2545
oriented|2546,2554
,|2554,2555
no|2556,2558
acute|2559,2564
distress|2565,2573
<EOL>|2575,2576
HEENT|2577,2582
:|2582,2583
Sclerae|2584,2591
anicteric|2592,2601
,|2601,2602
MMM|2603,2606
,|2606,2607
oropharynx|2608,2618
clear|2619,2624
<EOL>|2626,2627
CV|2628,2630
:|2630,2631
RRR|2632,2635
,|2635,2636
normal|2637,2643
S1|2644,2646
S2|2647,2649
,|2649,2650
systolic|2651,2659
murmur|2660,2666
RUBS|2667,2671
,|2671,2672
no|2673,2675
rubs|2676,2680
,|2680,2681
gallops|2682,2689
<EOL>|2691,2692
Lungs|2693,2698
:|2698,2699
Clear|2700,2705
to|2706,2708
auscultation|2709,2721
bilaterally|2722,2733
,|2733,2734
no|2735,2737
wheezes|2738,2745
,|2745,2746
rales|2747,2752
,|2752,2753
<EOL>|2754,2755
rhonchi|2755,2762
<EOL>|2764,2765
Abdomen|2766,2773
:|2773,2774
Soft|2775,2779
,|2779,2780
non-tender|2781,2791
,|2791,2792
non-distended|2793,2806
,|2806,2807
bowel|2808,2813
sounds|2814,2820
present|2821,2828
,|2828,2829
<EOL>|2830,2831
+|2831,2832
ileal|2832,2837
conduit|2838,2845
drain|2846,2851
in|2852,2854
RLQ|2855,2858
,|2858,2859
with|2860,2864
pigtail|2865,2872
drain|2873,2878
in|2879,2881
LLQ|2882,2885
draining|2886,2894
<EOL>|2895,2896
dark|2896,2900
/|2900,2901
sang|2901,2905
fluid|2906,2911
<EOL>|2913,2914
GU|2915,2917
:|2917,2918
No|2919,2921
foley|2922,2927
<EOL>|2929,2930
Ext|2931,2934
:|2934,2935
Warm|2936,2940
,|2940,2941
well|2942,2946
perfused|2947,2955
,|2955,2956
1|2957,2958
+|2958,2959
nonpitting|2960,2970
edema|2971,2976
LLE|2977,2980
<EOL>|2982,2983
Neuro|2984,2989
:|2989,2990
CN2|2991,2994
-|2994,2995
12|2995,2997
grossly|2998,3005
intact|3006,3012
,|3012,3013
moving|3014,3020
all|3021,3024
extremities|3025,3036
<EOL>|3037,3038
spontaneously|3038,3051
<EOL>|3051,3052
<EOL>|3052,3053
DISCHARGE|3053,3062
EXAM|3063,3067
:|3067,3068
<EOL>|3069,3070
=|3070,3071
=|3071,3072
=|3072,3073
=|3073,3074
=|3074,3075
=|3075,3076
=|3076,3077
=|3077,3078
=|3078,3079
=|3079,3080
=|3080,3081
=|3081,3082
=|3082,3083
=|3083,3084
=|3084,3085
<EOL>|3085,3086
Vital|3087,3092
signs|3093,3098
:|3098,3099
98.3|3100,3104
134|3106,3109
/|3109,3110
64|3110,3112
71|3114,3116
20|3118,3120
96|3122,3124
RA|3125,3127
<EOL>|3128,3129
General|3130,3137
:|3137,3138
AxO|3139,3142
x3|3143,3145
<EOL>|3145,3146
HEENT|3147,3152
:|3152,3153
Sclera|3154,3160
anicteric|3161,3170
<EOL>|3170,3171
Neck|3172,3176
:|3176,3177
supple|3178,3184
<EOL>|3185,3186
Lungs|3187,3192
:|3192,3193
Clear|3194,3199
to|3200,3202
auscultation|3203,3215
bilaterally|3216,3227
,|3227,3228
no|3229,3231
wheezes|3232,3239
,|3239,3240
rales|3241,3246
,|3246,3247
<EOL>|3248,3249
rhonchi|3249,3256
on|3257,3259
anterior|3260,3268
auscultation|3269,3281
<EOL>|3282,3283
CV|3284,3286
:|3286,3287
Regular|3288,3295
rate|3296,3300
and|3301,3304
rhythm|3305,3311
,|3311,3312
normal|3313,3319
S1|3320,3322
+|3323,3324
S2|3325,3327
,|3327,3328
III|3329,3332
/|3332,3333
VI|3333,3335
SEM|3336,3339
<EOL>|3339,3340
Abdomen|3341,3348
:|3348,3349
+|3350,3351
BS|3351,3353
,|3353,3354
ileal|3355,3360
conduit|3361,3368
draining|3369,3377
clear|3378,3383
yellow|3384,3390
urine|3391,3396
.|3396,3397
Has|3399,3402
<EOL>|3403,3404
one|3404,3407
LLQ|3408,3411
drain|3412,3417
in|3418,3420
place|3421,3426
draining|3427,3435
serosanguinous|3436,3450
fluid|3451,3456
.|3456,3457
<EOL>|3458,3459
Ext|3460,3463
:|3463,3464
Warm|3465,3469
,|3469,3470
well|3471,3475
perfused|3476,3484
,|3484,3485
2|3486,3487
+|3487,3488
pulses|3489,3495
,|3495,3496
no|3497,3499
clubbing|3500,3508
,|3508,3509
cyanosis|3510,3518
or|3519,3521
<EOL>|3522,3523
edema|3523,3528
<EOL>|3530,3531
<EOL>|3532,3533
Pertinent|3533,3542
Results|3543,3550
:|3550,3551
<EOL>|3551,3552
ADMISSION|3552,3561
LABS|3562,3566
:|3566,3567
<EOL>|3567,3568
=|3568,3569
=|3569,3570
=|3570,3571
=|3571,3572
=|3572,3573
=|3573,3574
=|3574,3575
=|3575,3576
=|3576,3577
=|3577,3578
=|3578,3579
=|3579,3580
=|3580,3581
=|3581,3582
=|3582,3583
<EOL>|3583,3584
_|3584,3585
_|3585,3586
_|3586,3587
07|3588,3590
:|3590,3591
10PM|3591,3595
BLOOD|3596,3601
WBC|3602,3605
-|3605,3606
19|3606,3608
.|3608,3609
4|3609,3610
*|3610,3611
#|3611,3612
RBC|3613,3616
-|3616,3617
2|3617,3618
.|3618,3619
53|3619,3621
*|3621,3622
Hgb|3623,3626
-|3626,3627
6|3627,3628
.|3628,3629
9|3629,3630
*|3630,3631
Hct|3632,3635
-|3635,3636
22|3636,3638
.|3638,3639
9|3639,3640
*|3640,3641
<EOL>|3642,3643
MCV|3643,3646
-|3646,3647
91|3647,3649
MCH|3650,3653
-|3653,3654
27.3|3654,3658
MCHC|3659,3663
-|3663,3664
30|3664,3666
.|3666,3667
1|3667,3668
*|3668,3669
RDW|3670,3673
-|3673,3674
15.1|3674,3678
RDWSD|3679,3684
-|3684,3685
49|3685,3687
.|3687,3688
5|3688,3689
*|3689,3690
Plt|3691,3694
_|3695,3696
_|3696,3697
_|3697,3698
<EOL>|3698,3699
_|3699,3700
_|3700,3701
_|3701,3702
07|3703,3705
:|3705,3706
10PM|3706,3710
BLOOD|3711,3716
Neuts|3717,3722
-|3722,3723
81|3723,3725
.|3725,3726
4|3726,3727
*|3727,3728
Lymphs|3729,3735
-|3735,3736
9|3736,3737
.|3737,3738
4|3738,3739
*|3739,3740
Monos|3741,3746
-|3746,3747
7.4|3747,3750
<EOL>|3751,3752
Eos|3752,3755
-|3755,3756
0|3756,3757
.|3757,3758
0|3758,3759
*|3759,3760
Baso|3761,3765
-|3765,3766
0.1|3766,3769
Im|3770,3772
_|3773,3774
_|3774,3775
_|3775,3776
AbsNeut|3777,3784
-|3784,3785
15|3785,3787
.|3787,3788
77|3788,3790
*|3790,3791
#|3791,3792
AbsLymp|3793,3800
-|3800,3801
1|3801,3802
.|3802,3803
81|3803,3805
<EOL>|3806,3807
AbsMono|3807,3814
-|3814,3815
1|3815,3816
.|3816,3817
43|3817,3819
*|3819,3820
AbsEos|3821,3827
-|3827,3828
0|3828,3829
.|3829,3830
00|3830,3832
*|3832,3833
AbsBaso|3834,3841
-|3841,3842
0|3842,3843
.|3843,3844
02|3844,3846
<EOL>|3846,3847
_|3847,3848
_|3848,3849
_|3849,3850
07|3851,3853
:|3853,3854
10PM|3854,3858
BLOOD|3859,3864
_|3865,3866
_|3866,3867
_|3867,3868
PTT|3869,3872
-|3872,3873
33.4|3873,3877
_|3878,3879
_|3879,3880
_|3880,3881
<EOL>|3881,3882
_|3882,3883
_|3883,3884
_|3884,3885
07|3886,3888
:|3888,3889
10PM|3889,3893
BLOOD|3894,3899
Ret|3900,3903
Aut|3904,3907
-|3907,3908
2|3908,3909
.|3909,3910
9|3910,3911
*|3911,3912
Abs|3913,3916
Ret|3917,3920
-|3920,3921
0.07|3921,3925
<EOL>|3925,3926
_|3926,3927
_|3927,3928
_|3928,3929
07|3930,3932
:|3932,3933
10PM|3933,3937
BLOOD|3938,3943
Glucose|3944,3951
-|3951,3952
118|3952,3955
*|3955,3956
UreaN|3957,3962
-|3962,3963
25|3963,3965
*|3965,3966
Creat|3967,3972
-|3972,3973
1.1|3973,3976
Na|3977,3979
-|3979,3980
133|3980,3983
<EOL>|3984,3985
K|3985,3986
-|3986,3987
5.0|3987,3990
Cl|3991,3993
-|3993,3994
97|3994,3996
HCO3|3997,4001
-|4001,4002
23|4002,4004
AnGap|4005,4010
-|4010,4011
18|4011,4013
<EOL>|4013,4014
_|4014,4015
_|4015,4016
_|4016,4017
07|4018,4020
:|4020,4021
10PM|4021,4025
BLOOD|4026,4031
ALT|4032,4035
-|4035,4036
9|4036,4037
AST|4038,4041
-|4041,4042
9|4042,4043
AlkPhos|4044,4051
-|4051,4052
56|4052,4054
TotBili|4055,4062
-|4062,4063
0.3|4063,4066
<EOL>|4066,4067
_|4067,4068
_|4068,4069
_|4069,4070
07|4071,4073
:|4073,4074
10PM|4074,4078
BLOOD|4079,4084
Lipase|4085,4091
-|4091,4092
9|4092,4093
<EOL>|4093,4094
_|4094,4095
_|4095,4096
_|4096,4097
07|4098,4100
:|4100,4101
10PM|4101,4105
BLOOD|4106,4111
Albumin|4112,4119
-|4119,4120
2|4120,4121
.|4121,4122
5|4122,4123
*|4123,4124
Iron|4125,4129
-|4129,4130
6|4130,4131
*|4131,4132
<EOL>|4132,4133
_|4133,4134
_|4134,4135
_|4135,4136
07|4137,4139
:|4139,4140
10PM|4140,4144
BLOOD|4145,4150
calTIBC|4151,4158
-|4158,4159
170|4159,4162
*|4162,4163
Hapto|4164,4169
-|4169,4170
518|4170,4173
*|4173,4174
Ferritn|4175,4182
-|4182,4183
489|4183,4186
*|4186,4187
<EOL>|4188,4189
TRF|4189,4192
-|4192,4193
131|4193,4196
*|4196,4197
<EOL>|4197,4198
_|4198,4199
_|4199,4200
_|4200,4201
07|4202,4204
:|4204,4205
13PM|4205,4209
BLOOD|4210,4215
Lactate|4216,4223
-|4223,4224
1.0|4224,4227
<EOL>|4227,4228
<EOL>|4228,4229
DISCHARGE|4229,4238
LABS|4239,4243
:|4243,4244
<EOL>|4244,4245
=|4245,4246
=|4246,4247
=|4247,4248
=|4248,4249
=|4249,4250
=|4250,4251
=|4251,4252
=|4252,4253
=|4253,4254
=|4254,4255
=|4255,4256
=|4256,4257
=|4257,4258
=|4258,4259
=|4259,4260
<EOL>|4260,4261
_|4261,4262
_|4262,4263
_|4263,4264
06|4265,4267
:|4267,4268
00AM|4268,4272
BLOOD|4273,4278
WBC|4279,4282
-|4282,4283
6.9|4283,4286
RBC|4287,4290
-|4290,4291
2|4291,4292
.|4292,4293
92|4293,4295
*|4295,4296
Hgb|4297,4300
-|4300,4301
8|4301,4302
.|4302,4303
3|4303,4304
*|4304,4305
Hct|4306,4309
-|4309,4310
26|4310,4312
.|4312,4313
8|4313,4314
*|4314,4315
<EOL>|4316,4317
MCV|4317,4320
-|4320,4321
92|4321,4323
MCH|4324,4327
-|4327,4328
28.4|4328,4332
MCHC|4333,4337
-|4337,4338
31|4338,4340
.|4340,4341
0|4341,4342
*|4342,4343
RDW|4344,4347
-|4347,4348
15.4|4348,4352
RDWSD|4353,4358
-|4358,4359
52|4359,4361
.|4361,4362
4|4362,4363
*|4363,4364
Plt|4365,4368
_|4369,4370
_|4370,4371
_|4371,4372
<EOL>|4372,4373
_|4373,4374
_|4374,4375
_|4375,4376
06|4377,4379
:|4379,4380
00AM|4380,4384
BLOOD|4385,4390
_|4391,4392
_|4392,4393
_|4393,4394
PTT|4395,4398
-|4398,4399
31.2|4399,4403
_|4404,4405
_|4405,4406
_|4406,4407
<EOL>|4407,4408
_|4408,4409
_|4409,4410
_|4410,4411
06|4412,4414
:|4414,4415
00AM|4415,4419
BLOOD|4420,4425
Plt|4426,4429
_|4430,4431
_|4431,4432
_|4432,4433
<EOL>|4433,4434
_|4434,4435
_|4435,4436
_|4436,4437
06|4438,4440
:|4440,4441
00AM|4441,4445
BLOOD|4446,4451
Glucose|4452,4459
-|4459,4460
86|4460,4462
UreaN|4463,4468
-|4468,4469
8|4469,4470
Creat|4471,4476
-|4476,4477
0.8|4477,4480
Na|4481,4483
-|4483,4484
143|4484,4487
K|4488,4489
-|4489,4490
3.6|4490,4493
<EOL>|4494,4495
Cl|4495,4497
-|4497,4498
106|4498,4501
HCO3|4502,4506
-|4506,4507
25|4507,4509
AnGap|4510,4515
-|4515,4516
16|4516,4518
<EOL>|4518,4519
_|4519,4520
_|4520,4521
_|4521,4522
06|4523,4525
:|4525,4526
00AM|4526,4530
BLOOD|4531,4536
Calcium|4537,4544
-|4544,4545
7|4545,4546
.|4546,4547
5|4547,4548
*|4548,4549
Phos|4550,4554
-|4554,4555
3.7|4555,4558
Mg|4559,4561
-|4561,4562
2.3|4562,4565
<EOL>|4565,4566
<EOL>|4566,4567
MICROBIOLOGY|4567,4579
:|4579,4580
<EOL>|4580,4581
=|4581,4582
=|4582,4583
=|4583,4584
=|4584,4585
=|4585,4586
=|4586,4587
=|4587,4588
=|4588,4589
=|4589,4590
=|4590,4591
=|4591,4592
=|4592,4593
=|4593,4594
<EOL>|4594,4595
Blood|4595,4600
cultures|4601,4609
x3|4610,4612
pending|4613,4620
<EOL>|4620,4621
<EOL>|4621,4622
_|4622,4623
_|4623,4624
_|4624,4625
4|4626,4627
:|4627,4628
35|4628,4630
pm|4631,4633
pelvic|4634,4640
aspiration|4641,4651
<EOL>|4651,4652
GRAM|4655,4659
STAIN|4660,4665
(|4666,4667
Final|4667,4672
_|4673,4674
_|4674,4675
_|4675,4676
:|4676,4677
<EOL>|4678,4679
1|4685,4686
+|4686,4687
(|4691,4692
<|4692,4693
1|4693,4694
per|4695,4698
1000X|4699,4704
FIELD|4705,4710
)|4710,4711
:|4711,4712
POLYMORPHONUCLEAR|4715,4732
<EOL>|4733,4734
LEUKOCYTES|4734,4744
.|4744,4745
<EOL>|4746,4747
NO|4753,4755
MICROORGANISMS|4756,4770
SEEN|4771,4775
.|4775,4776
<EOL>|4777,4778
FLUID|4781,4786
CULTURE|4787,4794
(|4795,4796
Final|4796,4801
_|4802,4803
_|4803,4804
_|4804,4805
:|4805,4806
NO|4810,4812
GROWTH|4813,4819
.|4819,4820
<EOL>|4821,4822
ANAEROBIC|4825,4834
CULTURE|4835,4842
(|4843,4844
Preliminary|4844,4855
)|4855,4856
:|4856,4857
NO|4861,4863
GROWTH|4864,4870
.|4870,4871
<EOL>|4872,4873
<EOL>|4873,4874
PERTINENT|4874,4883
IMAGING|4884,4891
:|4891,4892
<EOL>|4892,4893
=|4893,4894
=|4894,4895
=|4895,4896
=|4896,4897
=|4897,4898
=|4898,4899
=|4899,4900
=|4900,4901
=|4901,4902
=|4902,4903
=|4903,4904
=|4904,4905
=|4905,4906
=|4906,4907
=|4907,4908
=|4908,4909
=|4909,4910
=|4910,4911
<EOL>|4911,4912
CT|4912,4914
ABD|4915,4918
&|4918,4919
PEL|4919,4922
W|4923,4924
/|4924,4925
CONTRAST|4926,4934
<EOL>|4935,4936
_|4936,4937
_|4937,4938
_|4938,4939
<EOL>|4939,4940
1.|4940,4942
Interval|4943,4951
decrease|4952,4960
in|4961,4963
size|4964,4968
of|4969,4971
the|4972,4975
right|4976,4981
hemipelvis|4982,4992
fluid|4993,4998
<EOL>|4999,5000
collection|5000,5010
(|5011,5012
7.0|5012,5015
x|5016,5017
6.5|5018,5021
x|5022,5023
11.3|5024,5028
cm|5029,5031
,|5031,5032
previously|5033,5043
10.0|5044,5048
x|5049,5050
12.7|5051,5055
x|5056,5057
14.8|5058,5062
<EOL>|5063,5064
cm|5064,5066
)|5066,5067
with|5068,5072
the|5073,5076
anterior|5077,5085
approach|5086,5094
pigtail|5095,5102
catheter|5103,5111
unchanged|5112,5121
in|5122,5124
<EOL>|5125,5126
position|5126,5134
.|5134,5135
The|5137,5140
pigtail|5141,5148
is|5149,5151
again|5152,5157
located|5158,5165
partly|5166,5172
within|5173,5179
the|5180,5183
<EOL>|5184,5185
collection|5185,5195
and|5196,5199
partly|5200,5206
outside|5207,5214
its|5215,5218
wall|5219,5223
.|5223,5224
<EOL>|5225,5226
2.|5226,5228
Interval|5229,5237
increase|5238,5246
in|5247,5249
size|5250,5254
of|5255,5257
the|5258,5261
left|5262,5266
pelvic|5267,5273
fluid|5274,5279
<EOL>|5280,5281
collection|5281,5291
,|5291,5292
now|5293,5296
<EOL>|5297,5298
measuring|5298,5307
14.7|5308,5312
x|5313,5314
16.2|5315,5319
x|5320,5321
23.3|5322,5326
cm|5327,5329
(|5330,5331
previously|5331,5341
13.6|5342,5346
x|5347,5348
13.9|5349,5353
x|5354,5355
23.0|5356,5360
<EOL>|5361,5362
cm|5362,5364
)|5364,5365
.|5365,5366
Increased|5367,5376
peripheral|5377,5387
enhancement|5388,5399
may|5400,5403
suggest|5404,5411
superimposed|5412,5424
<EOL>|5425,5426
infection|5426,5435
.|5435,5436
<EOL>|5437,5438
3.|5438,5440
No|5441,5443
new|5444,5447
fluid|5448,5453
collection|5454,5464
identified|5465,5475
.|5475,5476
<EOL>|5477,5478
<EOL>|5480,5481
CTA|5481,5484
ABD|5485,5488
&|5489,5490
PELVIS|5491,5497
<EOL>|5497,5498
_|5498,5499
_|5499,5500
_|5500,5501
<EOL>|5501,5502
1.|5502,5504
Decrease|5505,5513
in|5514,5516
size|5517,5521
of|5522,5524
right|5525,5530
lower|5531,5536
quadrant|5537,5545
fluid|5546,5551
collection|5552,5562
<EOL>|5563,5564
that|5564,5568
has|5569,5572
<EOL>|5573,5574
percutaneous|5574,5586
drain|5587,5592
within|5593,5599
it|5600,5602
,|5602,5603
with|5604,5608
areas|5609,5614
of|5615,5617
high|5618,5622
attenuation|5623,5634
on|5635,5637
<EOL>|5638,5639
noncontrast|5639,5650
exam|5651,5655
consistent|5656,5666
with|5667,5671
blood|5672,5677
products|5678,5686
,|5686,5687
and|5688,5691
associated|5692,5702
<EOL>|5703,5704
hyperemia|5704,5713
which|5714,5719
is|5720,5722
likely|5723,5729
inflammatory|5730,5742
,|5742,5743
but|5744,5747
without|5748,5755
evidence|5756,5764
of|5765,5767
<EOL>|5768,5769
contrast|5769,5777
extravasation|5778,5791
.|5791,5792
<EOL>|5793,5794
2|5794,5795
.|5795,5796
There|5797,5802
is|5803,5805
large|5806,5811
stable|5812,5818
fluid|5819,5824
collection|5825,5835
in|5836,5838
the|5839,5842
low|5843,5846
left|5847,5851
<EOL>|5852,5853
abdomen|5853,5860
,|5860,5861
pelvis|5862,5868
with|5869,5873
mild|5874,5878
linear|5879,5885
peripheral|5886,5896
enhancement|5897,5908
,|5908,5909
<EOL>|5910,5911
infection|5911,5920
can|5921,5924
not|5924,5927
be|5928,5930
excluded|5931,5939
.|5939,5940
<EOL>|5941,5942
3|5942,5943
.|5943,5944
There|5945,5950
is|5951,5953
severe|5954,5960
left|5961,5965
,|5965,5966
and|5967,5970
moderate|5971,5979
to|5980,5982
severe|5983,5989
right|5990,5995
<EOL>|5996,5997
hydroureteronephrosis|5997,6018
,|6018,6019
with|6020,6024
delayed|6025,6032
left|6033,6037
nephrogram|6038,6048
,|6048,6049
stable|6050,6056
from|6057,6061
<EOL>|6062,6063
today|6063,6068
.|6068,6069
Mass|6071,6075
effect|6076,6082
about|6083,6088
anastomosis|6089,6100
between|6101,6108
distal|6109,6115
ureters|6116,6123
and|6124,6127
<EOL>|6128,6129
neobladder|6129,6139
has|6140,6143
resolved|6144,6152
all|6153,6156
since|6157,6162
_|6163,6164
_|6164,6165
_|6165,6166
,|6166,6167
and|6168,6171
while|6172,6177
<EOL>|6178,6179
hydronephrosis|6179,6193
may|6194,6197
be|6198,6200
from|6201,6205
residual|6206,6214
edema|6215,6220
,|6220,6221
if|6222,6224
this|6225,6229
does|6230,6234
not|6235,6238
<EOL>|6239,6240
resolve|6240,6247
,|6247,6248
alternative|6249,6260
etiologies|6261,6271
including|6272,6281
stenosis|6282,6290
,|6290,6291
tumor|6292,6297
<EOL>|6298,6299
infiltration|6299,6311
should|6312,6318
be|6319,6321
excluded|6322,6330
.|6330,6331
<EOL>|6332,6333
4.|6333,6335
Tiny|6336,6340
hepatic|6341,6348
lesion|6349,6355
segment|6356,6363
_|6364,6365
_|6365,6366
_|6366,6367
,|6367,6368
attention|6369,6378
to|6379,6381
this|6382,6386
area|6387,6391
on|6392,6394
<EOL>|6395,6396
subsequent|6396,6406
<EOL>|6407,6408
followups|6408,6417
recommended|6418,6429
.|6429,6430
<EOL>|6431,6432
<EOL>|6432,6433
CT|6433,6435
INTERVENTIONAL|6436,6450
PROCEDURE|6451,6460
<EOL>|6460,6461
_|6461,6462
_|6462,6463
_|6463,6464
<EOL>|6465,6466
1.|6466,6468
Complete|6470,6478
collapse|6479,6487
the|6488,6491
patient|6492,6499
has|6500,6503
recently|6504,6512
drained|6513,6520
left|6521,6525
<EOL>|6526,6527
lower|6527,6532
quadrant|6533,6541
<EOL>|6542,6543
collection|6543,6553
.|6553,6554
The|6556,6559
catheter|6560,6568
from|6569,6573
this|6574,6578
collection|6579,6589
was|6590,6593
removed|6594,6601
.|6601,6602
<EOL>|6603,6604
2.|6604,6606
Near|6608,6612
complete|6613,6621
collapse|6622,6630
of|6631,6633
the|6634,6637
patient|6638,6645
is|6646,6648
originally|6649,6659
drained|6660,6667
<EOL>|6668,6669
collection|6669,6679
in|6680,6682
the|6683,6686
mid|6687,6690
pelvis|6691,6697
,|6697,6698
with|6699,6703
pigtail|6704,6711
catheter|6712,6720
in|6721,6723
place|6724,6729
.|6729,6730
<EOL>|6731,6732
3.|6732,6734
Left|6736,6740
lower|6741,6746
quadrant|6747,6755
and|6756,6759
deep|6760,6764
pelvic|6765,6771
collections|6772,6783
as|6784,6786
above|6787,6792
.|6792,6793
<EOL>|6795,6796
These|6796,6801
findings|6802,6810
were|6811,6815
discussed|6816,6825
with|6826,6830
the|6831,6834
team|6835,6839
.|6839,6840
Given|6842,6847
the|6848,6851
<EOL>|6852,6853
patient|6853,6860
's|6860,6862
improving|6863,6872
clinical|6873,6881
status|6882,6888
,|6888,6889
the|6890,6893
decision|6894,6902
was|6903,6906
made|6907,6911
to|6912,6914
<EOL>|6915,6916
pursue|6916,6922
no|6923,6925
further|6926,6933
collection|6934,6944
drainage|6945,6953
at|6954,6956
this|6957,6961
time|6962,6966
.|6966,6967
<EOL>|6968,6969
4.|6969,6971
Severe|6973,6979
bilateral|6980,6989
hydronephrosis|6990,7004
,|7004,7005
as|7006,7008
on|7009,7011
prior|7012,7017
examinations|7018,7030
.|7030,7031
<EOL>|7032,7033
RECOMMENDATION|7033,7047
:|7047,7048
Given|7050,7055
persistence|7056,7067
of|7068,7070
severe|7071,7077
hydronephrosis|7078,7092
,|7092,7093
<EOL>|7094,7095
percutaneous|7095,7107
<EOL>|7108,7109
nephrostomy|7109,7120
tubes|7121,7126
should|7127,7133
be|7134,7136
considered|7137,7147
.|7147,7148
<EOL>|7149,7150
<EOL>|7150,7151
<EOL>|7152,7153
BRIEF|7176,7181
SUMMARY|7182,7189
:|7189,7190
<EOL>|7190,7191
=|7191,7192
=|7192,7193
=|7193,7194
=|7194,7195
=|7195,7196
=|7196,7197
=|7197,7198
=|7198,7199
=|7199,7200
=|7200,7201
=|7201,7202
=|7202,7203
=|7203,7204
=|7204,7205
<EOL>|7205,7206
_|7206,7207
_|7207,7208
_|7208,7209
year|7210,7214
old|7215,7218
women|7219,7224
with|7225,7229
a|7230,7231
history|7232,7239
of|7240,7242
bladder|7243,7250
cancer|7251,7257
s|7258,7259
/|7259,7260
p|7260,7261
<EOL>|7262,7263
cystectomy|7263,7273
,|7273,7274
hysterectomy|7275,7287
,|7287,7288
and|7289,7292
BSO|7293,7296
now|7297,7300
with|7301,7305
ileal|7306,7311
conduit|7312,7319
,|7319,7320
whose|7321,7326
<EOL>|7327,7328
post|7328,7332
operative|7333,7342
course|7343,7349
has|7350,7353
been|7354,7358
complicated|7359,7370
by|7371,7373
DVT|7374,7377
/|7377,7378
PE|7378,7380
,|7380,7381
ileus|7382,7387
,|7387,7388
and|7389,7392
<EOL>|7393,7394
pelvic|7394,7400
fluid|7401,7406
collections|7407,7418
w|7419,7420
/|7420,7421
one|7422,7425
LLQ|7426,7429
drain|7430,7435
presented|7436,7445
with|7446,7450
<EOL>|7451,7452
subjective|7452,7462
fevers|7463,7469
,|7469,7470
lethargy|7471,7479
,|7479,7480
and|7481,7484
bloody|7485,7491
drain|7492,7497
output|7498,7504
.|7504,7505
She|7506,7509
was|7510,7513
<EOL>|7514,7515
found|7515,7520
to|7521,7523
have|7524,7528
worsening|7529,7538
anemia|7539,7545
and|7546,7549
was|7550,7553
given|7554,7559
2|7560,7561
units|7562,7567
of|7568,7570
pRBC|7571,7575
<EOL>|7576,7577
with|7577,7581
appropriate|7582,7593
increase|7594,7602
in|7603,7605
hemoglobin|7606,7616
noted|7617,7622
.|7622,7623
She|7624,7627
was|7628,7631
also|7632,7636
<EOL>|7637,7638
found|7638,7643
on|7644,7646
CT|7647,7649
imaging|7650,7657
to|7658,7660
have|7661,7665
an|7666,7668
interval|7669,7677
increase|7678,7686
in|7687,7689
size|7690,7694
of|7695,7697
a|7698,7699
<EOL>|7700,7701
left|7701,7705
abdominal|7706,7715
fluid|7716,7721
collection|7722,7732
.|7732,7733
Decision|7734,7742
was|7743,7746
made|7747,7751
to|7752,7754
place|7755,7760
a|7761,7762
<EOL>|7763,7764
drain|7764,7769
per|7770,7773
ID|7774,7776
.|7776,7777
Fluid|7778,7783
was|7784,7787
sent|7788,7792
and|7793,7796
revealed|7797,7805
:|7805,7806
negative|7807,7815
cultures|7816,7824
,|7824,7825
<EOL>|7826,7827
negative|7827,7835
malignant|7836,7845
cells|7846,7851
,|7851,7852
no|7853,7855
evidence|7856,7864
of|7865,7867
lymphatic|7868,7877
or|7878,7880
urinary|7881,7888
<EOL>|7889,7890
fluid|7890,7895
.|7895,7896
This|7897,7901
new|7902,7905
drain|7906,7911
was|7912,7915
subsequently|7916,7928
removed|7929,7936
per|7937,7940
_|7941,7942
_|7942,7943
_|7943,7944
as|7945,7947
fluid|7948,7953
<EOL>|7954,7955
collection|7955,7965
was|7966,7969
completely|7970,7980
drained|7981,7988
.|7988,7989
The|7990,7993
prior|7994,7999
drain|8000,8005
was|8006,8009
still|8010,8015
<EOL>|8016,8017
draining|8017,8025
serosanguinous|8026,8040
fluid|8041,8046
and|8047,8050
was|8051,8054
kept|8055,8059
in|8060,8062
but|8063,8066
repositioned|8067,8079
.|8079,8080
<EOL>|8081,8082
ID|8082,8084
was|8085,8088
consulted|8089,8098
for|8099,8102
the|8103,8106
fevers|8107,8113
,|8113,8114
leukocytosis|8115,8127
and|8128,8131
fluid|8132,8137
<EOL>|8138,8139
collections|8139,8150
and|8151,8154
was|8155,8158
deemed|8159,8165
to|8166,8168
need|8169,8173
antibiotics|8174,8185
and|8186,8189
tranisitioned|8190,8203
<EOL>|8204,8205
from|8205,8209
broad|8210,8215
spectrum|8216,8224
to|8225,8227
IV|8228,8230
ertapenem|8231,8240
at|8241,8243
discharge|8244,8253
.|8253,8254
Will|8255,8259
require|8260,8267
<EOL>|8268,8269
multiple|8269,8277
follow|8278,8284
ups|8285,8288
and|8289,8292
imaging|8293,8300
as|8301,8303
specified|8304,8313
in|8314,8316
the|8317,8320
transitional|8321,8333
<EOL>|8334,8335
issues|8335,8341
.|8341,8342
<EOL>|8343,8344
<EOL>|8345,8346
ACUTE|8346,8351
ISSUES|8352,8358
:|8358,8359
<EOL>|8359,8360
=|8360,8361
=|8361,8362
=|8362,8363
=|8363,8364
=|8364,8365
=|8365,8366
=|8366,8367
=|8367,8368
=|8368,8369
=|8369,8370
=|8370,8371
=|8371,8372
=|8372,8373
<EOL>|8373,8374
#|8374,8375
Pelvic|8375,8381
fluid|8382,8387
collections|8388,8399
:|8399,8400
patient|8401,8408
arrived|8409,8416
with|8417,8421
one|8422,8425
anterior|8426,8434
<EOL>|8435,8436
drain|8436,8441
putting|8442,8449
out|8450,8453
serosanguinous|8454,8468
fluid|8469,8474
.|8474,8475
CT|8476,8478
abdomen|8479,8486
/|8486,8487
pelvis|8487,8493
<EOL>|8494,8495
revealed|8495,8503
enlarging|8504,8513
left|8514,8518
fluid|8519,8524
collection|8525,8535
,|8535,8536
and|8537,8540
decision|8541,8549
was|8550,8553
made|8554,8558
<EOL>|8559,8560
to|8560,8562
place|8563,8568
a|8569,8570
drain|8571,8576
per|8577,8580
_|8581,8582
_|8582,8583
_|8583,8584
.|8584,8585
The|8586,8589
fluid|8590,8595
was|8596,8599
negative|8600,8608
for|8609,8612
malignant|8613,8622
<EOL>|8623,8624
cells|8624,8629
.|8629,8630
The|8631,8634
fluid|8635,8640
had|8641,8644
Cr|8645,8647
1|8648,8649
and|8650,8653
triglycerides|8654,8667
<|8668,8669
9|8669,8670
suggesting|8671,8681
that|8682,8686
<EOL>|8687,8688
fluid|8688,8693
collection|8694,8704
is|8705,8707
neither|8708,8715
urine|8716,8721
nor|8722,8725
lymphatic|8726,8735
fluid|8736,8741
.|8741,8742
Fluid|8743,8748
<EOL>|8749,8750
culture|8750,8757
was|8758,8761
negative|8762,8770
for|8771,8774
bacteria|8775,8783
.|8783,8784
On|8785,8787
interval|8788,8796
imaging|8797,8804
,|8804,8805
the|8806,8809
new|8810,8813
<EOL>|8814,8815
enlarging|8815,8824
fluid|8825,8830
collection|8831,8841
had|8842,8845
completely|8846,8856
collapsed|8857,8866
and|8867,8870
the|8871,8874
<EOL>|8875,8876
drain|8876,8881
was|8882,8885
removed|8886,8893
.|8893,8894
As|8895,8897
for|8898,8901
the|8902,8905
other|8906,8911
fluid|8912,8917
collection|8918,8928
that|8929,8933
<EOL>|8934,8935
already|8935,8942
had|8943,8946
a|8947,8948
drain|8949,8954
putting|8955,8962
out|8963,8966
serosanguinous|8967,8981
fluid|8982,8987
,|8987,8988
it|8989,8991
<EOL>|8992,8993
continued|8993,9002
to|9003,9005
drain|9006,9011
serosanguinous|9012,9026
fluid|9027,9032
but|9033,9036
at|9037,9039
a|9040,9041
lower|9042,9047
rate|9048,9052
than|9053,9057
<EOL>|9058,9059
prior|9059,9064
to|9065,9067
admission|9068,9077
.|9077,9078
The|9079,9082
drain|9083,9088
was|9089,9092
left|9093,9097
in|9098,9100
place|9101,9106
as|9107,9109
the|9110,9113
fluid|9114,9119
<EOL>|9120,9121
collection|9121,9131
on|9132,9134
imaging|9135,9142
had|9143,9146
not|9147,9150
completely|9151,9161
collapsed|9162,9171
.|9171,9172
BID|9173,9176
-|9177,9178
N|9179,9180
<EOL>|9181,9182
cultures|9182,9190
for|9191,9194
the|9195,9198
aforementioned|9199,9213
fluid|9214,9219
collection|9220,9230
came|9231,9235
back|9236,9240
<EOL>|9241,9242
positive|9242,9250
for|9251,9254
MSSA|9255,9259
but|9260,9263
per|9264,9267
ID|9268,9270
,|9270,9271
does|9272,9276
not|9277,9280
reflect|9281,9288
rue|9289,9292
<EOL>|9293,9294
intra-abdominal|9294,9309
infection|9310,9319
.|9319,9320
Given|9321,9326
that|9327,9331
patient|9332,9339
had|9340,9343
a|9344,9345
fever|9346,9351
at|9352,9354
OSH|9355,9358
<EOL>|9359,9360
and|9360,9363
a|9364,9365
leukocytosis|9366,9378
,|9378,9379
she|9380,9383
was|9384,9387
placed|9388,9394
on|9395,9397
broad|9398,9403
spectrum|9404,9412
antibiotics|9413,9424
<EOL>|9425,9426
with|9426,9430
vanc|9431,9435
,|9435,9436
ceftaz|9437,9443
and|9444,9447
flagyl|9448,9454
.|9454,9455
This|9456,9460
was|9461,9464
tapered|9465,9472
per|9473,9476
ID|9477,9479
team|9480,9484
to|9485,9487
IV|9488,9490
<EOL>|9491,9492
zosyn|9492,9497
.|9497,9498
On|9499,9501
discharge|9502,9511
,|9511,9512
ID|9513,9515
recommended|9516,9527
ertapenem|9528,9537
for|9538,9541
approximately|9542,9555
<EOL>|9556,9557
4|9557,9558
weeks|9559,9564
with|9565,9569
final|9570,9575
length|9576,9582
of|9583,9585
treatment|9586,9595
to|9596,9598
be|9599,9601
determined|9602,9612
by|9613,9615
fluid|9616,9621
<EOL>|9622,9623
collection|9623,9633
changes|9634,9641
on|9642,9644
repeat|9645,9651
imaging|9652,9659
on|9660,9662
outpatient|9663,9673
basis|9674,9679
.|9679,9680
Mrs|9681,9684
.|9684,9685
<EOL>|9686,9687
_|9687,9688
_|9688,9689
_|9689,9690
remained|9691,9699
afebrile|9700,9708
,|9708,9709
and|9710,9713
leukocytosis|9714,9726
resolved|9727,9735
.|9735,9736
<EOL>|9737,9738
<EOL>|9738,9739
#|9739,9740
Pulmonary|9740,9749
embolism|9750,9758
:|9758,9759
Likely|9760,9766
developed|9767,9776
in|9777,9779
the|9780,9783
setting|9784,9791
of|9792,9794
being|9795,9800
<EOL>|9801,9802
diagnosed|9802,9811
with|9812,9816
a|9817,9818
post-op|9819,9826
DVT|9827,9830
.|9830,9831
She|9832,9835
was|9836,9839
placed|9840,9846
on|9847,9849
lovenox|9850,9857
.|9857,9858
She|9860,9863
<EOL>|9864,9865
was|9865,9868
transitioned|9869,9881
to|9882,9884
heparin|9885,9892
ggt|9893,9896
as|9897,9899
she|9900,9903
needed|9904,9910
_|9911,9912
_|9912,9913
_|9913,9914
procedures|9915,9925
and|9926,9929
<EOL>|9930,9931
was|9931,9934
transitioned|9935,9947
back|9948,9952
to|9953,9955
lovenox|9956,9963
but|9964,9967
at|9968,9970
a|9971,9972
lower|9973,9978
dose|9979,9983
per|9984,9987
weight|9988,9994
<EOL>|9995,9996
dosing|9996,10002
to|10003,10005
70mg|10006,10010
q12H|10011,10015
upon|10016,10020
discharge|10021,10030
.|10030,10031
<EOL>|10032,10033
<EOL>|10033,10034
#|10034,10035
Acute|10035,10040
renal|10041,10046
injury|10047,10053
:|10053,10054
SCr|10055,10058
has|10059,10062
been|10063,10067
steadily|10068,10076
rising|10077,10083
from|10084,10088
a|10089,10090
<EOL>|10091,10092
baseline|10092,10100
of|10101,10103
around|10104,10110
0.04|10111,10115
-|10115,10116
0.06|10116,10120
in|10121,10123
_|10124,10125
_|10125,10126
_|10126,10127
to|10128,10130
1.1|10131,10134
,|10134,10135
likely|10136,10142
<EOL>|10143,10144
_|10144,10145
_|10145,10146
_|10146,10147
obstructed|10148,10158
uropathy|10159,10167
_|10168,10169
_|10169,10170
_|10170,10171
large|10172,10177
pelbic|10178,10184
fluid|10185,10190
collections|10191,10202
.|10202,10203
_|10204,10205
_|10205,10206
_|10206,10207
<EOL>|10208,10209
resolved|10209,10217
over|10218,10222
the|10223,10226
course|10227,10233
of|10234,10236
her|10237,10240
hospital|10241,10249
stay|10250,10254
with|10255,10259
final|10260,10265
Cr|10266,10268
0.8|10269,10272
.|10272,10273
<EOL>|10274,10275
<EOL>|10275,10276
<EOL>|10276,10277
#|10277,10278
Hydronephrosis|10278,10292
:|10292,10293
bilateral|10294,10303
and|10304,10307
worsening|10308,10317
on|10318,10320
interval|10321,10329
imaging|10330,10337
<EOL>|10338,10339
from|10339,10343
prior|10344,10349
studies|10350,10357
.|10357,10358
Given|10359,10364
patient|10365,10372
's|10372,10374
age|10375,10378
,|10378,10379
adequate|10380,10388
urinary|10389,10396
<EOL>|10397,10398
output|10398,10404
,|10404,10405
adequate|10406,10414
creatinine|10415,10425
clearance|10426,10435
,|10435,10436
and|10437,10440
no|10441,10443
significant|10444,10455
<EOL>|10456,10457
electrolyte|10457,10468
abnormalities|10469,10482
,|10482,10483
patient|10484,10491
likely|10492,10498
would|10499,10504
not|10505,10508
<EOL>|10509,10510
significantly|10510,10523
benefit|10524,10531
from|10532,10536
intervention|10537,10549
at|10550,10552
this|10553,10557
time|10558,10562
.|10562,10563
Per|10564,10567
<EOL>|10568,10569
urology|10569,10576
consult|10577,10584
,|10584,10585
deemed|10586,10592
stable|10593,10599
for|10600,10603
discharge|10604,10613
and|10614,10617
recommended|10618,10629
<EOL>|10630,10631
outpatient|10631,10641
urology|10642,10649
followup|10650,10658
.|10658,10659
<EOL>|10660,10661
<EOL>|10661,10662
#|10662,10663
Anemia|10663,10669
:|10669,10670
likely|10671,10677
a|10678,10679
combination|10680,10691
of|10692,10694
anemia|10695,10701
of|10702,10704
chronic|10705,10712
inflammation|10713,10725
<EOL>|10726,10727
and|10727,10730
acute|10731,10736
blood|10737,10742
loss|10743,10747
_|10748,10749
_|10749,10750
_|10750,10751
to|10752,10754
anterior|10755,10763
abdominal|10764,10773
drain|10774,10779
showing|10780,10787
<EOL>|10788,10789
serosanguinous|10789,10803
fluid|10804,10809
.|10809,10810
Labs|10811,10815
not|10816,10819
consistent|10820,10830
with|10831,10835
hemolysis|10836,10845
.|10845,10846
<EOL>|10847,10848
Received|10848,10856
2|10857,10858
units|10859,10864
of|10865,10867
pRBC|10868,10872
with|10873,10877
appropriate|10878,10889
response|10890,10898
.|10898,10899
Patient|10900,10907
was|10908,10911
<EOL>|10912,10913
discharged|10913,10923
with|10924,10928
Hgb|10929,10932
of|10933,10935
8.3|10936,10939
per|10940,10943
hem|10944,10947
/|10947,10948
onc|10948,10951
recommendation|10952,10966
for|10967,10970
<EOL>|10971,10972
threshold|10972,10981
Hgb|10982,10985
>|10985,10986
8|10986,10987
as|10988,10990
patient|10991,10998
feels|10999,11004
and|11005,11008
functionally|11009,11021
performs|11022,11030
<EOL>|11031,11032
better|11032,11038
with|11039,11043
higher|11044,11050
blood|11051,11056
counts|11057,11063
.|11063,11064
<EOL>|11065,11066
<EOL>|11066,11067
#|11067,11068
Hypokalemia|11068,11079
:|11079,11080
was|11081,11084
hypokalemic|11085,11096
and|11097,11100
was|11101,11104
repleted|11105,11113
with|11114,11118
oral|11119,11123
KCl|11124,11127
<EOL>|11128,11129
PRN|11129,11132
.|11132,11133
<EOL>|11134,11135
<EOL>|11135,11136
CHRONIC|11136,11143
ISSUES|11144,11150
:|11150,11151
<EOL>|11151,11152
=|11152,11153
=|11153,11154
=|11154,11155
=|11155,11156
=|11156,11157
=|11157,11158
=|11158,11159
=|11159,11160
=|11160,11161
=|11161,11162
=|11162,11163
=|11163,11164
=|11164,11165
=|11165,11166
=|11166,11167
<EOL>|11167,11168
#|11168,11169
Invasive|11169,11177
high|11178,11182
-|11182,11183
grade|11183,11188
urothelial|11189,11199
carcinoma|11200,11209
,|11209,11210
involving|11211,11220
the|11221,11224
deep|11225,11229
<EOL>|11230,11231
muscularis|11231,11241
propria|11242,11249
<EOL>|11249,11250
S|11250,11251
/|11251,11252
p|11252,11253
cystectomy|11254,11264
,|11264,11265
hysterectomy|11266,11278
,|11278,11279
and|11280,11283
BSO|11284,11287
now|11288,11291
with|11292,11296
ileal|11297,11302
conduit|11303,11310
,|11310,11311
<EOL>|11312,11313
whose|11313,11318
post|11319,11323
operative|11324,11333
course|11334,11340
has|11341,11344
been|11345,11349
complicated|11350,11361
by|11362,11364
DVT|11365,11368
/|11368,11369
PE|11369,11371
,|11371,11372
<EOL>|11373,11374
ileus|11374,11379
,|11379,11380
and|11381,11384
pelvic|11385,11391
fluid|11392,11397
collections|11398,11409
.|11409,11410
Patient|11412,11419
stating|11420,11427
that|11428,11432
there|11433,11438
<EOL>|11439,11440
is|11440,11442
no|11443,11445
plan|11446,11450
for|11451,11454
chemo|11455,11460
and|11461,11464
radiation|11465,11474
,|11474,11475
her|11476,11479
PET|11480,11483
scan|11484,11488
does|11489,11493
show|11494,11498
<EOL>|11499,11500
concerning|11500,11510
foci|11511,11515
of|11516,11518
metastatic|11519,11529
disease|11530,11537
in|11538,11540
the|11541,11544
lung|11545,11549
and|11550,11553
<EOL>|11554,11555
peritoneum|11555,11565
.|11565,11566
Per|11567,11570
patient|11571,11578
's|11578,11580
son|11581,11584
,|11584,11585
Mrs.|11586,11590
_|11591,11592
_|11592,11593
_|11593,11594
has|11595,11598
seen|11599,11603
a|11604,11605
doctor|11606,11612
<EOL>|11613,11614
to|11614,11616
work|11617,11621
up|11622,11624
the|11625,11628
lung|11629,11633
mass|11634,11638
.|11638,11639
Will|11640,11644
need|11645,11649
ongoing|11650,11657
discussion|11658,11668
with|11669,11673
<EOL>|11674,11675
outpatient|11675,11685
hem|11686,11689
/|11689,11690
onc|11690,11693
regarding|11694,11703
how|11704,11707
to|11708,11710
best|11711,11715
manage|11716,11722
concerning|11723,11733
<EOL>|11734,11735
lesions|11735,11742
.|11742,11743
<EOL>|11744,11745
<EOL>|11745,11746
#|11746,11747
Breast|11747,11753
mass|11754,11758
_|11759,11760
_|11760,11761
_|11761,11762
mammogram|11763,11772
showing|11773,11780
BI-RADS|11781,11788
5|11789,11790
,|11790,11791
Solid|11792,11797
mass|11798,11802
<EOL>|11803,11804
in|11804,11806
the|11807,11810
3|11811,11812
o|11813,11814
'|11814,11815
clock|11815,11820
left|11821,11825
breast|11826,11832
with|11833,11837
features|11838,11846
of|11847,11849
a|11850,11851
highly|11852,11858
<EOL>|11859,11860
suspicious|11860,11870
for|11871,11874
malignancy|11875,11885
.|11885,11886
Per|11887,11890
patient|11891,11898
's|11898,11900
son|11901,11904
,|11904,11905
she|11906,11909
has|11910,11913
seen|11914,11918
a|11919,11920
<EOL>|11921,11922
doctor|11922,11928
for|11929,11932
evaluating|11933,11943
the|11944,11947
new|11948,11951
breast|11952,11958
mass|11959,11963
.|11963,11964
Would|11965,11970
recommend|11971,11980
<EOL>|11981,11982
ongoing|11982,11989
discussion|11990,12000
with|12001,12005
aforementioned|12006,12020
doctor|12021,12027
and|12028,12031
outpatient|12032,12042
<EOL>|12043,12044
hem|12044,12047
/|12047,12048
onc|12048,12051
about|12052,12057
plan|12058,12062
to|12063,12065
manage|12066,12072
.|12072,12073
<EOL>|12073,12074
<EOL>|12074,12075
#|12075,12076
HLD|12077,12080
:|12080,12081
continued|12082,12091
atorvastatin|12092,12104
without|12105,12112
changes|12113,12120
.|12120,12121
Consider|12122,12130
<EOL>|12131,12132
evaluation|12132,12142
regarding|12143,12152
stopping|12153,12161
atorvastatin|12162,12174
on|12175,12177
outpatient|12178,12188
basis|12189,12194
<EOL>|12195,12196
<EOL>|12197,12198
#|12198,12199
Hypothyroidism|12200,12214
:|12214,12215
continued|12216,12225
levothyroxine|12226,12239
without|12240,12247
changes|12248,12255
.|12255,12256
<EOL>|12259,12260
<EOL>|12262,12263
#|12263,12264
HCP|12264,12267
:|12267,12268
Dr.|12270,12273
_|12274,12275
_|12275,12276
_|12276,12277
(|12278,12279
son|12279,12282
,|12282,12283
_|12284,12285
_|12285,12286
_|12286,12287
physician|12288,12297
)|12297,12298
_|12299,12300
_|12300,12301
_|12301,12302
<EOL>|12302,12303
#|12303,12304
Code|12304,12308
status|12309,12315
:|12315,12316
full|12317,12321
code|12322,12326
(|12327,12328
confirmed|12328,12337
with|12338,12342
patient|12343,12350
on|12351,12353
_|12354,12355
_|12355,12356
_|12356,12357
<EOL>|12358,12359
<EOL>|12359,12360
TRANSITIONAL|12360,12372
ISSUES|12373,12379
:|12379,12380
<EOL>|12380,12381
=|12381,12382
=|12382,12383
=|12383,12384
=|12384,12385
=|12385,12386
=|12386,12387
=|12387,12388
=|12388,12389
=|12389,12390
=|12390,12391
=|12391,12392
=|12392,12393
=|12393,12394
=|12394,12395
=|12395,12396
=|12396,12397
=|12397,12398
=|12398,12399
=|12399,12400
=|12400,12401
<EOL>|12401,12402
[|12402,12403
]|12404,12405
Will|12406,12410
need|12411,12415
infectious|12416,12426
disease|12427,12434
follow|12435,12441
up|12442,12444
.|12444,12445
If|12446,12448
ID|12449,12451
has|12452,12455
not|12456,12459
<EOL>|12460,12461
contacted|12461,12470
Mrs|12471,12474
_|12475,12476
_|12476,12477
_|12477,12478
by|12479,12481
_|12482,12483
_|12483,12484
_|12484,12485
,|12485,12486
she|12487,12490
should|12491,12497
call|12498,12502
_|12503,12504
_|12504,12505
_|12505,12506
<EOL>|12507,12508
to|12508,12510
set|12511,12514
up|12515,12517
an|12518,12520
appointment|12521,12532
.|12532,12533
The|12534,12537
ID|12538,12540
appointment|12541,12552
needs|12553,12558
to|12559,12561
be|12562,12564
AFTER|12565,12570
<EOL>|12571,12572
her|12572,12575
CT|12576,12578
abdomen|12579,12586
/|12586,12587
pelvis|12587,12593
has|12594,12597
already|12598,12605
been|12606,12610
done|12611,12615
<EOL>|12616,12617
[|12617,12618
]|12619,12620
Assure|12621,12627
that|12628,12632
Mrs|12633,12636
_|12637,12638
_|12638,12639
_|12639,12640
has|12641,12644
her|12645,12648
CT|12649,12651
abdomen|12652,12659
&|12660,12661
pelvis|12662,12668
with|12669,12673
<EOL>|12674,12675
contrast|12675,12683
in|12684,12686
the|12687,12690
week|12691,12695
of|12696,12698
_|12699,12700
_|12700,12701
_|12701,12702
<EOL>|12702,12703
[|12703,12704
]|12705,12706
She|12707,12710
should|12711,12717
get|12718,12721
weekly|12722,12728
lab|12729,12732
draws|12733,12738
of|12739,12741
the|12742,12745
following|12746,12755
:|12755,12756
CBC|12757,12760
with|12761,12765
<EOL>|12766,12767
differential|12767,12779
,|12779,12780
BUN|12781,12784
,|12784,12785
Cr|12786,12788
,|12788,12789
AST|12790,12793
,|12793,12794
ALT|12795,12798
,|12798,12799
TB|12800,12802
,|12802,12803
ALK|12804,12807
PHOS|12808,12812
.|12812,12813
ALL|12814,12817
LAB|12818,12821
REQUESTS|12822,12830
<EOL>|12831,12832
SHOULD|12832,12838
BE|12839,12841
ANNOTATED|12842,12851
WITH|12852,12856
:|12856,12857
*|12858,12859
*|12859,12860
ATTN|12860,12864
:|12864,12865
_|12866,12867
_|12867,12868
_|12868,12869
CLINIC|12870,12876
-|12877,12878
FAX|12879,12882
:|12882,12883
<EOL>|12884,12885
_|12885,12886
_|12886,12887
_|12887,12888
<EOL>|12888,12889
[|12889,12890
]|12891,12892
If|12893,12895
possible|12896,12904
,|12904,12905
please|12906,12912
give|12913,12917
ertapenem|12918,12927
at|12928,12930
night|12931,12936
-|12936,12937
time|12937,12941
so|12942,12944
it|12945,12947
does|12948,12952
<EOL>|12953,12954
not|12954,12957
interfere|12958,12967
with|12968,12972
her|12973,12976
daily|12977,12982
activities|12983,12993
.|12993,12994
Tentatively|12995,13006
,|13006,13007
she|13008,13011
will|13012,13016
<EOL>|13017,13018
be|13018,13020
receiving|13021,13030
ertapenem|13031,13040
for|13041,13044
_|13045,13046
_|13046,13047
_|13047,13048
weeks|13049,13054
but|13055,13058
with|13059,13063
final|13064,13069
treatment|13070,13079
<EOL>|13080,13081
length|13081,13087
determined|13088,13098
by|13099,13101
the|13102,13105
infectious|13106,13116
disease|13117,13124
team|13125,13129
.|13129,13130
<EOL>|13131,13132
[|13132,13133
]|13134,13135
Will|13136,13140
need|13141,13145
ongoing|13146,13153
discussion|13154,13164
with|13165,13169
outpatient|13170,13180
PCP|13181,13184
and|13185,13188
hem|13189,13192
/|13192,13193
onc|13193,13196
<EOL>|13197,13198
regarding|13198,13207
how|13208,13211
to|13212,13214
manage|13215,13221
new|13222,13225
breast|13226,13232
lesion|13233,13239
and|13240,13243
lung|13244,13248
/|13248,13249
peritoneum|13249,13259
<EOL>|13260,13261
lesions|13261,13268
.|13268,13269
<EOL>|13270,13271
[|13271,13272
]|13273,13274
Reevaluate|13275,13285
need|13286,13290
for|13291,13294
atorvastatin|13295,13307
<EOL>|13307,13308
[|13308,13309
]|13310,13311
Will|13312,13316
need|13317,13321
outpatient|13322,13332
follow|13333,13339
up|13340,13342
with|13343,13347
urology|13348,13355
,|13355,13356
Dr.|13357,13360
_|13361,13362
_|13362,13363
_|13363,13364
<EOL>|13365,13366
his|13366,13369
team|13370,13374
regarding|13375,13384
worsening|13385,13394
hydronephrosis|13395,13409
<EOL>|13409,13410
<EOL>|13410,13411
<EOL>|13412,13413
Medications|13413,13424
on|13425,13427
Admission|13428,13437
:|13437,13438
<EOL>|13438,13439
The|13439,13442
Preadmission|13443,13455
Medication|13456,13466
list|13467,13471
is|13472,13474
accurate|13475,13483
and|13484,13487
complete|13488,13496
.|13496,13497
<EOL>|13497,13498
1.|13498,13500
Acetaminophen|13501,13514
650|13515,13518
mg|13519,13521
PO|13522,13524
Q6H|13525,13528
<EOL>|13529,13530
2.|13530,13532
Atorvastatin|13533,13545
10|13546,13548
mg|13549,13551
PO|13552,13554
QPM|13555,13558
<EOL>|13559,13560
3.|13560,13562
Enoxaparin|13563,13573
Sodium|13574,13580
90|13581,13583
mg|13584,13586
SC|13587,13589
Q12H|13590,13594
<EOL>|13595,13596
Start|13596,13601
:|13601,13602
_|13603,13604
_|13604,13605
_|13605,13606
,|13606,13607
First|13608,13613
Dose|13614,13618
:|13618,13619
Next|13620,13624
Routine|13625,13632
Administration|13633,13647
Time|13648,13652
<EOL>|13653,13654
4.|13654,13656
Levothyroxine|13657,13670
Sodium|13671,13677
175|13678,13681
mcg|13682,13685
PO|13686,13688
DAILY|13689,13694
<EOL>|13695,13696
5.|13696,13698
LORazepam|13699,13708
0.25|13709,13713
-|13713,13714
0|13714,13715
.|13715,13716
5|13716,13717
mg|13718,13720
PO|13721,13723
DAILY|13724,13729
:|13729,13730
PRN|13730,13733
anxiety|13734,13741
<EOL>|13742,13743
<EOL>|13743,13744
<EOL>|13745,13746
Discharge|13746,13755
Medications|13756,13767
:|13767,13768
<EOL>|13768,13769
1.|13769,13771
Ertapenem|13773,13782
Sodium|13783,13789
1|13790,13791
g|13792,13793
IV|13794,13796
1X|13797,13799
Duration|13800,13808
:|13808,13809
1|13810,13811
Dose|13812,13816
<EOL>|13817,13818
please|13818,13824
give|13825,13829
ertapenem|13830,13839
daily|13840,13845
,|13845,13846
preferably|13847,13857
at|13858,13860
nighttime|13861,13870
to|13871,13873
not|13874,13877
<EOL>|13878,13879
interfere|13879,13888
with|13889,13893
her|13894,13897
daily|13898,13903
activities|13904,13914
<EOL>|13916,13917
2.|13917,13919
Milk|13921,13925
of|13926,13928
Magnesia|13929,13937
30|13938,13940
mL|13941,13943
PO|13944,13946
Q6H|13947,13950
:|13950,13951
PRN|13951,13954
constipation|13955,13967
<EOL>|13969,13970
3.|13970,13972
Enoxaparin|13974,13984
Sodium|13985,13991
70|13992,13994
mg|13995,13997
SC|13998,14000
Q12H|14001,14005
<EOL>|14006,14007
Start|14007,14012
:|14012,14013
Today|14014,14019
-|14020,14021
_|14022,14023
_|14023,14024
_|14024,14025
,|14025,14026
First|14027,14032
Dose|14033,14037
:|14037,14038
Next|14039,14043
Routine|14044,14051
Administration|14052,14066
<EOL>|14067,14068
Time|14068,14072
<EOL>|14074,14075
4.|14075,14077
Acetaminophen|14079,14092
650|14093,14096
mg|14097,14099
PO|14100,14102
Q6H|14103,14106
<EOL>|14108,14109
5.|14109,14111
Atorvastatin|14113,14125
10|14126,14128
mg|14129,14131
PO|14132,14134
QPM|14135,14138
<EOL>|14140,14141
6.|14141,14143
Levothyroxine|14145,14158
Sodium|14159,14165
175|14166,14169
mcg|14170,14173
PO|14174,14176
DAILY|14177,14182
<EOL>|14184,14185
7.|14185,14187
LORazepam|14189,14198
0.25|14199,14203
-|14203,14204
0|14204,14205
.|14205,14206
5|14206,14207
mg|14208,14210
PO|14211,14213
DAILY|14214,14219
:|14219,14220
PRN|14220,14223
anxiety|14224,14231
<EOL>|14233,14234
<EOL>|14234,14235
<EOL>|14236,14237
Discharge|14237,14246
Disposition|14247,14258
:|14258,14259
<EOL>|14259,14260
Extended|14260,14268
Care|14269,14273
<EOL>|14273,14274
<EOL>|14275,14276
Facility|14276,14284
:|14284,14285
<EOL>|14285,14286
_|14286,14287
_|14287,14288
_|14288,14289
<EOL>|14289,14290
<EOL>|14291,14292
Discharge|14292,14301
Diagnosis|14302,14311
:|14311,14312
<EOL>|14312,14313
Primary|14313,14320
diagnosis|14321,14330
:|14330,14331
Pelvic|14332,14338
fluid|14339,14344
collection|14345,14355
infection|14356,14365
,|14365,14366
_|14367,14368
_|14368,14369
_|14369,14370
,|14370,14371
acute|14372,14377
<EOL>|14378,14379
blood|14379,14384
loss|14385,14389
anemia|14390,14396
<EOL>|14396,14397
<EOL>|14397,14398
Secondary|14398,14407
diagnosis|14408,14417
:|14417,14418
acute|14419,14424
renal|14425,14430
failure|14431,14438
,|14438,14439
acute|14440,14445
on|14446,14448
chronic|14449,14456
<EOL>|14457,14458
anemia|14458,14464
,|14464,14465
recent|14466,14472
pulmonary|14473,14482
embolism|14483,14491
,|14491,14492
invasive|14493,14501
high|14502,14506
-|14506,14507
grade|14507,14512
<EOL>|14513,14514
urothelial|14514,14524
carcinoma|14525,14534
,|14534,14535
left|14536,14540
breast|14541,14547
mass|14548,14552
(|14553,14554
BIRADS|14554,14560
5|14561,14562
)|14562,14563
,|14563,14564
<EOL>|14565,14566
hypothyroidism|14566,14580
<EOL>|14582,14583
<EOL>|14583,14584
<EOL>|14585,14586
Mental|14607,14613
Status|14614,14620
:|14620,14621
Clear|14622,14627
and|14628,14631
coherent|14632,14640
.|14640,14641
<EOL>|14641,14642
Level|14642,14647
of|14648,14650
Consciousness|14651,14664
:|14664,14665
Alert|14666,14671
and|14672,14675
interactive|14676,14687
.|14687,14688
<EOL>|14688,14689
Activity|14689,14697
Status|14698,14704
:|14704,14705
Ambulatory|14706,14716
-|14717,14718
requires|14719,14727
assistance|14728,14738
or|14739,14741
aid|14742,14745
(|14746,14747
walker|14747,14753
<EOL>|14754,14755
or|14755,14757
cane|14758,14762
)|14762,14763
.|14763,14764
<EOL>|14764,14765
<EOL>|14765,14766
<EOL>|14767,14768
Dear|14792,14796
_|14797,14798
_|14798,14799
_|14799,14800
,|14800,14801
<EOL>|14801,14802
<EOL>|14802,14803
_|14803,14804
_|14804,14805
_|14805,14806
did|14807,14810
you|14811,14814
come|14815,14819
to|14820,14822
the|14823,14826
hospital|14827,14835
?|14835,14836
<EOL>|14836,14837
-|14837,14838
You|14839,14842
were|14843,14847
feeling|14848,14855
tired|14856,14861
and|14862,14865
your|14866,14870
drain|14871,14876
output|14877,14883
was|14884,14887
bloody|14888,14894
.|14894,14895
<EOL>|14896,14897
<EOL>|14897,14898
What|14898,14902
happened|14903,14911
at|14912,14914
the|14915,14918
hospital|14919,14927
?|14927,14928
<EOL>|14928,14929
-|14929,14930
A|14931,14932
CT|14933,14935
scan|14936,14940
showed|14941,14947
very|14948,14952
large|14953,14958
fluid|14959,14964
collections|14965,14976
in|14977,14979
your|14980,14984
pelvis|14985,14991
<EOL>|14992,14993
-|14993,14994
The|14995,14998
radiologists|14999,15011
placed|15012,15018
another|15019,15026
drain|15027,15032
and|15033,15036
removed|15037,15044
it|15045,15047
once|15048,15052
it|15053,15055
<EOL>|15056,15057
appeared|15057,15065
that|15066,15070
the|15071,15074
large|15075,15080
fluid|15081,15086
collection|15087,15097
was|15098,15101
gone|15102,15106
<EOL>|15106,15107
-|15107,15108
You|15109,15112
were|15113,15117
given|15118,15123
a|15124,15125
blood|15126,15131
transfusion|15132,15143
<EOL>|15143,15144
-|15144,15145
We|15146,15148
placed|15149,15155
a|15156,15157
PICC|15158,15162
(|15163,15164
a|15164,15165
long|15166,15170
IV|15171,15173
)|15173,15174
so|15175,15177
that|15178,15182
you|15183,15186
can|15187,15190
receive|15191,15198
<EOL>|15199,15200
antibiotics|15200,15211
after|15212,15217
you|15218,15221
get|15222,15225
discharged|15226,15236
from|15237,15241
the|15242,15245
hospital|15246,15254
<EOL>|15254,15255
<EOL>|15255,15256
What|15256,15260
needs|15261,15266
to|15267,15269
happen|15270,15276
when|15277,15281
you|15282,15285
leave|15286,15291
the|15292,15295
hospital|15296,15304
?|15304,15305
<EOL>|15305,15306
-|15306,15307
Please|15308,15314
continue|15315,15323
seeing|15324,15330
the|15331,15334
doctors|15335,15342
that|15343,15347
are|15348,15351
_|15352,15353
_|15353,15354
_|15354,15355
your|15356,15360
<EOL>|15361,15362
lung|15362,15366
and|15367,15370
breast|15371,15377
lesions|15378,15385
and|15386,15389
follow|15390,15396
their|15397,15402
recommendations|15403,15418
.|15418,15419
<EOL>|15420,15421
-|15421,15422
Continue|15423,15431
taking|15432,15438
Lovenox|15439,15446
every|15447,15452
day|15453,15456
to|15457,15459
treat|15460,15465
the|15466,15469
blood|15470,15475
clot|15476,15480
in|15481,15483
<EOL>|15484,15485
your|15485,15489
lung|15490,15494
.|15494,15495
<EOL>|15496,15497
-|15497,15498
If|15499,15501
the|15502,15505
infectious|15506,15516
disease|15517,15524
doctor|15525,15531
has|15532,15535
not|15536,15539
contacted|15540,15549
you|15550,15553
by|15554,15556
_|15557,15558
_|15558,15559
_|15559,15560
,|15560,15561
please|15562,15568
call|15569,15573
the|15574,15577
following|15578,15587
number|15588,15594
to|15595,15597
set|15598,15601
up|15602,15604
an|15605,15607
appointment|15608,15619
:|15619,15620
<EOL>|15621,15622
_|15622,15623
_|15623,15624
_|15624,15625
.|15625,15626
<EOL>|15627,15628
-|15628,15629
Please|15630,15636
make|15637,15641
sure|15642,15646
you|15647,15650
have|15651,15655
a|15656,15657
repeat|15658,15664
CT|15665,15667
scan|15668,15672
done|15673,15677
BEFORE|15678,15684
your|15685,15689
<EOL>|15690,15691
appointment|15691,15702
with|15703,15707
the|15708,15711
infectious|15712,15722
disease|15723,15730
doctor|15731,15737
<EOL>|15737,15738
-|15738,15739
You|15740,15743
will|15744,15748
be|15749,15751
getting|15752,15759
IV|15760,15762
antibiotics|15763,15774
for|15775,15778
several|15779,15786
weeks|15787,15792
.|15792,15793
The|15794,15797
<EOL>|15798,15799
infectious|15799,15809
disease|15810,15817
doctor|15818,15824
_|15825,15826
_|15826,15827
_|15827,15828
determine|15829,15838
how|15839,15842
long|15843,15847
you|15848,15851
will|15852,15856
need|15857,15861
<EOL>|15862,15863
to|15863,15865
be|15866,15868
on|15869,15871
it|15872,15874
.|15874,15875
<EOL>|15876,15877
<EOL>|15877,15878
It|15878,15880
was|15881,15884
a|15885,15886
pleasure|15887,15895
taking|15896,15902
care|15903,15907
of|15908,15910
you|15911,15914
.|15914,15915
<EOL>|15916,15917
Your|15917,15921
_|15922,15923
_|15923,15924
_|15924,15925
team|15926,15930
<EOL>|15931,15932
<EOL>|15933,15934
Followup|15934,15942
Instructions|15943,15955
:|15955,15956
<EOL>|15956,15957
_|15957,15958
_|15958,15959
_|15959,15960
<EOL>|15960,15961

