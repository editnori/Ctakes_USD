 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|34,38
No|39,41
:|41,42
_|45,46
_|46,47
_|47,48
<EOL>|48,49
<EOL>|50,51
Admission|51,60
Date|61,65
:|65,66
_|68,69
_|69,70
_|70,71
Discharge|85,94
Date|95,99
:|99,100
_|103,104
_|104,105
_|105,106
<EOL>|106,107
<EOL>|108,109
Date|109,113
of|114,116
Birth|117,122
:|122,123
_|125,126
_|126,127
_|127,128
Sex|141,144
:|144,145
M|148,149
<EOL>|149,150
<EOL>|151,152
Service|152,159
:|159,160
MEDICINE|161,169
<EOL>|169,170
<EOL>|171,172
Allergies|172,181
:|181,182
<EOL>|183,184
No|184,186
Known|187,192
Allergies|193,202
/|203,204
Adverse|205,212
Drug|213,217
Reactions|218,227
<EOL>|227,228
<EOL>|229,230
Attending|230,239
:|239,240
_|241,242
_|242,243
_|243,244
.|244,245
<EOL>|245,246
<EOL>|247,248
Chief|248,253
Complaint|254,263
:|263,264
<EOL>|264,265
Right|265,270
flank|271,276
bruising|277,285
and|286,289
pain|290,294
s|295,296
/|296,297
p|297,298
fall|299,303
<EOL>|303,304
<EOL>|305,306
Major|306,311
Surgical|312,320
or|321,323
Invasive|324,332
Procedure|333,342
:|342,343
<EOL>|343,344
None|344,348
<EOL>|348,349
<EOL>|349,350
<EOL>|351,352
History|352,359
of|360,362
Present|363,370
Illness|371,378
:|378,379
<EOL>|379,380
Mr.|380,383
_|384,385
_|385,386
_|386,387
is|388,390
a|391,392
_|393,394
_|394,395
_|395,396
with|397,401
history|402,409
of|410,412
factor|413,419
VIII|420,424
deficiency|425,435
who|436,439
<EOL>|440,441
presents|441,449
with|450,454
right|455,460
neck|461,465
swelling|466,474
after|475,480
snowboarding|481,493
accident|494,502
.|502,503
<EOL>|504,505
The|505,508
patient|509,516
reports|517,524
that|525,529
he|530,532
fell|533,537
while|538,543
snowboarding|544,556
with|557,561
loss|562,566
of|567,569
<EOL>|570,571
consciousness|571,584
on|585,587
_|588,589
_|589,590
_|590,591
.|591,592
He|593,595
was|596,599
initially|600,609
seen|610,614
at|615,617
<EOL>|618,619
_|619,620
_|620,621
_|621,622
where|623,628
CT|629,631
imaging|632,639
of|640,642
head|643,647
/|647,648
neck|648,652
showed|653,659
no|660,662
<EOL>|663,664
intracranial|664,676
hemorrhage|677,687
.|687,688
A|689,690
CTA|691,694
neck|695,699
showed|700,706
a|707,708
thickened|709,718
right|719,724
<EOL>|725,726
platysma|726,734
muscle|735,741
with|742,746
surrounding|747,758
hematoma|759,767
and|768,771
a|772,773
focus|774,779
of|780,782
active|783,789
<EOL>|790,791
contrast|791,799
extravasation|800,813
within|814,820
the|821,824
right|825,830
platysma|831,839
muscle|840,846
.|846,847
He|848,850
also|851,855
<EOL>|856,857
developed|857,866
a|867,868
right|869,874
shoulder|875,883
hematoma|884,892
although|893,901
shoulder|902,910
plain|911,916
<EOL>|917,918
films|918,923
did|924,927
n't|927,930
show|931,935
acute|936,941
abnormality|942,953
.|953,954
He|955,957
was|958,961
seen|962,966
by|967,969
_|970,971
_|971,972
_|972,973
<EOL>|974,975
Hematology|975,985
and|986,989
gave|990,994
him|995,998
one|999,1002
dose|1003,1007
of|1008,1010
DDAVP|1011,1016
IV|1017,1019
.|1019,1020
A|1021,1022
factor|1023,1029
VIII|1030,1034
<EOL>|1035,1036
assay|1036,1041
was|1042,1045
139|1046,1049
and|1050,1053
vW|1054,1056
level|1057,1062
was|1063,1066
>|1067,1068
200|1068,1071
per|1072,1075
report|1076,1082
.|1082,1083
Per|1084,1087
report|1088,1094
,|1094,1095
his|1096,1099
<EOL>|1100,1101
hemoglobin|1101,1111
decreased|1112,1121
from|1122,1126
13.2|1127,1131
on|1132,1134
_|1135,1136
_|1136,1137
_|1137,1138
to|1139,1141
11.6|1142,1146
on|1147,1149
_|1150,1151
_|1151,1152
_|1152,1153
.|1153,1154
<EOL>|1155,1156
Repeat|1156,1162
imaging|1163,1170
in|1171,1173
the|1174,1177
morning|1178,1185
showed|1186,1192
stable|1193,1199
injuries|1200,1208
.|1208,1209
The|1210,1213
<EOL>|1214,1215
patient|1215,1222
saw|1223,1226
his|1227,1230
hematologist|1231,1243
on|1244,1246
_|1247,1248
_|1248,1249
_|1249,1250
and|1251,1254
was|1255,1258
found|1259,1264
to|1265,1267
have|1268,1272
a|1273,1274
<EOL>|1275,1276
hemoglobin|1276,1286
of|1287,1289
10.4|1290,1294
.|1294,1295
Because|1296,1303
of|1304,1306
the|1307,1310
continued|1311,1320
mild|1321,1325
decrease|1326,1334
,|1334,1335
the|1336,1339
<EOL>|1340,1341
patient|1341,1348
followed|1349,1357
up|1358,1360
with|1361,1365
his|1366,1369
PCP|1370,1373
_|1374,1375
_|1375,1376
_|1376,1377
_|1378,1379
_|1379,1380
_|1380,1381
at|1382,1384
which|1385,1390
time|1391,1395
his|1396,1399
<EOL>|1400,1401
hemoglobin|1401,1411
was|1412,1415
9.9|1416,1419
.|1419,1420
He|1421,1423
was|1424,1427
found|1428,1433
to|1434,1436
have|1437,1441
an|1442,1444
enlarging|1445,1454
flank|1455,1460
<EOL>|1461,1462
hematoma|1462,1470
,|1470,1471
thus|1472,1476
was|1477,1480
referred|1481,1489
given|1490,1495
concern|1496,1503
for|1504,1507
retroperitoneal|1508,1523
<EOL>|1524,1525
bleed|1525,1530
.|1530,1531
The|1532,1535
patient|1536,1543
has|1544,1547
been|1548,1552
using|1553,1558
DDAVP|1559,1564
intranasally|1565,1577
<EOL>|1578,1579
intermittently|1579,1593
since|1594,1599
the|1600,1603
accident|1604,1612
.|1612,1613
He|1614,1616
denies|1617,1623
lightheadedness|1624,1639
or|1640,1642
<EOL>|1643,1644
palpitations|1644,1656
,|1656,1657
any|1658,1661
increase|1662,1670
in|1671,1673
neck|1674,1678
swelling|1679,1687
over|1688,1692
the|1693,1696
course|1697,1703
of|1704,1706
<EOL>|1707,1708
the|1708,1711
week|1712,1716
.|1716,1717
He|1718,1720
does|1721,1725
endorse|1726,1733
pain|1734,1738
in|1739,1741
his|1742,1745
right|1746,1751
shoulder|1752,1760
_|1761,1762
_|1762,1763
_|1763,1764
<EOL>|1765,1766
resting|1766,1773
,|1773,1774
_|1775,1776
_|1776,1777
_|1777,1778
moving|1779,1785
)|1785,1786
,|1786,1787
though|1788,1794
this|1795,1799
has|1800,1803
improved|1804,1812
over|1813,1817
the|1818,1821
course|1822,1828
<EOL>|1829,1830
of|1830,1832
the|1833,1836
week|1837,1841
.|1841,1842
<EOL>|1844,1845
In|1845,1847
the|1848,1851
ED|1852,1854
,|1854,1855
initial|1856,1863
vital|1864,1869
signs|1870,1875
were|1876,1880
99.2|1881,1885
87|1886,1888
124|1889,1892
/|1892,1893
75|1893,1895
18|1896,1898
100|1899,1902
%|1902,1903
/|1903,1904
RA|1904,1906
.|1906,1907
<EOL>|1908,1909
Initial|1909,1916
labs|1917,1921
demonstrated|1922,1934
hemoglobin|1935,1945
10.6|1946,1950
,|1950,1951
though|1952,1958
repeat|1959,1965
was|1966,1969
<EOL>|1970,1971
9.7|1971,1974
.|1974,1975
Chemistries|1976,1987
and|1988,1991
coags|1992,1997
were|1998,2002
unremarkable|2003,2015
.|2015,2016
FVIII|2017,2022
activity|2023,2031
was|2032,2035
<EOL>|2036,2037
103|2037,2040
.|2040,2041
A|2042,2043
CTAP|2044,2048
was|2049,2052
performed|2053,2062
which|2063,2068
demonstrated|2069,2081
muscular|2082,2090
hemorrhage|2091,2101
<EOL>|2102,2103
along|2103,2108
the|2109,2112
flank|2113,2118
,|2118,2119
but|2120,2123
no|2124,2126
retroperitoneal|2127,2142
bleed|2143,2148
on|2149,2151
preliminary|2152,2163
<EOL>|2164,2165
read|2165,2169
.|2169,2170
The|2171,2174
patient|2175,2182
's|2182,2184
outpatient|2185,2195
hematologist|2196,2208
,|2208,2209
Dr.|2210,2213
_|2214,2215
_|2215,2216
_|2216,2217
,|2217,2218
was|2219,2222
<EOL>|2223,2224
contacted|2224,2233
and|2234,2237
it|2238,2240
was|2241,2244
decided|2245,2252
to|2253,2255
give|2256,2260
the|2261,2264
patient|2265,2272
desmopressin|2273,2285
<EOL>|2286,2287
0.3|2287,2290
mg|2290,2292
/|2292,2293
kg|2293,2295
IV|2296,2298
.|2298,2299
The|2300,2303
patient|2304,2311
was|2312,2315
then|2316,2320
admitted|2321,2329
for|2330,2333
futher|2334,2340
<EOL>|2341,2342
management|2342,2352
.|2352,2353
<EOL>|2355,2356
Per|2356,2359
review|2360,2366
of|2367,2369
records|2370,2377
,|2377,2378
the|2379,2382
patient|2383,2390
has|2391,2394
a|2395,2396
history|2397,2404
of|2405,2407
significant|2408,2419
<EOL>|2420,2421
bleeding|2421,2429
after|2430,2435
his|2436,2439
circumcision|2440,2452
,|2452,2453
requiring|2454,2463
blood|2464,2469
transfusion|2470,2481
.|2481,2482
<EOL>|2483,2484
Throughout|2484,2494
childhood|2495,2504
,|2504,2505
he|2506,2508
also|2509,2513
had|2514,2517
a|2518,2519
tendency|2520,2528
to|2529,2531
bruise|2532,2538
easily|2539,2545
.|2545,2546
<EOL>|2547,2548
He|2548,2550
was|2551,2554
tested|2555,2561
and|2562,2565
found|2566,2571
to|2572,2574
have|2575,2579
_|2580,2581
_|2581,2582
_|2582,2583
disease|2584,2591
.|2591,2592
Later|2593,2598
,|2598,2599
<EOL>|2600,2601
after|2601,2606
wisdom|2607,2613
tooth|2614,2619
extraction|2620,2630
,|2630,2631
the|2632,2635
patient|2636,2643
experienced|2644,2655
late|2656,2660
<EOL>|2661,2662
(|2662,2663
e|2663,2664
.|2664,2665
g|2665,2666
.|2666,2667
_|2668,2669
_|2669,2670
_|2670,2671
days|2672,2676
later|2677,2682
)|2682,2683
bleeding|2684,2692
despite|2693,2700
treatment|2701,2710
with|2711,2715
DDAVP|2716,2721
.|2721,2722
The|2723,2726
<EOL>|2727,2728
patient|2728,2735
was|2736,2739
retested|2740,2748
by|2749,2751
a|2752,2753
hematologist|2754,2766
associated|2767,2777
with|2778,2782
the|2783,2786
<EOL>|2787,2788
_|2788,2789
_|2789,2790
_|2790,2791
and|2792,2795
was|2796,2799
diagnosed|2800,2809
<EOL>|2810,2811
with|2811,2815
hemophilia|2816,2826
A.|2827,2829
His|2830,2833
FVIII|2834,2839
activity|2840,2848
has|2849,2852
been|2853,2857
checked|2858,2865
on|2866,2868
<EOL>|2869,2870
multiple|2870,2878
occasions|2879,2888
,|2888,2889
sometimes|2890,2899
testing|2900,2907
normal|2908,2914
,|2914,2915
though|2916,2922
has|2923,2926
been|2927,2931
as|2932,2934
<EOL>|2935,2936
low|2936,2939
as|2940,2942
~|2943,2944
50|2944,2946
.|2946,2947
<EOL>|2949,2950
Upon|2950,2954
arrival|2955,2962
to|2963,2965
the|2966,2969
floor|2970,2975
,|2975,2976
the|2977,2980
patient|2981,2988
is|2989,2991
comfortable|2992,3003
without|3004,3011
<EOL>|3012,3013
complaint|3013,3022
.|3022,3023
<EOL>|3025,3026
Review|3026,3032
of|3033,3035
Systems|3036,3043
:|3043,3044
<EOL>|3046,3047
(|3047,3048
+|3048,3049
)|3049,3050
per|3051,3054
HPI|3055,3058
<EOL>|3060,3061
(|3061,3062
-|3062,3063
)|3063,3064
fever|3065,3070
,|3070,3071
chills|3072,3078
,|3078,3079
night|3080,3085
sweats|3086,3092
,|3092,3093
headache|3094,3102
,|3102,3103
vision|3104,3110
changes|3111,3118
,|3118,3119
<EOL>|3120,3121
rhinorrhea|3121,3131
,|3131,3132
congestion|3133,3143
,|3143,3144
sore|3145,3149
throat|3150,3156
,|3156,3157
cough|3158,3163
,|3163,3164
shortness|3165,3174
of|3175,3177
breath|3178,3184
,|3184,3185
<EOL>|3186,3187
chest|3187,3192
pain|3193,3197
,|3197,3198
abdominal|3199,3208
pain|3209,3213
,|3213,3214
nausea|3215,3221
,|3221,3222
vomiting|3223,3231
,|3231,3232
diarrhea|3233,3241
,|3241,3242
<EOL>|3243,3244
constipation|3244,3256
,|3256,3257
BRBPR|3258,3263
,|3263,3264
melena|3265,3271
,|3271,3272
hematochezia|3273,3285
,|3285,3286
dysuria|3287,3294
,|3294,3295
hematuria|3296,3305
.|3305,3306
<EOL>|3306,3307
<EOL>|3308,3309
Past|3309,3313
Medical|3314,3321
History|3322,3329
:|3329,3330
<EOL>|3330,3331
-|3331,3332
Factor|3332,3338
VIII|3339,3343
deficiency|3344,3354
(|3355,3356
mild|3356,3360
)|3360,3361
<EOL>|3363,3364
<EOL>|3364,3365
<EOL>|3366,3367
Social|3367,3373
History|3374,3381
:|3381,3382
<EOL>|3382,3383
_|3383,3384
_|3384,3385
_|3385,3386
<EOL>|3386,3387
Family|3387,3393
History|3394,3401
:|3401,3402
<EOL>|3402,3403
The|3403,3406
patient|3407,3414
's|3414,3416
mother|3417,3423
had|3424,3427
tendency|3428,3436
to|3437,3439
bleed|3440,3445
.|3445,3446
<EOL>|3448,3449
<EOL>|3449,3450
<EOL>|3451,3452
Physical|3452,3460
Exam|3461,3465
:|3465,3466
<EOL>|3466,3467
ON|3467,3469
ADMISSION|3470,3479
<EOL>|3479,3480
VS|3480,3482
:|3482,3483
98|3483,3485
120|3486,3489
/|3489,3490
40|3490,3492
64|3493,3495
20|3496,3498
100RA|3499,3504
<EOL>|3506,3507
GENERAL|3507,3514
:|3514,3515
lying|3516,3521
flat|3522,3526
in|3527,3529
bed|3530,3533
,|3533,3534
no|3535,3537
acute|3538,3543
distress|3544,3552
<EOL>|3554,3555
HEENT|3555,3560
:|3560,3561
NCAT|3562,3566
,|3566,3567
MMM|3568,3571
,|3571,3572
OP|3573,3575
clear|3576,3581
<EOL>|3583,3584
NECK|3584,3588
:|3588,3589
Supple|3590,3596
<EOL>|3598,3599
CARDIAC|3599,3606
:|3606,3607
RRR|3608,3611
,|3611,3612
S1|3613,3615
/|3615,3616
S2|3616,3618
,|3618,3619
no|3620,3622
murmurs|3623,3630
,|3630,3631
gallops|3632,3639
,|3639,3640
or|3641,3643
rubs|3644,3648
<EOL>|3650,3651
LUNG|3651,3655
:|3655,3656
Generally|3657,3666
CTA|3667,3670
b|3671,3672
/|3672,3673
l|3673,3674
<EOL>|3676,3677
ABDOMEN|3677,3684
:|3684,3685
Soft|3686,3690
,|3690,3691
non-tender|3692,3702
,|3702,3703
non-distended|3704,3717
<EOL>|3719,3720
EXTREMITIES|3720,3731
:|3731,3732
Warm|3733,3737
,|3737,3738
well|3739,3743
-|3743,3744
perfused|3744,3752
<EOL>|3754,3755
PULSES|3755,3761
:|3761,3762
2|3763,3764
+|3764,3765
DP|3766,3768
pulses|3769,3775
bilaterally|3776,3787
<EOL>|3789,3790
NEURO|3790,3795
:|3795,3796
CN|3797,3799
II|3800,3802
-|3802,3803
XII|3803,3806
intact|3807,3813
<EOL>|3815,3816
SKIN|3816,3820
:|3820,3821
Hematomas|3822,3831
on|3832,3834
right|3835,3840
aspect|3841,3847
of|3848,3850
neck|3851,3855
and|3856,3859
flank|3860,3865
<EOL>|3866,3867
<EOL>|3867,3868
ON|3868,3870
DISCHARGE|3871,3880
<EOL>|3880,3881
Vitals|3881,3887
:|3887,3888
98.0|3889,3893
,|3893,3894
100|3895,3898
-|3898,3899
120|3899,3902
/|3902,3903
40|3903,3905
-|3905,3906
58|3906,3908
,|3908,3909
66|3910,3912
,|3912,3913
20|3914,3916
,|3916,3917
99|3918,3920
on|3921,3923
RA|3924,3926
<EOL>|3928,3929
GENERAL|3929,3936
:|3936,3937
lying|3938,3943
flat|3944,3948
in|3949,3951
bed|3952,3955
,|3955,3956
no|3957,3959
acute|3960,3965
distress|3966,3974
<EOL>|3976,3977
HEENT|3977,3982
:|3982,3983
NCAT|3984,3988
,|3988,3989
MMM|3990,3993
,|3993,3994
OP|3995,3997
clear|3998,4003
<EOL>|4005,4006
NECK|4006,4010
:|4010,4011
Supple|4012,4018
<EOL>|4020,4021
CARDIAC|4021,4028
:|4028,4029
RRR|4030,4033
,|4033,4034
S1|4035,4037
/|4037,4038
S2|4038,4040
,|4040,4041
no|4042,4044
murmurs|4045,4052
,|4052,4053
gallops|4054,4061
,|4061,4062
or|4063,4065
rubs|4066,4070
<EOL>|4072,4073
LUNG|4073,4077
:|4077,4078
Generally|4079,4088
CTA|4089,4092
b|4093,4094
/|4094,4095
l|4095,4096
<EOL>|4098,4099
ABDOMEN|4099,4106
:|4106,4107
Soft|4108,4112
,|4112,4113
non-tender|4114,4124
,|4124,4125
non-distended|4126,4139
<EOL>|4141,4142
EXTREMITIES|4142,4153
:|4153,4154
Warm|4155,4159
,|4159,4160
well|4161,4165
-|4165,4166
perfused|4166,4174
<EOL>|4176,4177
PULSES|4177,4183
:|4183,4184
2|4185,4186
+|4186,4187
DP|4188,4190
pulses|4191,4197
bilaterally|4198,4209
<EOL>|4211,4212
NEURO|4212,4217
:|4217,4218
CN|4219,4221
II|4222,4224
-|4224,4225
XII|4225,4228
intact|4229,4235
<EOL>|4237,4238
SKIN|4238,4242
:|4242,4243
Hematomas|4244,4253
on|4254,4256
right|4257,4262
aspect|4263,4269
of|4270,4272
neck|4273,4277
and|4278,4281
flank|4282,4287
<EOL>|4287,4288
<EOL>|4288,4289
<EOL>|4290,4291
Pertinent|4291,4300
Results|4301,4308
:|4308,4309
<EOL>|4309,4310
ADMISSION|4310,4319
,|4319,4320
DISCHARGE|4321,4330
,|4330,4331
PERTINENT|4332,4341
LABS|4342,4346
:|4346,4347
<EOL>|4347,4348
<EOL>|4348,4349
_|4349,4350
_|4350,4351
_|4351,4352
07|4353,4355
:|4355,4356
03PM|4356,4360
BLOOD|4361,4366
WBC|4367,4370
-|4370,4371
6.6|4371,4374
RBC|4375,4378
-|4378,4379
3|4379,4380
.|4380,4381
58|4381,4383
*|4383,4384
Hgb|4385,4388
-|4388,4389
10|4389,4391
.|4391,4392
6|4392,4393
*|4393,4394
#|4394,4395
Hct|4396,4399
-|4399,4400
29|4400,4402
.|4402,4403
8|4403,4404
*|4404,4405
#|4405,4406
<EOL>|4407,4408
MCV|4408,4411
-|4411,4412
83|4412,4414
MCH|4415,4418
-|4418,4419
29.6|4419,4423
MCHC|4424,4428
-|4428,4429
35|4429,4431
.|4431,4432
6|4432,4433
*|4433,4434
RDW|4435,4438
-|4438,4439
14.7|4439,4443
Plt|4444,4447
_|4448,4449
_|4449,4450
_|4450,4451
<EOL>|4451,4452
_|4452,4453
_|4453,4454
_|4454,4455
07|4456,4458
:|4458,4459
03PM|4459,4463
BLOOD|4464,4469
Neuts|4470,4475
-|4475,4476
69.7|4476,4480
_|4481,4482
_|4482,4483
_|4483,4484
Monos|4485,4490
-|4490,4491
7.2|4491,4494
Eos|4495,4498
-|4498,4499
2.4|4499,4502
<EOL>|4503,4504
Baso|4504,4508
-|4508,4509
0.2|4509,4512
<EOL>|4512,4513
_|4513,4514
_|4514,4515
_|4515,4516
07|4517,4519
:|4519,4520
03PM|4520,4524
BLOOD|4525,4530
_|4531,4532
_|4532,4533
_|4533,4534
PTT|4535,4538
-|4538,4539
35.2|4539,4543
_|4544,4545
_|4545,4546
_|4546,4547
<EOL>|4547,4548
_|4548,4549
_|4549,4550
_|4550,4551
07|4552,4554
:|4554,4555
03PM|4555,4559
BLOOD|4560,4565
Plt|4566,4569
_|4570,4571
_|4571,4572
_|4572,4573
<EOL>|4573,4574
_|4574,4575
_|4575,4576
_|4576,4577
07|4578,4580
:|4580,4581
03PM|4581,4585
BLOOD|4586,4591
FacVIII|4592,4599
-|4599,4600
103|4600,4603
<EOL>|4603,4604
_|4604,4605
_|4605,4606
_|4606,4607
07|4608,4610
:|4610,4611
03PM|4611,4615
BLOOD|4616,4621
Glucose|4622,4629
-|4629,4630
93|4630,4632
UreaN|4633,4638
-|4638,4639
15|4639,4641
Creat|4642,4647
-|4647,4648
0.8|4648,4651
Na|4652,4654
-|4654,4655
139|4655,4658
<EOL>|4659,4660
K|4660,4661
-|4661,4662
4.1|4662,4665
Cl|4666,4668
-|4668,4669
101|4669,4672
HCO3|4673,4677
-|4677,4678
28|4678,4680
AnGap|4681,4686
-|4686,4687
14|4687,4689
<EOL>|4689,4690
_|4690,4691
_|4691,4692
_|4692,4693
11|4694,4696
:|4696,4697
00PM|4697,4701
BLOOD|4702,4707
WBC|4708,4711
-|4711,4712
6.6|4712,4715
RBC|4716,4719
-|4719,4720
3|4720,4721
.|4721,4722
30|4722,4724
*|4724,4725
Hgb|4726,4729
-|4729,4730
9|4730,4731
.|4731,4732
7|4732,4733
*|4733,4734
Hct|4735,4738
-|4738,4739
27|4739,4741
.|4741,4742
0|4742,4743
*|4743,4744
<EOL>|4745,4746
MCV|4746,4749
-|4749,4750
82|4750,4752
MCH|4753,4756
-|4756,4757
29.4|4757,4761
MCHC|4762,4766
-|4766,4767
36|4767,4769
.|4769,4770
0|4770,4771
*|4771,4772
RDW|4773,4776
-|4776,4777
14.7|4777,4781
Plt|4782,4785
_|4786,4787
_|4787,4788
_|4788,4789
<EOL>|4789,4790
_|4790,4791
_|4791,4792
_|4792,4793
07|4794,4796
:|4796,4797
25AM|4797,4801
BLOOD|4802,4807
WBC|4808,4811
-|4811,4812
5.2|4812,4815
RBC|4816,4819
-|4819,4820
3|4820,4821
.|4821,4822
14|4822,4824
*|4824,4825
Hgb|4826,4829
-|4829,4830
9|4830,4831
.|4831,4832
3|4832,4833
*|4833,4834
Hct|4835,4838
-|4838,4839
26|4839,4841
.|4841,4842
2|4842,4843
*|4843,4844
<EOL>|4845,4846
MCV|4846,4849
-|4849,4850
83|4850,4852
MCH|4853,4856
-|4856,4857
29.7|4857,4861
MCHC|4862,4866
-|4866,4867
35|4867,4869
.|4869,4870
7|4870,4871
*|4871,4872
RDW|4873,4876
-|4876,4877
14.6|4877,4881
Plt|4882,4885
_|4886,4887
_|4887,4888
_|4888,4889
<EOL>|4889,4890
_|4890,4891
_|4891,4892
_|4892,4893
03|4894,4896
:|4896,4897
25PM|4897,4901
BLOOD|4902,4907
WBC|4908,4911
-|4911,4912
6.3|4912,4915
RBC|4916,4919
-|4919,4920
3|4920,4921
.|4921,4922
27|4922,4924
*|4924,4925
Hgb|4926,4929
-|4929,4930
9|4930,4931
.|4931,4932
9|4932,4933
*|4933,4934
Hct|4935,4938
-|4938,4939
27|4939,4941
.|4941,4942
1|4942,4943
*|4943,4944
<EOL>|4945,4946
MCV|4946,4949
-|4949,4950
83|4950,4952
MCH|4953,4956
-|4956,4957
30.3|4957,4961
MCHC|4962,4966
-|4966,4967
36|4967,4969
.|4969,4970
5|4970,4971
*|4971,4972
RDW|4973,4976
-|4976,4977
14.7|4977,4981
Plt|4982,4985
_|4986,4987
_|4987,4988
_|4988,4989
<EOL>|4989,4990
_|4990,4991
_|4991,4992
_|4992,4993
07|4994,4996
:|4996,4997
50PM|4997,5001
URINE|5002,5007
Color|5008,5013
-|5013,5014
Yellow|5014,5020
Appear|5021,5027
-|5027,5028
Clear|5028,5033
Sp|5034,5036
_|5037,5038
_|5038,5039
_|5039,5040
<EOL>|5040,5041
_|5041,5042
_|5042,5043
_|5043,5044
07|5045,5047
:|5047,5048
50PM|5048,5052
URINE|5053,5058
Blood|5059,5064
-|5064,5065
NEG|5065,5068
Nitrite|5069,5076
-|5076,5077
NEG|5077,5080
Protein|5081,5088
-|5088,5089
30|5089,5091
<EOL>|5092,5093
Glucose|5093,5100
-|5100,5101
NEG|5101,5104
Ketone|5105,5111
-|5111,5112
NEG|5112,5115
Bilirub|5116,5123
-|5123,5124
NEG|5124,5127
Urobiln|5128,5135
-|5135,5136
NEG|5136,5139
pH|5140,5142
-|5142,5143
6.0|5143,5146
Leuks|5147,5152
-|5152,5153
NEG|5153,5156
<EOL>|5156,5157
_|5157,5158
_|5158,5159
_|5159,5160
07|5161,5163
:|5163,5164
50PM|5164,5168
URINE|5169,5174
RBC|5175,5178
-|5178,5179
<|5179,5180
1|5180,5181
WBC|5182,5185
-|5185,5186
1|5186,5187
Bacteri|5188,5195
-|5195,5196
FEW|5196,5199
Yeast|5200,5205
-|5205,5206
NONE|5206,5210
Epi|5211,5214
-|5214,5215
0|5215,5216
<EOL>|5216,5217
_|5217,5218
_|5218,5219
_|5219,5220
07|5221,5223
:|5223,5224
50PM|5224,5228
URINE|5229,5234
Mucous|5235,5241
-|5241,5242
RARE|5242,5246
<EOL>|5246,5247
<EOL>|5247,5248
IMAGING|5248,5255
/|5255,5256
STUDIES|5256,5263
:|5263,5264
<EOL>|5264,5265
<EOL>|5266,5267
_|5267,5268
_|5268,5269
_|5269,5270
CT|5271,5273
A|5274,5275
/|5275,5276
P|5276,5277
<EOL>|5277,5278
Acute|5278,5283
hemorrhage|5284,5294
along|5295,5300
right|5301,5306
posterior|5307,5316
flank|5317,5322
musculature|5323,5334
and|5335,5338
<EOL>|5339,5340
probably|5340,5348
layering|5349,5357
over|5358,5362
it|5363,5365
,|5365,5366
only|5367,5371
partly|5372,5378
imaged|5379,5385
and|5386,5389
hard|5390,5394
to|5395,5397
<EOL>|5398,5399
distinguish|5399,5410
musculature|5411,5422
from|5423,5427
hemorrhage|5428,5438
.|5438,5439
No|5440,5442
active|5443,5449
extravasation|5450,5463
<EOL>|5464,5465
seen|5465,5469
.|5469,5470
Probable|5471,5479
old|5480,5483
hematoma|5484,5492
along|5493,5498
posterior|5499,5508
left|5509,5513
flank|5514,5519
.|5519,5520
<EOL>|5521,5522
<EOL>|5522,5523
<EOL>|5524,5525
Brief|5525,5530
Hospital|5531,5539
Course|5540,5546
:|5546,5547
<EOL>|5547,5548
Mr.|5548,5551
_|5552,5553
_|5553,5554
_|5554,5555
is|5556,5558
a|5559,5560
_|5561,5562
_|5562,5563
_|5563,5564
with|5565,5569
history|5570,5577
of|5578,5580
mild|5581,5585
FVIII|5586,5591
deficiency|5592,5602
who|5603,5606
<EOL>|5607,5608
presents|5608,5616
after|5617,5622
snowboarding|5623,5635
accident|5636,5644
with|5645,5649
multiple|5650,5658
hematomas|5659,5668
and|5669,5672
<EOL>|5673,5674
falling|5674,5681
hemoglobin|5682,5692
concerning|5693,5703
for|5704,5707
ongoing|5708,5715
bleeding|5716,5724
.|5724,5725
<EOL>|5725,5726
<EOL>|5726,5727
#|5727,5728
FACTOR|5729,5735
VIII|5736,5740
DEFICIENCY|5741,5751
,|5751,5752
MULTIPLE|5753,5761
HEMATOMAS|5762,5771
:|5771,5772
Patient|5773,5780
presented|5781,5790
<EOL>|5791,5792
after|5792,5797
recent|5798,5804
snowboarding|5805,5817
accident|5818,5826
.|5826,5827
At|5828,5830
_|5831,5832
_|5832,5833
_|5833,5834
<EOL>|5835,5836
_|5836,5837
_|5837,5838
_|5838,5839
,|5839,5840
imaging|5841,5848
was|5849,5852
notable|5853,5860
for|5861,5864
neck|5865,5869
and|5870,5873
shoulder|5874,5882
hematomas|5883,5892
.|5892,5893
<EOL>|5894,5895
Upon|5895,5899
reevaluation|5900,5912
by|5913,5915
his|5916,5919
PCP|5920,5923
,|5923,5924
the|5925,5928
patient|5929,5936
was|5937,5940
found|5941,5946
to|5947,5949
have|5950,5954
a|5955,5956
<EOL>|5957,5958
flank|5958,5963
hematoma|5964,5972
.|5972,5973
Given|5974,5979
falling|5980,5987
hemoglobin|5988,5998
,|5998,5999
there|6000,6005
was|6006,6009
concern|6010,6017
for|6018,6021
<EOL>|6022,6023
retroperitoneal|6023,6038
bleed|6039,6044
.|6044,6045
CTAP|6046,6050
in|6051,6053
the|6054,6057
ED|6058,6060
demonstrated|6061,6073
hematoma|6074,6082
over|6083,6087
<EOL>|6088,6089
his|6089,6092
flank|6093,6098
musculature|6099,6110
,|6110,6111
but|6112,6115
no|6116,6118
active|6119,6125
extravasation|6126,6139
.|6139,6140
He|6141,6143
was|6144,6147
given|6148,6153
<EOL>|6154,6155
IV|6155,6157
DDAVP|6158,6163
,|6163,6164
but|6165,6168
FVIII|6169,6174
activity|6175,6183
was|6184,6187
103|6188,6191
(|6192,6193
wnl|6193,6196
)|6196,6197
.|6197,6198
CBC|6199,6202
remained|6203,6211
stable|6212,6218
<EOL>|6219,6220
and|6220,6223
patient|6224,6231
declined|6232,6240
further|6241,6248
inpatient|6249,6258
monitoring|6259,6269
.|6269,6270
Atrius|6271,6277
<EOL>|6278,6279
hematology|6279,6289
recommended|6290,6301
continued|6302,6311
outpatient|6312,6322
hemoglobin|6323,6333
<EOL>|6334,6335
monitoring|6335,6345
,|6345,6346
but|6347,6350
did|6351,6354
not|6355,6358
think|6359,6364
further|6365,6372
DDAVP|6373,6378
was|6379,6382
indicated|6383,6392
given|6393,6398
<EOL>|6399,6400
normal|6400,6406
FVIII|6407,6412
level|6413,6418
.|6418,6419
<EOL>|6420,6421
<EOL>|6423,6424
<EOL>|6424,6425
#|6425,6426
TRANISTIONAL|6427,6439
ISSUES|6440,6446
:|6446,6447
<EOL>|6447,6448
-|6448,6449
PCP|6450,6453
_|6454,6455
_|6455,6456
_|6456,6457
_|6458,6459
_|6459,6460
_|6460,6461
<EOL>|6461,6462
-|6462,6463
CBC|6464,6467
_|6468,6469
_|6469,6470
_|6470,6471
-|6472,6473
_|6474,6475
_|6475,6476
_|6476,6477
at|6478,6480
_|6481,6482
_|6482,6483
_|6483,6484
<EOL>|6484,6485
-|6485,6486
Caution|6487,6494
to|6495,6497
avoid|6498,6503
dangerous|6504,6513
activity|6514,6522
<EOL>|6522,6523
-|6523,6524
Code|6525,6529
:|6529,6530
presumed|6531,6539
full|6540,6544
<EOL>|6546,6547
-|6547,6548
Emergency|6549,6558
Contact|6559,6566
:|6566,6567
_|6568,6569
_|6569,6570
_|6570,6571
_|6572,6573
_|6573,6574
_|6574,6575
-|6576,6577
wife|6578,6582
)|6582,6583
<EOL>|6584,6585
<EOL>|6586,6587
Medications|6587,6598
on|6599,6601
Admission|6602,6611
:|6611,6612
<EOL>|6612,6613
The|6613,6616
Preadmission|6617,6629
Medication|6630,6640
list|6641,6645
is|6646,6648
accurate|6649,6657
and|6658,6661
complete|6662,6670
.|6670,6671
<EOL>|6671,6672
1.|6672,6674
Desmopressin|6675,6687
Nasal|6688,6693
_|6694,6695
_|6695,6696
_|6696,6697
mcg|6698,6701
NAS|6702,6705
PRN|6706,6709
bleeding|6710,6718
<EOL>|6719,6720
<EOL>|6720,6721
<EOL>|6722,6723
Discharge|6723,6732
Medications|6733,6744
:|6744,6745
<EOL>|6745,6746
1.|6746,6748
Acetaminophen|6749,6762
1000|6763,6767
mg|6768,6770
PO|6771,6773
Q8H|6774,6777
pain|6778,6782
<EOL>|6783,6784
2.|6784,6786
Desmopressin|6787,6799
Nasal|6800,6805
_|6806,6807
_|6807,6808
_|6808,6809
mcg|6810,6813
NAS|6814,6817
PRN|6818,6821
bleeding|6822,6830
<EOL>|6831,6832
3.|6832,6834
Outpatient|6835,6845
Lab|6846,6849
Work|6850,6854
<EOL>|6854,6855
CBC|6855,6858
on|6859,6861
_|6862,6863
_|6863,6864
_|6864,6865
or|6866,6868
_|6869,6870
_|6870,6871
_|6871,6872
.|6872,6873
Last|6874,6878
hemoglobin|6879,6889
9.9|6890,6893
_|6894,6895
_|6895,6896
_|6896,6897
_|6898,6899
_|6899,6900
_|6900,6901
.|6901,6902
<EOL>|6902,6903
<EOL>|6903,6904
<EOL>|6905,6906
Discharge|6906,6915
Disposition|6916,6927
:|6927,6928
<EOL>|6928,6929
Home|6929,6933
<EOL>|6933,6934
<EOL>|6935,6936
Discharge|6936,6945
Diagnosis|6946,6955
:|6955,6956
<EOL>|6956,6957
PRIMARY|6957,6964
:|6964,6965
<EOL>|6965,6966
-|6966,6967
Acute|6968,6973
muscular|6974,6982
hematoma|6983,6991
,|6991,6992
right|6993,6998
flank|6999,7004
<EOL>|7004,7005
-|7005,7006
Hemophilia|7007,7017
,|7017,7018
factor|7019,7025
VIII|7026,7030
deficiency|7031,7041
<EOL>|7041,7042
<EOL>|7042,7043
<EOL>|7044,7045
Discharge|7045,7054
Condition|7055,7064
:|7064,7065
<EOL>|7065,7066
Mental|7066,7072
Status|7073,7079
:|7079,7080
Clear|7081,7086
and|7087,7090
coherent|7091,7099
.|7099,7100
<EOL>|7100,7101
Level|7101,7106
of|7107,7109
Consciousness|7110,7123
:|7123,7124
Alert|7125,7130
and|7131,7134
interactive|7135,7146
.|7146,7147
<EOL>|7147,7148
Activity|7148,7156
Status|7157,7163
:|7163,7164
Ambulatory|7165,7175
-|7176,7177
Independent|7178,7189
.|7189,7190
<EOL>|7190,7191
<EOL>|7191,7192
<EOL>|7193,7194
Discharge|7194,7203
Instructions|7204,7216
:|7216,7217
<EOL>|7217,7218
Mr.|7218,7221
_|7222,7223
_|7223,7224
_|7224,7225
,|7225,7226
<EOL>|7226,7227
<EOL>|7227,7228
It|7228,7230
was|7231,7234
our|7235,7238
pleasure|7239,7247
caring|7248,7254
for|7255,7258
you|7259,7262
at|7263,7265
_|7266,7267
_|7267,7268
_|7268,7269
<EOL>|7270,7271
_|7271,7272
_|7272,7273
_|7273,7274
.|7274,7275
You|7276,7279
were|7280,7284
admitted|7285,7293
with|7294,7298
bruising|7299,7307
on|7308,7310
your|7311,7315
right|7316,7321
<EOL>|7322,7323
side|7323,7327
and|7328,7331
low|7332,7335
blood|7336,7341
counts|7342,7348
after|7349,7354
a|7355,7356
snowboarding|7357,7369
fall|7370,7374
.|7374,7375
With|7376,7380
your|7381,7385
<EOL>|7386,7387
history|7387,7394
of|7395,7397
hemophilia|7398,7408
,|7408,7409
it|7410,7412
was|7413,7416
important|7417,7426
to|7427,7429
evaluate|7430,7438
internal|7439,7447
<EOL>|7448,7449
bleeding|7449,7457
which|7458,7463
did|7464,7467
show|7468,7472
a|7473,7474
right|7475,7480
muscular|7481,7489
flank|7490,7495
blood|7496,7501
collection|7502,7512
.|7512,7513
<EOL>|7514,7515
Your|7515,7519
facotr|7520,7526
VIII|7527,7531
level|7532,7537
was|7538,7541
103|7542,7545
and|7546,7549
you|7550,7553
received|7554,7562
IV|7563,7565
DDAVP|7566,7571
under|7572,7577
<EOL>|7578,7579
our|7579,7582
care|7583,7587
.|7587,7588
Your|7589,7593
blood|7594,7599
counts|7600,7606
were|7607,7611
stable|7612,7618
to|7619,7621
improved|7622,7630
on|7631,7633
the|7634,7637
day|7638,7641
<EOL>|7642,7643
of|7643,7645
admission|7646,7655
.|7655,7656
<EOL>|7657,7658
<EOL>|7658,7659
It|7659,7661
is|7662,7664
important|7665,7674
that|7675,7679
you|7680,7683
not|7684,7687
participate|7688,7699
in|7700,7702
any|7703,7706
dangerous|7707,7716
<EOL>|7717,7718
activities|7718,7728
given|7729,7734
your|7735,7739
recent|7740,7746
bleed|7747,7752
and|7753,7756
your|7757,7761
hemophilia|7762,7772
.|7772,7773
Bleeding|7774,7782
<EOL>|7783,7784
in|7784,7786
hemophiliacs|7787,7799
has|7800,7803
more|7804,7808
potential|7809,7818
to|7819,7821
be|7822,7824
life|7825,7829
-|7829,7830
threatening|7830,7841
.|7841,7842
<EOL>|7842,7843
<EOL>|7843,7844
Please|7844,7850
get|7851,7854
your|7855,7859
blood|7860,7865
counts|7866,7872
checked|7873,7880
at|7881,7883
_|7884,7885
_|7885,7886
_|7886,7887
site|7888,7892
on|7893,7895
either|7896,7902
<EOL>|7903,7904
_|7904,7905
_|7905,7906
_|7906,7907
or|7908,7910
_|7911,7912
_|7912,7913
_|7913,7914
.|7914,7915
Follow|7916,7922
up|7923,7925
with|7926,7930
your|7931,7935
<EOL>|7936,7937
regular|7937,7944
doctor|7945,7951
early|7952,7957
next|7958,7962
week|7963,7967
.|7967,7968
<EOL>|7968,7969
<EOL>|7969,7970
Best|7970,7974
wishes|7975,7981
,|7981,7982
<EOL>|7982,7983
Your|7983,7987
_|7988,7989
_|7989,7990
_|7990,7991
Care|7992,7996
Team|7997,8001
<EOL>|8001,8002
<EOL>|8003,8004
Followup|8004,8012
Instructions|8013,8025
:|8025,8026
<EOL>|8026,8027
_|8027,8028
_|8028,8029
_|8029,8030
<EOL>|8030,8031

