CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Neurology speciality|Title|false|false||NEUROLOGYnull|sulfa|Drug|false|false||Sulfanull|Sulfonamides, ophthalmologic antiinfectives|Drug|false|false||Sulfonamides
null|Sulfonamide Anti-Infective Agents|Drug|false|false||Sulfonamides
null|Sulfonamide Anti-Infective Agents|Drug|false|false||Sulfonamides
null|Sulfonamides, topical|Drug|false|false||Sulfonamides
null|Sulfonamides|Drug|false|false||Sulfonamides
null|Sulfonamides|Drug|false|false||Sulfonamides
null|Sulfonamides, ophthalmologic antiinfectives|Drug|false|false||Sulfonamides
null|Sulfonamides, Gynecological|Drug|false|false||Sulfonamides
null|Sulfonamides, Gynecological|Drug|false|false||Sulfonamides
null|Sulfonamides, intestinal antiinfectives|Drug|false|false||Sulfonamides
null|Sulfonamides, intestinal antiinfectives|Drug|false|false||Sulfonamidesnull|Poisoning by, adverse effect of and underdosing of sulfonamides|Disorder|false|false||Sulfonamides
null|Poisoning by sulfonamide|Disorder|false|false||Sulfonamidesnull|Adverse reaction to sulfonamides|Finding|false|false||Sulfonamidesnull|penicillins|Drug|false|false||Penicillins
null|penicillins|Drug|false|false||Penicillinsnull|Poisoning by, adverse effect of and underdosing of penicillins|Disorder|false|false||Penicillins
null|Poisoning by penicillin|Disorder|false|false||Penicillinsnull|Adverse reaction to penicillins|Finding|false|false||Penicillinsnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Facial Paresis|Disorder|false|false||Facial weaknessnull|Face|Anatomy|false|false||Facialnull|Facial|Modifier|false|false||Facialnull|Weakness|Finding|false|false||weakness
null|Asthenia|Finding|false|false||weaknessnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Proline dehydrogenase deficiency|Disorder|false|false||HPInull|History of present illness (finding)|Finding|false|false||HPI
null|allene oxide synthase activity|Finding|false|false||HPInull|Rhomboid fossa structure|Anatomy|false|false||RHFnull|Gastroesophageal reflux disease|Disorder|false|false||GERDnull|Mild depression|Disorder|false|false||mild depressionnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Cancer patients and suicide and depression|Disorder|false|false||depression
null|Mental Depression|Disorder|false|false||depression
null|Depressive disorder|Disorder|false|false||depression
null|Depressed mood|Disorder|false|false||depressionnull|Depression - motion|Finding|false|false||depression
null|null|Finding|false|false||depressionnull|Depression - recess|Modifier|false|false||depressionnull|null|Time|false|false||priornull|Migraine Disorders|Disorder|false|false||migrainesnull|Episode of|Time|false|false||episode ofnull|Episode of|Time|false|false||episodenull|Numbness of face|Finding|false|false||facial numbnessnull|Face|Anatomy|false|false||facialnull|Facial|Modifier|false|false||facialnull|Numbness|Finding|false|false||numbness
null|Hypesthesia|Finding|false|false||numbnessnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|FANCONI ANEMIA, COMPLEMENTATION GROUP E|Disorder|false|false||facenull|FANCE wt Allele|Finding|false|false||face
null|FANCE gene|Finding|false|false||face
null|ELOVL6 gene|Finding|false|false||facenull|Head>Face|Anatomy|false|false||face
null|Face|Anatomy|false|false||facenull|Face (spatial concept)|Modifier|false|false||facenull|Watching TV|Finding|false|false||watching TVnull|Watching|Finding|false|false||watchingnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|FANCONI ANEMIA, COMPLEMENTATION GROUP E|Disorder|false|false||facenull|FANCE wt Allele|Finding|false|false||face
null|FANCE gene|Finding|false|false||face
null|ELOVL6 gene|Finding|false|false||facenull|Head>Face|Anatomy|false|false||face
null|Face|Anatomy|false|false||facenull|Face (spatial concept)|Modifier|false|false||facenull|Numb (emotional response)|Finding|false|false||numb
null|NUMB gene|Finding|false|false||numbnull|Distribution [PK]|Finding|false|false||distribution
null|Distribution|Finding|false|false||distributionnull|Spatial Distribution|Modifier|false|false||distributionnull|Jaw|Anatomy|false|false||jawnull|Jaw Device|Device|false|false||jawnull|Line Specimen|Drug|false|false||line
null|Long Interspersed Elements|Drug|false|false||line
null|Long Interspersed Elements|Drug|false|false||linenull|line source specimen code|Finding|false|false||linenull|Intravascular line|Device|false|false||linenull|Linear|Modifier|false|false||linenull|Line Unit of Length|LabModifier|false|false||linenull|Initially|Time|false|false||initiallynull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Diffuse|Modifier|false|false||diffusenull|Dull pain|Finding|false|false||dullnull|Dull sensation quality|Modifier|false|false||dull
null|Dull|Modifier|false|false||dullnull|Unusual|Modifier|false|false||unusualnull|Migraine Disorders|Disorder|false|false||migrainenull|Usual|Modifier|false|false||typicalnull|Migraine Disorders|Disorder|false|false||migrainesnull|Numbness|Finding|false|false||numbness
null|Hypesthesia|Finding|false|false||numbnessnull|Minute of time|Time|false|false||minutesnull|Minute Unit of Plane Angle|LabModifier|false|false||minutes
null|Minute (diminutive)|LabModifier|false|false||minutes
null|Small|LabModifier|false|false||minutesnull|Completely - dosing instruction fragment|Finding|false|false||completelynull|Complete|Modifier|false|false||completelynull|Associated with|Modifier|false|false||associatednull|Weakness|Finding|false|false||weakness
null|Asthenia|Finding|false|false||weaknessnull|Sensory (qualifier value)|Modifier|false|false||sensorynull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|FANCONI ANEMIA, COMPLEMENTATION GROUP E|Disorder|false|false||facenull|FANCE wt Allele|Finding|false|false||face
null|FANCE gene|Finding|false|false||face
null|ELOVL6 gene|Finding|false|false||facenull|Head>Face|Anatomy|false|false||face
null|Face|Anatomy|false|false||facenull|Face (spatial concept)|Modifier|false|false||facenull|Vertigo as late effect of cerebrovascular disease|Disorder|false|false||vertigonull|Vertigo|Finding|false|false||vertigonull|Vertigo <Vertiginidae>|Entity|false|false||vertigonull|Language Disorders|Disorder|false|false||language impairmentnull|Programming Languages|Finding|false|false||languagenull|null|Attribute|false|false||languagenull|Languages|Entity|false|false||languagenull|Impaired health|Finding|false|false||impairment
null|Impaired|Finding|false|false||impairmentnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Extended Priority Codes - Routine|Finding|false|false||routine
null|Report priority - Routine|Finding|false|false||routine
null|Admission Type - Routine|Finding|false|false||routine
null|Level of Care - Routine|Finding|false|false||routine
null|Processing priority - Routine|Finding|false|false||routine
null|Referral priority - Routine|Finding|false|false||routinenull|Routine coag|Procedure|false|false||routinenull|Priority - Routine|Time|false|false||routinenull|Routine|Modifier|false|false||routinenull|Reactive Oxygen Species|Drug|false|false||ROS
null|rosiglitazone|Drug|false|false||ROS
null|rosiglitazone|Drug|false|false||ROS
null|Reactive Oxygen Species|Drug|false|false||ROSnull|ROS1 wt Allele|Finding|false|false||ROS
null|ROS1 gene|Finding|false|false||ROSnull|Review of systems (procedure)|Procedure|false|false||ROSnull|rostral sulcus|Anatomy|false|false||ROSnull|2 Weeks|Time|false|false||2 weeksnull|week|Time|false|false||weeksnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|rectal discharge diarrhea (physical finding)|Finding|false|false||diarrhea
null|Diarrhea|Finding|false|false||diarrheanull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Feelings|Finding|false|false||feelingnull|4 days ago|Time|false|false||4 days agonull|4 Days|Time|false|false||4 daysnull|day|Time|false|false||daysnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|Health|Finding|false|false||healthnull|Gastroesophageal reflux disease|Disorder|false|false||GERDnull|Mild depression|Disorder|false|false||mild depressionnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Cancer patients and suicide and depression|Disorder|false|false||depression
null|Mental Depression|Disorder|false|false||depression
null|Depressive disorder|Disorder|false|false||depression
null|Depressed mood|Disorder|false|false||depressionnull|Depression - motion|Finding|false|false||depression
null|null|Finding|false|false||depressionnull|Depression - recess|Modifier|false|false||depressionnull|Migraine Disorders|Disorder|false|false||migrainesnull|Mental association|Finding|false|false||assocnull|Associated with|Modifier|false|false||assocnull|Photopsia|Disorder|false|false||visual flashesnull|Visual|Finding|false|false||visualnull|Photopsia|Disorder|false|false||flashes of lightnull|Photopsia|Disorder|false|false||flashesnull|Light Sources, Flash|Device|false|false||flashesnull|Natural flashes|Phenomenon|false|false||flashesnull|TNFSF14 protein, human|Drug|false|false||light
null|TNFSF14 protein, human|Drug|false|false||lightnull|Light - subjective measurement|Finding|false|false||light
null|TNFSF14 wt Allele|Finding|false|false||light
null|TNFSF14 gene|Finding|false|false||light
null|Light color|Finding|false|false||lightnull|Phototherapy|Procedure|false|false||lightnull|Light|Phenomenon|false|false||lightnull|Light (qualifier)|Modifier|false|false||lightnull|Last|Modifier|false|false||lastnull|year|Time|false|false||yearsnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|Bunion|Disorder|false|false||bunionsnull|Indirect exposure mechanism - Father|Finding|false|false||Father
null|Relationship - Father|Finding|false|false||Father
null|Father - courtesy title|Finding|false|false||Fathernull|Father (person)|Subject|false|false||Fathernull|Cerebrovascular accident|Disorder|false|false||strokenull|Stroke (heart beat)|Finding|false|false||strokenull|Cardiac Catheterization Procedures|Procedure|false|false||cardiac cathnull|Cardiac attachment|Finding|false|false||cardiacnull|Heart|Anatomy|false|false||cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||cardiacnull|Catheterization|Procedure|false|false||cathnull|Late|Time|false|false||Laternull|Life|Finding|false|false||lifenull|Laser-Induced Fluorescence Endoscopy|Procedure|false|false||lifenull|Indirect exposure mechanism - Father|Finding|false|false||father
null|Relationship - Father|Finding|false|false||father
null|Father - courtesy title|Finding|false|false||fathernull|Father (person)|Subject|false|false||fathernull|Benign Meningioma|Disorder|false|false||meningioma
null|Meningioma|Disorder|false|false||meningiomanull|Following|Time|false|false||subsequentnull|Seizures|Finding|false|false||seizuresnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Gen
null|GEN1 wt Allele|Finding|false|false||Gen
null|GEN1 gene|Finding|false|false||Gennull|Lying in bed|Modifier|false|false||Lying in bednull|Telling untruths|Finding|false|false||Lyingnull|Supine Position|Modifier|false|false||Lyingnull|BORNHOLM EYE DISEASE|Disorder|false|false||bednull|Bachelor of Education|Finding|false|false||bednull|Beds|Device|false|false||bednull|Patient Location - Bed|Modifier|false|false||bednull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|HEENT|Anatomy|false|false||HEENTnull|Moist oral mucosa|Finding|false|false||moist oral mucosanull|Moist|Modifier|false|false||moistnull|Oral mucous membrane structure|Anatomy|false|false||oral mucosanull|Oral Dosage Form|Drug|false|false||oralnull|Oral Route of Administration|Finding|false|false||oral
null|Oral (intended site)|Finding|false|false||oralnull|Oral cavity|Anatomy|false|false||oralnull|Oral|Modifier|false|false||oralnull|null|Finding|false|false||mucosanull|Mucous Membrane|Anatomy|false|false||mucosanull|Passive joint movement of neck (finding)|Finding|false|false||Neck
null|Neck problem|Finding|false|false||Necknull|dendritic spine neck|Anatomy|false|false||Neck
null|Neck|Anatomy|false|false||Necknull|Emotional tenderness|Finding|true|false||tenderness
null|Sore to touch|Finding|true|false||tendernessnull|Palpation|Procedure|false|false||palpationnull|Rupture of Membranes|Finding|false|false||ROM
null|ROM1 gene|Finding|false|false||ROMnull|Range of motion technique (procedure)|Procedure|false|false||ROMnull|Read Only Memory Device|Device|false|false||ROMnull|Romani Language|Entity|false|false||ROMnull|Supple|Finding|false|false||supplenull|Carotid Arteries|Anatomy|false|false||carotidnull|Bone structure of spine|Anatomy|false|false||vertebralnull|Bruit|Finding|false|false||bruitnull|Heart murmur|Finding|true|false||murmursnull|Pericardial friction rub|Finding|true|false||rubsnull|Lung diseases|Disorder|false|false||Lungnull|Lung Problem|Finding|false|false||Lungnull|Chest>Lung|Anatomy|false|false||Lung
null|Lung|Anatomy|false|false||Lungnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Auscultation|Procedure|false|false||auscultationnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false||aBdnull|ABD (body structure)|Anatomy|false|false||aBd
null|Abdomen|Anatomy|false|false||aBdnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|Hereditary Multiple Exostoses|Disorder|false|false||extnull|EXT1 wt Allele|Finding|false|false||ext
null|EXT1 gene|Finding|false|false||extnull|Relational Operator - Equal|Finding|false|false||equalnull|Equal|Modifier|false|false||equalnull|Radial|Finding|false|false||radial
null|Circumpennate|Finding|false|false||radialnull|Pedal pulse|Finding|false|false||pedal pulsesnull|Foot|Anatomy|false|false||pedal
null|Paw|Anatomy|false|false||pedalnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Neurologic Examination|Procedure|false|false||Neurologic examinationnull|Neurologic (qualifier value)|Modifier|false|false||Neurologicnull|Physical Examination|Procedure|false|false||examination
null|Medical Examination|Procedure|false|false||examinationnull|Examination|Event|false|false||examinationnull|Mental state|Finding|false|false||Mental statusnull|null|Attribute|false|false||Mental status
null|null|Attribute|false|false||Mental statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|Alert brand of caffeine|Drug|false|false||alert
null|Alert brand of caffeine|Drug|false|false||alertnull|Mentally alert|Finding|false|false||alert
null|Consciousness clear|Finding|false|false||alert
null|Alert note|Finding|false|false||alert
null|Alert|Finding|false|false||alertnull|null|Attribute|false|false||alertnull|cooperative|Entity|false|false||cooperativenull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Affect (mental function)|Finding|false|false||affectnull|assessment of affect|Procedure|false|false||affectnull|Oriented to person|Finding|false|false||Oriented to personnull|Oriented to place|Finding|false|false||Orientednull|Orientation, Spatial|Modifier|false|false||Orientednull|Person Info|Finding|false|false||personnull|null|Attribute|false|false||personnull|Persons|Subject|false|false||personnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Backward (qualifier value)|Modifier|false|false||backwardsnull|Speech|Finding|false|false||Speechnull|Speech assessment|Procedure|false|false||Speechnull|Comprehension|Finding|false|false||comprehensionnull|speech fluency repetition (physical finding)|Finding|false|false||repetition
null|Repeat|Finding|false|false||repetitionnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Dysarthria|Disorder|true|false||dysarthrianull|Reading (datum presentation)|Finding|false|false||Reading
null|Reading (activity)|Finding|false|false||Reading
null|Reading Ability question|Finding|false|false||Readingnull|null|Attribute|false|false||Readingnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Confusion|Disorder|false|false||confusionnull|Clouded consciousness|Finding|false|false||confusionnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Apraxias|Disorder|true|false||apraxianull|Victim of neglect (finding)|Finding|true|false||neglectnull|Neglect (event)|Event|true|false||neglectnull|Neoplasm of uncertain or unknown behavior of cranial nerves|Disorder|false|false||Cranial Nerves
null|Benign neoplasm of cranial nerves|Disorder|false|false||Cranial Nervesnull|Cranial Nerves|Anatomy|false|false||Cranial Nervesnull|Bone structure of cranium|Anatomy|false|false||Cranialnull|Cranial|Modifier|false|false||Cranialnull|Nerve|Anatomy|false|false||Nervesnull|Pupil|Anatomy|false|false||Pupilsnull|Round shape|Modifier|false|false||roundnull|Reactive to light|Finding|false|false||reactive to lightnull|Reactive Therapy|Procedure|false|false||reactivenull|Reactive|Modifier|false|false||reactivenull|TNFSF14 protein, human|Drug|false|false||light
null|TNFSF14 protein, human|Drug|false|false||lightnull|Light - subjective measurement|Finding|false|false||light
null|TNFSF14 wt Allele|Finding|false|false||light
null|TNFSF14 gene|Finding|false|false||light
null|Light color|Finding|false|false||lightnull|Phototherapy|Procedure|false|false||lightnull|Light|Phenomenon|false|false||lightnull|Light (qualifier)|Modifier|false|false||lightnull|Visual Fields|Modifier|false|false||Visual fieldsnull|Visual|Finding|false|false||Visualnull|Full|Modifier|false|false||fullnull|Social confrontation skill|Finding|false|false||confrontationnull|Confrontation visual field test|Procedure|false|false||confrontation
null|Confrontation|Procedure|false|false||confrontationnull|Retina|Anatomy|false|false||Retinasnull|Sharp sensation quality|Finding|false|false||sharp
null|SPEN wt Allele|Finding|false|false||sharp
null|SPEN gene|Finding|false|false||sharpnull|Disk Drug Form|Drug|false|false||discnull|Disc (List bullets)|Finding|false|false||disc
null|Discontinued|Finding|false|false||discnull|Disc - Body Part|Anatomy|false|false||disc
null|death-inducing signaling complex location|Anatomy|false|false||discnull|Disk Device|Device|false|false||discnull|Disk Shape|Modifier|false|false||discnull|Disk Dosing Unit|LabModifier|false|false||discnull|examination of extraocular movements|Procedure|false|false||Extraocular movementsnull|Extraocular|Finding|false|false||Extraocularnull|Movement|Finding|false|false||movementsnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Nystagmus|Disorder|true|false||nystagmusnull|Observation of Sensation|Finding|false|false||Sensation
null|Sensory perception|Finding|false|false||Sensationnull|sensory exam|Procedure|false|false||Sensationnull|Sensation quality|Modifier|false|false||Sensationnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Face|Anatomy|false|false||Facialnull|Facial|Modifier|false|false||Facialnull|Movement|Finding|false|false||movementnull|Symmetric Relationship|Finding|false|false||symmetric
null|Symmetrical|Finding|false|false||symmetricnull|outcomes otolaryngology hearing|Finding|false|false||Hearing
null|Hearing finding|Finding|false|false||Hearing
null|Hearing|Finding|false|false||Hearingnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Upper extremity>Finger|Anatomy|false|false||finger
null|Fingers|Anatomy|false|false||finger
null|Fingers not including thumb|Anatomy|false|false||fingernull|Palate|Anatomy|false|false||Palatenull|Elevation procedure|Procedure|false|false||elevationnull|Elevation|Modifier|false|false||elevationnull|Symmetrical|Finding|false|false||symmetricalnull|Structure of sternocleidomastoid muscle|Anatomy|false|false||Sternocleidomastoidnull|Structure of trapezius muscle|Anatomy|false|false||trapeziusnull|tongue midline|Finding|false|false||Tongue midlinenull|Benign neoplasm of tongue|Disorder|false|false||Tonguenull|Procedure on tongue|Procedure|false|false||Tonguenull|Tongue|Anatomy|false|false||Tonguenull|midline cell component|Anatomy|false|false||midlinenull|Midline (qualifier value)|Modifier|false|false||midlinenull|Movement|Finding|false|false||movementsnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|motor movement|Finding|false|false||Motornull|Motor Device|Device|false|false||Motornull|Bulk (conceptual)|Drug|false|false||bulk
null|Dietary Fiber|Drug|false|false||bulknull|Myoclonus|Finding|true|false||myoclonusnull|Tremor|Finding|false|false||tremornull|Pronator drift|Finding|true|false||pronator driftnull|Double-Expressor Lymphoma|Disorder|false|false||Del
null|Chromosome Deletion|Disorder|false|false||Del
null|Deletion Mutation|Disorder|false|false||Delnull|Delaware Language|Entity|false|false||Delnull|Bistris|Drug|false|false||Tri Binull|TRI-AAT9-1 gene|Finding|false|false||Tri
null|Temptation and Restraint Inventory|Finding|false|false||Trinull|Observation of Sensation|Finding|false|false||Sensation
null|Sensory perception|Finding|false|false||Sensationnull|sensory exam|Procedure|false|false||Sensationnull|Sensation quality|Modifier|false|false||Sensationnull|Gender Status - Intact|Finding|false|false||Intactnull|Intact|Modifier|false|false||Intactnull|Light touch|Finding|false|false||light touchnull|TNFSF14 protein, human|Drug|false|false||light
null|TNFSF14 protein, human|Drug|false|false||lightnull|Light - subjective measurement|Finding|false|false||light
null|TNFSF14 wt Allele|Finding|false|false||light
null|TNFSF14 gene|Finding|false|false||light
null|Light color|Finding|false|false||lightnull|Phototherapy|Procedure|false|false||lightnull|Light|Phenomenon|false|false||lightnull|Light (qualifier)|Modifier|false|false||lightnull|Touch Perception|Finding|false|false||touch
null|Touch sensation|Finding|false|false||touchnull|Therapeutic Touch|Procedure|false|false||touchnull|Tactile|Modifier|false|false||touchnull|Proprioception|Finding|false|false||proprioceptionnull|Observation of reflex|Finding|false|false||Reflexes
null|Reflex action|Finding|false|false||Reflexesnull|Examination of reflexes|Procedure|false|false||Reflexesnull|Symmetric Relationship|Finding|false|false||symmetric
null|Symmetrical|Finding|false|false||symmetricnull|Lower extremity>Toes|Anatomy|false|false||Toes
null|Toes|Anatomy|false|false||Toesnull|Coordination of Benefits - Coordination|Finding|false|false||Coordination
null|Coordinated|Finding|false|false||Coordination
null|Physiologic Coordination|Finding|false|false||Coordinationnull|Upper extremity>Finger|Anatomy|false|false||finger
null|Fingers|Anatomy|false|false||finger
null|Fingers not including thumb|Anatomy|false|false||fingernull|Upper extremity>Finger|Anatomy|false|false||finger
null|Fingers|Anatomy|false|false||finger
null|Fingers not including thumb|Anatomy|false|false||fingernull|Heel|Anatomy|false|false||heelnull|Shin|Anatomy|false|false||shinnull|rams|Entity|false|false||RAMsnull|Gait|Finding|false|false||Gaitnull|Narrow face|Finding|false|false||Narrownull|Narrow|Modifier|false|false||Narrow
null|Narrowed structure|Modifier|false|false||Narrownull|Steady|Modifier|false|false||steadynull|Able (qualifier value)|Finding|false|false||Ablenull|Ability|Subject|false|false||Ablenull|Walking (function)|Finding|false|false||walknull|Has difficulty doing (qualifier value)|Finding|false|false||difficultynull|Facial Hemiatrophy|Disorder|false|false||Rombergnull|Rh Negative Blood Group|Finding|false|false||Negative
null|Negative|Finding|false|false||Negative
null|Negative Finding|Finding|false|false||Negativenull|Expression Negative|Lab|false|false||Negativenull|Negative - qualifier|Modifier|false|false||Negative
null|Negative Charge|Modifier|false|false||Negativenull|Negative Number|LabModifier|false|false||Negativenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Maxillary left first molar mesial prosthesis|Device|false|false||14PMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Monos|Drug|false|false||Monos
null|Mono-S|Drug|false|false||Monos
null|Monos|Drug|false|false||Monosnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||Eos
null|Familial eosinophilia|Disorder|false|false||Eosnull|PRSS33 gene|Finding|false|false||Eos
null|IKZF4 gene|Finding|false|false||Eosnull|Eos <Loriini>|Entity|false|false||Eosnull|Maxillary left first molar mesial prosthesis|Device|false|false||14PMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Maxillary left first molar mesial prosthesis|Device|false|false||14PMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||ASTnull|Atypical Spitz Nevus|Disorder|false|false||ASTnull|SLC17A5 wt Allele|Finding|false|false||AST
null|SLC17A5 gene|Finding|false|false||AST
null|GOT1 gene|Finding|false|false||ASTnull|Asterion|Anatomy|false|false||ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Creatine Kinase|Drug|false|false||CPK
null|Creatine Kinase|Drug|false|false||CPKnull|PIK3C2A gene|Finding|false|false||CPKnull|Creatine kinase measurement|Procedure|false|false||CPKnull|Alkaline Phosphatase|Drug|false|false||AlkPhos
null|Alkaline Phosphatase|Drug|false|false||AlkPhosnull|Maxillary left first molar mesial prosthesis|Device|false|false||14PMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MB
null|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MBnull|creatine kinase activity|Finding|false|false||CK-MBnull|Serum creatine phosphokinase MB isoenzyme measurement|Procedure|false|false||CK-MB
null|Creatine kinase MB measurement|Procedure|false|false||CK-MBnull|Maxillary left first molar mesial prosthesis|Device|false|false||14PMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Albumin|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumin|Drug|false|false||Albuminnull|Albumin metabolic function|Finding|false|false||Albumin
null|ALB gene|Finding|false|false||Albuminnull|Albumin measurement|Procedure|false|false||Albuminnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Glycosylated hemoglobin A|Drug|false|false||HbA1c
null|Glycosylated hemoglobin A|Drug|false|false||HbA1cnull|Glucohemoglobin measurement|Procedure|false|false||HbA1cnull|Maxillary left first molar mesial prosthesis|Device|false|false||14PMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Arylsulfatase A, human|Drug|false|false||ASA
null|Arylsulfatase A, human|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASAnull|ARSA gene|Finding|false|false||ASAnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|CNS depressants ethanol|Drug|false|false||Ethanol
null|CNS depressants ethanol|Drug|false|false||Ethanol
null|antiseptics ethanol|Drug|false|false||Ethanol
null|antiseptics ethanol|Drug|false|false||Ethanol
null|ethanol|Drug|false|false||Ethanol
null|ethanol|Drug|false|false||Ethanolnull|Toxic effect of ethyl alcohol|Disorder|false|false||Ethanolnull|Ethanol measurement|Procedure|false|false||Ethanolnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Radiology report|Finding|false|false||Radiology Reportnull|radiology referral type|Finding|false|false||Radiology
null|Radiology Section ID|Finding|false|false||Radiology
null|Encounter due to radiological examination|Finding|false|false||Radiologynull|Radiology studies|Procedure|false|false||Radiology
null|Diagnostic radiologic examination|Procedure|false|false||Radiology
null|Radiographic imaging procedure|Procedure|false|false||Radiologynull|Radiology Specialty|Title|false|false||Radiologynull|Report (document)|Finding|false|false||Reportnull|Reporting|Procedure|false|false||Reportnull|null|Attribute|false|false||Reportnull|tocilizumab|Drug|false|false||MRA
null|tocilizumab|Drug|false|false||MRA
null|tocilizumab|Drug|false|false||MRAnull|Magnetic Resonance Angiography|Procedure|false|false||MRAnull|MRI-Based Angiogram|Lab|false|false||MRAnull|Brain Diseases|Disorder|false|false||BRAINnull|Head>Brain|Anatomy|false|false||BRAIN
null|Brain|Anatomy|false|false||BRAINnull|Contrast Media|Drug|false|false||CONTRASTnull|Contrast|Modifier|false|false||CONTRASTnull|Study Object|Finding|false|false||Studynull|Scientific Study|Procedure|false|false||Study
null|Study|Procedure|false|false||Study
null|Clinical Research|Procedure|false|false||Studynull|Room of building - Study|Device|false|false||Studynull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|false|false||acutenull|Intracranial Route of Administration|Finding|false|false||intracranialnull|Intracranial|Anatomy|false|false||intracranialnull|Congenital Abnormality|Disorder|true|false||abnormalitynull|Abnormality|Finding|true|false||abnormalitynull|Evidence of (contextual qualifier)|Finding|false|false||evidence ofnull|Evidence|Finding|false|false||evidencenull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Act Relationship Subset - previous|Time|false|false||previous
null|Previous|Time|false|false||previousnull|Ischemic|Finding|false|false||ischemicnull|Event|Event|false|false||eventnull|Bone structure of cranium|Anatomy|false|false||cranialnull|Cranial|Modifier|false|false||cranialnull|Neck|Anatomy|false|false||cervicalnull|Cervical|Modifier|false|false||cervicalnull|tocilizumab|Drug|false|false||MRA
null|tocilizumab|Drug|false|false||MRA
null|tocilizumab|Drug|false|false||MRAnull|Magnetic Resonance Angiography|Procedure|false|false||MRAnull|MRI-Based Angiogram|Lab|false|false||MRAnull|Significant|Finding|true|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Mural|Modifier|false|false||muralnull|Flow|Phenomenon|false|false||flownull|Stenosis|Finding|false|false||stenosisnull|Stenosis <Pimeliinae>|Entity|false|false||stenosisnull|Stenosis Morphology|Modifier|false|false||stenosisnull|Woman|Subject|false|false||woman
null|Human, Female adult|Subject|false|false||womannull|Cancer patients and suicide and depression|Disorder|false|false||depression
null|Mental Depression|Disorder|false|false||depression
null|Depressive disorder|Disorder|false|false||depression
null|Depressed mood|Disorder|false|false||depressionnull|Depression - motion|Finding|false|false||depression
null|null|Finding|false|false||depressionnull|Depression - recess|Modifier|false|false||depressionnull|Gastroesophageal reflux disease|Disorder|false|false||GERDnull|Migraine Disorders|Disorder|false|false||migrainesnull|Episode of|Time|false|false||episode ofnull|Episode of|Time|false|false||episodenull|Numbness of face|Finding|false|false||facial numbnessnull|Face|Anatomy|false|false||facialnull|Facial|Modifier|false|false||facialnull|Numbness|Finding|false|false||numbness
null|Hypesthesia|Finding|false|false||numbnessnull|Numbness of face|Finding|false|false||Facial numbnessnull|Face|Anatomy|false|false||Facialnull|Facial|Modifier|false|false||Facialnull|Numbness|Finding|false|false||numbness
null|Hypesthesia|Finding|false|false||numbnessnull|Episode of|Time|false|false||episodenull|Headache|Finding|false|false||headachenull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Migraine Disorders|Disorder|false|false||migrainenull|Equal|Modifier|false|false||equivalentnull|Equivalent Weight|LabModifier|false|false||equivalentnull|Episode of|Time|false|false||episodenull|Transient Cerebral Ischemia|Disorder|false|false||TIA
null|Transient Ischemic Attack|Disorder|false|false||TIAnull|Tacca leontopetaloides|Entity|false|false||TIAnull|Thalamic structure|Anatomy|false|false||thalamusnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|Aspects of signs|Finding|true|false||signs
null|Physical findings|Finding|true|false||signsnull|Manufactured sign|Device|true|false||signsnull|Ischemia|Finding|true|false||ischemianull|Ischemia Procedure|Procedure|true|false||ischemianull|Vasculature|Anatomy|false|false||vasculaturenull|Blood supply aspects|Modifier|false|false||vasculaturenull|Migraine Disorders|Disorder|false|false||migrainenull|Much|Finding|false|false||muchnull|More|LabModifier|false|false||morenull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Diagnosis Classification - Diagnosis|Finding|false|false||diagnosis
null|diagnosis aspects|Finding|false|false||diagnosisnull|Diagnosis|Procedure|false|false||diagnosisnull|null|Attribute|false|false||diagnosisnull|Transient Cerebral Ischemia|Disorder|false|false||TIA
null|Transient Ischemic Attack|Disorder|false|false||TIAnull|Tacca leontopetaloides|Entity|false|false||TIAnull|Daily|Time|false|false||dailynull|aspirin|Drug|false|false||aspirin
null|aspirin|Drug|false|false||aspirinnull|Future|Time|false|false||futurenull|Cerebrovascular accident|Disorder|false|false||strokenull|Stroke (heart beat)|Finding|false|false||strokenull|Prophylactic treatment|Procedure|false|false||prophylaxisnull|prevention & control|Modifier|false|false||prophylaxisnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|On discharge|Time|false|false||on dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Symmetric Relationship|Finding|false|false||symmetric
null|Symmetrical|Finding|false|false||symmetricnull|Hyperreflexia|Finding|false|false||hyperreflexianull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|Neurologic Examination|Procedure|false|false||neurological examnull|Neurologic (qualifier value)|Modifier|false|false||neurologicalnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Residual|Modifier|false|false||residualnull|Sensory deficit|Finding|false|false||sensory deficitsnull|Sensory (qualifier value)|Modifier|false|false||sensorynull|Deficit|Modifier|false|false||deficitsnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|Nexium|Drug|false|false||NEXIUM
null|Nexium|Drug|false|false||NEXIUMnull|capsule (pharmacologic)|Drug|false|false||capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||capsule
null|Structure of organ capsule|Anatomy|false|false||capsulenull|Capsule Shape|Modifier|false|false||capsulenull|Capsule (unit of presentation)|LabModifier|false|false||capsule
null|Capsule Dosing Unit|LabModifier|false|false||capsulenull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Prozac|Drug|false|false||PROZAC
null|Prozac|Drug|false|false||PROZACnull|capsule (pharmacologic)|Drug|false|false||capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||capsule
null|Structure of organ capsule|Anatomy|false|false||capsulenull|Capsule Shape|Modifier|false|false||capsulenull|Capsule (unit of presentation)|LabModifier|false|false||capsule
null|Capsule Dosing Unit|LabModifier|false|false||capsulenull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|pantoprazole|Drug|false|false||Pantoprazole
null|pantoprazole|Drug|false|false||Pantoprazolenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Delayed Release Dosage Form|Drug|false|false||Delayed Releasenull|Views delayed|Attribute|false|false||Delayednull|Deferred|Time|false|false||Delayednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Delayed Release Dosage Form|Drug|false|false||Delayed Releasenull|Views delayed|Attribute|false|false||Delayednull|Deferred|Time|false|false||Delayednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Every twenty four hours|Time|false|false||Q24Hnull|24 Hours|Time|false|false||24 hoursnull|Hour|Time|false|false||hoursnull|fluoxetine|Drug|false|false||Fluoxetine
null|fluoxetine|Drug|false|false||Fluoxetinenull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Delayed Release Dosage Form|Drug|false|false||Delayed Releasenull|Views delayed|Attribute|false|false||Delayednull|Deferred|Time|false|false||Delayednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Delayed Release Dosage Form|Drug|false|false||Delayed Releasenull|Views delayed|Attribute|false|false||Delayednull|Deferred|Time|false|false||Delayednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Migraine Disorders|Disorder|false|false||Migrainenull|Mild Severity of Illness Code|Finding|false|false||Mildnull|Mild (qualifier value)|Modifier|false|false||Mild
null|Mild Allergy Severity|Modifier|false|false||Mildnull|Symmetric Relationship|Finding|false|false||symmetric
null|Symmetrical|Finding|false|false||symmetricnull|Hyperreflexia in the lower extremities|Finding|false|false||hyperreflexia in the lower extremitiesnull|Hyperreflexia|Finding|false|false||hyperreflexianull|Lower Extremity|Anatomy|false|false||lower extremitiesnull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|Neurologic Examination|Procedure|false|false||neurological examnull|Neurologic (qualifier value)|Modifier|false|false||neurologicalnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Left sided|Modifier|false|false||left sided
null|Left|Modifier|false|false||left sidednull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Numbness of face|Finding|false|false||facial numbnessnull|Face|Anatomy|false|false||facialnull|Facial|Modifier|false|false||facialnull|Numbness|Finding|false|false||numbness
null|Hypesthesia|Finding|false|false||numbnessnull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|Aspects of signs|Finding|true|false||signs
null|Physical findings|Finding|true|false||signsnull|Manufactured sign|Device|true|false||signsnull|Ischemia|Finding|true|false||ischemianull|Ischemia Procedure|Procedure|true|false||ischemianull|Relate - vinyl resin|Drug|false|false||relatednull|Role Link Type - related|Finding|false|false||related
null|Related (finding)|Finding|false|false||relatednull|Definitely Related to Intervention|Modifier|false|false||related
null|Relationships|Modifier|false|false||relatednull|Migraine Disorders|Disorder|false|false||migraine headachesnull|Migraine Disorders|Disorder|false|false||migrainenull|Headache|Finding|false|false||headachesnull|Full|Modifier|false|false||fullnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|aspirin|Drug|false|false||aspirin
null|aspirin|Drug|false|false||aspirinnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Numbness|Finding|false|false||numbness
null|Hypesthesia|Finding|false|false||numbnessnull|Weakness|Finding|false|false||weakness
null|Asthenia|Finding|false|false||weaknessnull|Headache|Finding|false|false||headachesnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Proximal|Modifier|false|false||nearestnull|Further|Modifier|false|false||furthernull|Processing type - Evaluation|Finding|false|false||evaluationnull|Evaluation procedure|Procedure|false|false||evaluation
null|Evaluation|Procedure|false|false||evaluationnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions