CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Level of Care - Surgery|Finding|false|false||SURGERY
null|Surgical procedure finding|Finding|false|false||SURGERY
null|Surgical aspects|Finding|false|false||SURGERYnull|Operative Surgical Procedures|Procedure|false|false||SURGERYnull|General surgery specialty|Title|false|false||SURGERY
null|Surgery specialty|Title|false|false||SURGERYnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Dyes|Drug|false|false||Dyenull|Iodine, Homeopathic preparation|Drug|false|false||Iodine
null|iodine|Drug|false|false||Iodine
null|iodine|Drug|false|false||Iodine
null|iodine|Drug|false|false||Iodinenull|Containing (qualifier value)|Finding|false|false||Containingnull|Contain (action)|Event|false|false||Containingnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Chief complaint (finding)|Finding|false|false||Chief Complaintnull|Complaint (finding)|Finding|false|false||Complaintnull|null|Attribute|false|false||Complaintnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Vomiting|Finding|false|false||vomitingnull|1 Day|Time|false|false||1 daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|History of present illness (finding)|Finding|false|false||History of Present Illnessnull|null|Attribute|false|false||History of Present Illnessnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Present illness|Finding|false|false||Present Illnessnull|Present|Finding|false|false||Present
null|Presentation|Finding|false|false||Presentnull|Illness (finding)|Finding|false|false||Illnessnull|Sigmoid colectomy|Procedure|false|false|C0227391|sigmoid colectomynull|Sigmoid colon|Anatomy|false|false|C0009274;C0012813;C0192866|sigmoidnull|Colectomy|Procedure|false|false|C0227391|colectomynull|Recurrent|Time|false|false||recurrent
null|Episodic|Time|false|false||recurrentnull|Diverticulitis|Disorder|false|false|C0227391|diverticulitisnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Low residue diet|Procedure|false|false||low residue dietnull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Residue|Finding|false|false||residuenull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|Wound Infection|Finding|false|false||wound infectionnull|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic Wound|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|1 Week|Time|false|false||one weeknull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|1 Day|Time|false|false||1 daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|With intensity|Modifier|false|false||intensenull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Emesis [PE]|Finding|false|false||emesis
null|Vomiting|Finding|false|false||emesis
null|Vomitus|Finding|false|false||emesisnull|Emesis <Emesidini>|Entity|false|false||emesis
null|Emesis <subgenus>|Entity|false|false||emesisnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Intensity and Distress 1|Finding|false|false||slightnull|Slight (qualifier value)|Modifier|false|false||slight
null|Mild (qualifier value)|Modifier|false|false||slightnull|Increase|Finding|false|false||increasenull|Epigastric pain|Finding|false|false|C0521440;C0000726|epigastric abdominal painnull|Epigastric|Anatomy|false|false|C0232493|epigastricnull|Abdominal Pain|Finding|false|false|C0000726|abdominal painnull|Abdomen|Anatomy|false|false|C0000737;C1549543;C0030193;C0232493|abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Administration Method - Pain|Finding|false|false|C0000726|pain
null|Pain|Finding|false|false|C0000726|painnull|null|Attribute|false|false||painnull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Emotional tenderness|Finding|false|false||tenderness
null|Sore to touch|Finding|false|false||tendernessnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Diverticulitis|Disorder|false|false||diverticulitisnull|ACP2 protein, human|Drug|false|false||lap
null|ACP2 protein, human|Drug|false|false||lapnull|Congenital laryngeal adductor palsy|Disorder|false|false|C0227391|lapnull|Left atrial pressure|Finding|false|false|C0227391|lap
null|ACP2 gene|Finding|false|false|C0227391|lap
null|PICALM wt Allele|Finding|false|false|C0227391|lap
null|LAP3 wt Allele|Finding|false|false|C0227391|lap
null|ACP2 wt Allele|Finding|false|false|C0227391|lap
null|LAP3 gene|Finding|false|false|C0227391|lap
null|CENPJ gene|Finding|false|false|C0227391|lap
null|CEBPB wt Allele|Finding|false|false|C0227391|lap
null|PICALM gene|Finding|false|false|C0227391|lap
null|CEBPB gene|Finding|false|false|C0227391|lapnull|Laparoscopy|Procedure|false|false|C0227391|lapnull|Lap - unit|LabModifier|false|false||lapnull|Sigmoid colectomy|Procedure|false|false|C0227391|sigmoid colectomynull|Sigmoid colon|Anatomy|false|false|C0396060;C0456170;C1424863;C1425522;C1423544;C1413323;C2827449;C5575443;C3540509;C5890955;C1412132;C0031150;C0009274;C0192866|sigmoidnull|Colectomy|Procedure|false|false|C0227391|colectomynull|Wound Infection|Finding|false|false||wound infectionnull|Traumatic Wound|Disorder|false|false||wound
null|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Migraine Disorders|Disorder|false|false||Migrainesnull|Table Cell Horizontal Align - left|Finding|false|false|C4299059;C0851278;C0016129|Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Upper extremity>Finger|Anatomy|false|false|C0007642;C1552822;C2025995|finger
null|Fingers|Anatomy|false|false|C0007642;C1552822;C2025995|finger
null|Fingers not including thumb|Anatomy|false|false|C0007642;C1552822;C2025995|fingernull|Cellulitis|Disorder|false|false|C4299059;C0851278;C0016129|cellulitisnull|cellulitis on exam (physical finding)|Finding|false|false|C4299059;C0851278;C0016129|cellulitisnull|Social and personal history|Finding|false|false||Social History
null|Social History|Finding|false|false||Social Historynull|Social|Finding|false|false||Socialnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Family Medical History|Finding|false|false||Family Historynull|Entity Name Part Type - family|Finding|false|false||Family
null|Last Name|Finding|false|false||Family
null|Living Arrangement - Family|Finding|false|false||Family
null|Family (taxonomic)|Finding|false|false||Family
null|Family Collection|Finding|false|false||Familynull|Family|Subject|false|false||Familynull|History of present illness (finding)|Finding|false|true||History
null|History of previous events|Finding|false|true||History
null|Historical aspects qualifier|Finding|false|true||History
null|Medical History|Finding|false|true||History
null|Concept History|Finding|false|true||Historynull|History|Subject|false|false||Historynull|Indirect exposure mechanism - Father|Finding|false|false||father
null|Relationship - Father|Finding|false|false||father
null|Father - courtesy title|Finding|false|false||fathernull|Father (person)|Subject|false|false||fathernull|Colitis|Disorder|false|false||colitisnull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|Apyrexial|Finding|false|false||afebrilenull|Taking vital signs|Procedure|false|false||vital signsnull|null|Attribute|false|false||vital signs
null|Vital signs|Attribute|false|false||vital signsnull|Vital High Nitrogen Enteral Nutrition|Drug|false|false||vitalnull|Vital (qualifier value)|Modifier|false|false||vitalnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|null|Finding|false|false||within normal limitsnull|Limited (extensiveness)|Finding|false|false||limitsnull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|talkative|Finding|false|false||talkativenull|Extraocular|Finding|false|false|C0028863|EOMnull|Muscle of orbit|Anatomy|false|false|C0241886;C1642390;C0205180|EOMnull|Full|Modifier|false|false||fullnull|Pupil equal round and reacting to light|Finding|false|false|C0028863|PERRLnull|Anicteric|Finding|false|false|C0028863;C0036410|anictericnull|Scleral Diseases|Disorder|false|false|C0036410|scleranull|examination of sclera|Procedure|false|false|C0036410|scleranull|Sclera|Anatomy|false|false|C2228481;C0036412;C0205180|scleranull|chest clear|Finding|false|false|C1527391;C0817096|Chest clearnull|Chest problem|Finding|false|false|C1527391;C0817096|Chestnull|Chest|Anatomy|false|false|C0578395;C0741025;C1550016|Chest
null|Anterior thoracic region|Anatomy|false|false|C0578395;C0741025;C1550016|Chestnull|Remote control command - Clear|Finding|false|false|C1527391;C0817096|clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Heart murmur|Finding|true|false||murmursnull|Abdomen soft|Finding|false|false|C0230168;C0000726|Abdomen softnull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|Abdomennull|Abdomen problem|Finding|false|false|C0230168;C0000726|Abdomennull|Abdomen|Anatomy|false|false|C0941288;C0426663;C3542022;C0153662|Abdomen
null|Abdominal Cavity|Anatomy|false|false|C0941288;C0426663;C3542022;C0153662|Abdomennull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false|C0230168;C0000726|softnull|Soft|Modifier|false|false||softnull|Round shape|Modifier|false|false||roundnull|Open|Modifier|false|false||opennull|Transverse incision|Procedure|false|false|C0222331;C0278403;C2338258|transverse incisionnull|Anatomical transverse plane|Modifier|false|false||transverse
null|Transverse plane|Modifier|false|false||transversenull|Surgical wound|Disorder|false|false|C2338258;C0222331;C0278403|incisionnull|Surgical incisions|Procedure|false|false|C0222331;C0278403;C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0332803;C0184898;C1261209|incisionnull|Subcutaneous Tissue|Anatomy|false|false|C0184898;C0332803;C1554187;C1261209|subcutis
null|Subcutaneous Fat|Anatomy|false|false|C0184898;C0332803;C1554187;C1261209|subcutisnull|Gender Status - Intact|Finding|false|false|C0222331;C0278403|intactnull|Intact|Modifier|false|false||intactnull|Deep Resection Margin|Attribute|false|false||deepnull|Deep (qualifier value)|Modifier|false|false||deepnull|Fascia|Anatomy|false|false||fascianull|Erythema|Disorder|true|false||erythemanull|Induration|Finding|true|false||indurationnull|Minimal|Modifier|false|false||minimal
null|Mild (qualifier value)|Modifier|false|false||minimal
null|Minimum|Modifier|false|false||minimalnull|Serous|Modifier|false|false||serousnull|system output|Finding|false|false||outputnull|Measurement of fluid output|Procedure|false|false||outputnull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Computed tomography, abdomen; without contrast material|Procedure|false|false|C0230168;C0000726|CT ABDOMEN W/O CONTRASTnull|CT of abdomen|Procedure|false|false|C0230168;C0000726|CT ABDOMENnull|null|Attribute|false|false|C0230168;C0000726|CT ABDOMENnull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|ABDOMENnull|Abdomen problem|Finding|false|false|C0230168;C0000726|ABDOMENnull|Abdomen|Anatomy|false|false|C0941288;C0153662;C0202838;C1644645;C0412620|ABDOMEN
null|Abdominal Cavity|Anatomy|false|false|C0941288;C0153662;C0202838;C1644645;C0412620|ABDOMENnull|Contrast Media|Drug|false|false||CONTRASTnull|Contrast|Modifier|false|false||CONTRASTnull|Contrast Media|Drug|false|false||CONTRASTnull|Contrast|Modifier|false|false||CONTRASTnull|Computed tomography of pelvis|Procedure|false|false|C4266535;C0030797;C0559769|CT PELVISnull|null|Attribute|false|false|C4266535;C0030797;C0559769|CT PELVISnull|Malignant neoplasm of pelvis|Disorder|false|false|C4266535;C0030797;C0559769|PELVISnull|Pelvis problem|Finding|false|false|C4266535;C0030797;C0559769|PELVISnull|Pelvis+|Anatomy|false|false|C0812455;C0153663;C0882057;C0412628|PELVIS
null|Pelvic cavity structure|Anatomy|false|false|C0812455;C0153663;C0882057;C0412628|PELVIS
null|Pelvis|Anatomy|false|false|C0812455;C0153663;C0882057;C0412628|PELVISnull|Contrast Media|Drug|false|false||CONTRASTnull|Contrast|Modifier|false|false||CONTRASTnull|Indication of (contextual qualifier)|Finding|false|false||Reasonnull|Abscess|Disorder|false|false||abscessnull|null|Finding|false|false||abscessnull|IV contrast|Drug|true|false||IV contrastnull|Contrast Media|Drug|true|false||contrastnull|Contrast|Modifier|false|false||contrastnull|Field of View|Modifier|false|false||Field of viewnull|Knowledge Field|Finding|false|false||Field
null|Force Field|Finding|false|false||Field
null|Field|Finding|false|false||Fieldnull|field - patient encounter|Procedure|false|false||Fieldnull|View|Modifier|false|false||viewnull|Medical Condition|Finding|false|false||MEDICAL CONDITIONnull|Medical referral type|Finding|false|false||MEDICAL
null|Medical|Finding|false|false||MEDICAL
null|Medical school type|Finding|false|false||MEDICALnull|Medical service|Procedure|false|false||MEDICALnull|Disease|Disorder|false|false||CONDITIONnull|Logical Condition|Finding|false|false||CONDITIONnull|null|Attribute|false|false||CONDITIONnull|Condition|Modifier|false|false||CONDITIONnull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Old|Time|false|false||oldnull|Woman|Subject|false|false||woman
null|Human, Female adult|Subject|false|false||womannull|Colectomy|Procedure|false|false||colectomynull|Elevated|Modifier|false|false||elevated
null|High|Modifier|false|false||elevatednull|Leukocytes|Anatomy|false|false|C0027497|WBCnull|Nausea|Finding|false|false|C0023516|nauseanull|null|Attribute|false|false||nauseanull|Indication of (contextual qualifier)|Finding|false|false||REASON FORnull|Indication of (contextual qualifier)|Finding|false|false||REASONnull|Physical Examination|Procedure|false|false||EXAMINATION
null|Medical Examination|Procedure|false|false||EXAMINATIONnull|Examination|Event|false|false||EXAMINATIONnull|Abscess|Disorder|false|false||abscessnull|null|Finding|false|false||abscessnull|IV contrast|Drug|true|false||IV contrastnull|Contrast Media|Drug|true|false||contrastnull|Contrast|Modifier|false|false||contrastnull|Medical contraindication|Finding|false|false||CONTRAINDICATIONSnull|IV contrast|Drug|false|false||IV CONTRASTnull|Contrast Media|Drug|false|false||CONTRASTnull|Contrast|Modifier|false|false||CONTRASTnull|Indication of (contextual qualifier)|Finding|false|false||INDICATION
null|Indication|Finding|false|false||INDICATIONnull|null|Attribute|false|false||INDICATIONnull|Woman|Subject|false|false||woman
null|Human, Female adult|Subject|false|false||womannull|Elevated|Modifier|false|false||elevated
null|High|Modifier|false|false||elevatednull|Leukocytes|Anatomy|false|false|C0851353;C1413336;C1413337|white blood cellnull|White (population group)|Subject|false|false||white
null|Caucasian|Subject|false|false||white
null|Caucasians|Subject|false|false||whitenull|White color|Modifier|false|false||whitenull|Blood Cells|Anatomy|false|false||blood cellnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516;C0007634|bloodnull|peripheral blood|Finding|false|false|C0007634|blood
null|Blood|Finding|false|false|C0007634|blood
null|In Blood|Finding|false|false|C0007634|bloodnull|CELP gene|Finding|false|false|C0023516;C0007634|cell
null|CEL gene|Finding|false|false|C0023516;C0007634|cellnull|Cells|Anatomy|false|false|C0005768;C0229664;C0005767;C1413336;C1413337;C0851353|cellnull|Cell Device|Device|false|false||cell
null|Cellular Phone|Device|false|false||cellnull|Cell (compartment)|Modifier|false|false||cellnull|Count Dosing Unit|LabModifier|false|false||count
null|Count|LabModifier|false|false||countnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Recent|Time|false|false||recentnull|Colectomy|Procedure|false|false||colectomynull|Recurrent|Time|false|false||recurrent
null|Episodic|Time|false|false||recurrentnull|Diverticulitis|Disorder|false|false||diverticulitisnull|Comparison|Event|false|false||COMPARISONnull|null|Attribute|false|false|C4266535;C0030797;C0559769|CT abdomen and pelvisnull|CT of abdomen|Procedure|false|false|C0000726;C1508499;C0230168;C0000726;C4266535;C0030797;C0559769|CT abdomennull|null|Attribute|false|false|C0230168;C0000726|CT abdomennull|Abdominopelvic structure|Anatomy|false|false|C0153662;C0412620|abdomen and pelvisnull|Abdomen|Anatomy|false|false|C0412620|abdomen andnull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726;C1508499|abdomennull|Abdomen problem|Finding|false|false|C0230168;C0000726|abdomennull|Abdomen|Anatomy|false|false|C1644645;C0941288;C0153662;C0412620|abdomen
null|Abdominal Cavity|Anatomy|false|false|C1644645;C0941288;C0153662;C0412620|abdomennull|Malignant neoplasm of pelvis|Disorder|false|false|C4266535;C0030797;C0559769|pelvisnull|Pelvis problem|Finding|false|false|C4266535;C0030797;C0559769|pelvisnull|Pelvis+|Anatomy|false|false|C1715387;C0153663;C0812455;C0412620|pelvis
null|Pelvic cavity structure|Anatomy|false|false|C1715387;C0153663;C0812455;C0412620|pelvis
null|Pelvis|Anatomy|false|false|C1715387;C0153663;C0812455;C0412620|pelvisnull|Techniques|Finding|false|false||TECHNIQUEnull|Multidetector Computed Tomography|Procedure|false|false||MDCTnull|Acquired Name|Finding|false|false||acquirednull|Acquired (qualifier value)|Modifier|false|false||acquirednull|Axial|Modifier|false|false||axialnull|Abdominopelvic structure|Anatomy|false|false|C1527415;C4521986;C0009924;C0812455;C1533734;C0941288;C0153662;C0153663|abdomen and pelvisnull|Abdomen|Anatomy|false|false|C0153663;C0941288;C1527415;C4521986;C0812455;C0153662|abdomen andnull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726;C1508499;C4266535;C0030797;C0559769;C0000726|abdomennull|Abdomen problem|Finding|false|false|C0000726;C0230168;C0000726;C1508499|abdomennull|Abdomen|Anatomy|false|false|C0153662;C0812455;C0941288;C1527415;C4521986;C0153663|abdomen
null|Abdominal Cavity|Anatomy|false|false|C0153662;C0812455;C0941288;C1527415;C4521986;C0153663|abdomennull|Malignant neoplasm of pelvis|Disorder|false|false|C0000726;C4266535;C0030797;C0559769;C1508499;C0230168;C0000726|pelvisnull|Pelvis problem|Finding|false|false|C4266535;C0030797;C0559769;C0230168;C0000726;C0000726;C1508499|pelvisnull|Pelvis+|Anatomy|false|false|C0812455;C0153663;C0153662|pelvis
null|Pelvic cavity structure|Anatomy|false|false|C0812455;C0153663;C0153662|pelvis
null|Pelvis|Anatomy|false|false|C0812455;C0153663;C0153662|pelvisnull|Administration (procedure)|Procedure|false|false|C1508499|administrationnull|Administration occupational activities|Event|false|false||administrationnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896;C1508499;C0000726;C0230168;C0000726|oral
null|Oral (intended site)|Finding|false|false|C0226896;C1508499;C0000726;C0230168;C0000726|oralnull|Oral cavity|Anatomy|false|false|C1272919;C1527415;C4521986|oralnull|Oral|Modifier|false|false||oralnull|Contrast Media|Drug|false|false|C1508499|contrastnull|Contrast|Modifier|false|false||contrastnull|IV contrast|Drug|false|false||intravenous contrastnull|Intravenous Route of Administration|Finding|false|false||intravenousnull|Intravenous|Modifier|false|false||intravenousnull|Contrast Media|Drug|false|false||contrastnull|Contrast|Modifier|false|false||contrastnull|findings aspects|Finding|false|false||FINDINGSnull|null|Attribute|false|false||FINDINGSnull|Lung diseases|Disorder|false|false|C4037972;C0024109|lungnull|Lung Problem|Finding|false|false|C4037972;C0024109|lungnull|Chest>Lung|Anatomy|false|false|C0740941;C1550016;C0024115|lung
null|Lung|Anatomy|false|false|C0740941;C1550016;C0024115|lungnull|Base|Drug|false|false||basesnull|Base - unit of product usage|LabModifier|false|false||basesnull|Remote control command - Clear|Finding|false|false|C4037972;C0024109|clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Calcified granuloma|Finding|false|false||calcified granulomanull|Calcified (qualifier value)|Modifier|false|false||calcifiednull|null|Finding|false|false||granuloma
null|Granuloma|Finding|false|false||granulomanull|Structure of base of right lung|Anatomy|false|false|C1704464;C0178499;C1550601;C1880279;C0740941;C1549548;C1705938;C1843354;C1552823;C0024115;C0442739|right lung basenull|Right lung|Anatomy|false|false|C1549548;C1705938;C1843354;C0442739;C1552823;C0024115;C1704464;C0178499;C1550601;C1880279;C0740941|right lungnull|Table Cell Horizontal Align - right|Finding|false|false|C0225706;C2987514;C0225704;C0225708|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Basal segment of lung|Anatomy|false|false|C1549548;C1705938;C1843354;C0024115;C0740941;C1704464;C0178499;C1550601;C1880279;C1552823;C0442739|lung basenull|Lung diseases|Disorder|false|false|C2987514;C0225706;C0225704;C4037972;C0024109;C0225708|lungnull|Lung Problem|Finding|false|false|C0225704;C0225708;C0225706;C4037972;C0024109;C2987514|lungnull|Chest>Lung|Anatomy|false|false|C1549548;C1705938;C1843354;C0024115;C0740941;C1704464;C0178499;C1550601;C1880279|lung
null|Lung|Anatomy|false|false|C1549548;C1705938;C1843354;C0024115;C0740941;C1704464;C0178499;C1550601;C1880279|lungnull|nitrogenous base|Drug|false|false|C2987514;C0225708;C0225706;C0225704;C4037972;C0024109|base
null|Base|Drug|false|false|C2987514;C0225708;C0225706;C0225704;C4037972;C0024109|base
null|Dental Base|Drug|false|false|C2987514;C0225708;C0225706;C0225704;C4037972;C0024109|base
null|base - RoleClass|Drug|false|false|C2987514;C0225708;C0225706;C0225704;C4037972;C0024109|basenull|Base - General Qualifier|Finding|false|false|C2987514;C0225706;C0225704;C4037972;C0024109;C0225708|base
null|BPIFA4P gene|Finding|false|false|C2987514;C0225706;C0225704;C4037972;C0024109;C0225708|base
null|Base - RX Component Type|Finding|false|false|C2987514;C0225706;C0225704;C4037972;C0024109;C0225708|basenull|Anatomical base|Anatomy|false|false|C0024115;C1549548;C1705938;C1843354;C1704464;C0178499;C1550601;C1880279;C1552823;C0740941;C0442739|basenull|Base - unit of product usage|LabModifier|false|false||basenull|null|Finding|false|false|C0225706;C2987514;C0225704;C0225708|unchangednull|About The Same|Modifier|false|false||unchangednull|Limited component (foundation metadata concept)|Finding|false|false|C4037974;C0018787|Limited
null|Limited (extensiveness)|Finding|false|false|C4037974;C0018787|Limitednull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C0795691;C0439801;C3542948;C0153957;C0153500|heart
null|Heart|Anatomy|false|false|C0795691;C0439801;C3542948;C0153957;C0153500|heartnull|null|Modifier|false|false||unremarkablenull|Pericardial effusion|Disorder|true|false|C0031050;C0442031|pericardial effusionnull|Pericardial effusion body substance|Finding|true|false|C0031050;C0442031|pericardial effusionnull|Pericardial (qualifier value)|Anatomy|false|false|C2317432;C1546613;C0013687;C1253937;C0031039|pericardial
null|Pericardial sac structure|Anatomy|false|false|C2317432;C1546613;C0013687;C1253937;C0031039|pericardialnull|Effusion (substance)|Finding|true|false|C0031050;C0442031|effusion
null|null|Finding|true|false|C0031050;C0442031|effusion
null|effusion|Finding|true|false|C0031050;C0442031|effusionnull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|abdomennull|Abdomen problem|Finding|false|false|C0230168;C0000726|abdomennull|Abdomen|Anatomy|false|false|C0941288;C2032932;C0577060;C0872387;C0023895;C0496870;C0153662|abdomen
null|Abdominal Cavity|Anatomy|false|false|C0941288;C2032932;C0577060;C0872387;C0023895;C0496870;C0153662|abdomennull|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|false|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|false|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|livernull|Benign neoplasm of liver|Disorder|false|false|C0230168;C0000726;C4037986;C1278929;C0023884|liver
null|Liver diseases|Disorder|false|false|C0230168;C0000726;C4037986;C1278929;C0023884|livernull|Liver problem|Finding|false|false|C0230168;C0000726;C4037986;C1278929;C0023884|livernull|Procedures on liver|Procedure|false|false|C4037986;C1278929;C0023884;C0230168;C0000726|livernull|Abdomen>Liver|Anatomy|false|false|C0153470;C0872387;C0577060;C0812414;C0023895;C0496870;C0721399;C0023899;C2032932;C0869677|liver
null|null|Anatomy|false|false|C0153470;C0872387;C0577060;C0812414;C0023895;C0496870;C0721399;C0023899;C2032932;C0869677|liver
null|Liver|Anatomy|false|false|C0153470;C0872387;C0577060;C0812414;C0023895;C0496870;C0721399;C0023899;C2032932;C0869677|livernull|examination of gallbladder|Procedure|false|false|C4071903;C0016976;C1524055;C0230168;C0000726;C4037986;C1278929;C0023884|gallbladdernull|Abdomen>Gallbladder|Anatomy|false|false|C2032932;C0812414;C0153470;C0869677|gallbladder
null|Gallbladder|Anatomy|false|false|C2032932;C0812414;C0153470;C0869677|gallbladder
null|Gallbladder (MMHCC)|Anatomy|false|false|C2032932;C0812414;C0153470;C0869677|gallbladdernull|Malignant neoplasm of spleen|Disorder|false|false|C4037986;C1278929;C0023884;C4071903;C0016976;C1524055;C4037984;C0037993|spleennull|Spleen problem|Finding|false|false|C4071903;C0016976;C1524055;C4037984;C0037993;C4037986;C1278929;C0023884|spleennull|Procedures on Spleen|Procedure|false|false|C4037984;C0037993;C4071903;C0016976;C1524055;C4037986;C1278929;C0023884|spleennull|Abdomen>Spleen|Anatomy|false|false|C0869677;C0812414;C0153470|spleen
null|Spleen|Anatomy|false|false|C0869677;C0812414;C0153470|spleennull|Both kidneys|Anatomy|false|false||kidneys
null|Kidney|Anatomy|false|false||kidneysnull|Adrenal|Finding|false|false|C0001625|adrenalnull|Adrenal Glands|Anatomy|false|false|C0521428|adrenalnull|Gland|Anatomy|false|false|C0771711;C0869826;C1512911;C0347284;C0030286;C0577027;C0872393;C0038354;C0496905;C0153943;C0154060;C0813176|glandsnull|pancreas extract|Drug|false|false|C1285092;C4037927;C0030274|pancreas
null|pancreas extract|Drug|false|false|C1285092;C4037927;C0030274|pancreasnull|Benign tumor of pancreas|Disorder|false|false|C4037927;C0030274;C1285092|pancreas
null|Pancreatic Diseases|Disorder|false|false|C4037927;C0030274;C1285092|pancreasnull|Pancreas problem|Finding|false|false|C4037927;C0030274;C1285092|pancreasnull|Procedures on Pancreas|Procedure|false|false|C4037927;C0030274;C1285092|pancreasnull|Abdomen>Pancreas|Anatomy|false|false|C0869826;C0347284;C0030286;C0813176;C0771711|pancreas
null|Pancreas|Anatomy|false|false|C0869826;C0347284;C0030286;C0813176;C0771711|pancreasnull|Neoplasm of uncertain or unknown behavior of stomach|Disorder|false|false|C1285092;C3714551;C0038351;C4266636|stomach
null|Stomach Diseases|Disorder|false|false|C1285092;C3714551;C0038351;C4266636|stomach
null|Benign neoplasm of stomach|Disorder|false|false|C1285092;C3714551;C0038351;C4266636|stomach
null|Carcinoma in situ of stomach|Disorder|false|false|C1285092;C3714551;C0038351;C4266636|stomachnull|Stomach problem|Finding|false|false|C1285092;C3714551;C0038351;C4266636|stomachnull|Procedure on stomach|Procedure|false|false|C3714551;C0038351;C4266636;C1285092|stomachnull|Stomach structure|Anatomy|false|false|C0872393;C0577027;C0038354;C0496905;C0153943;C0154060|stomach
null|Abdomen>Stomach|Anatomy|false|false|C0872393;C0577027;C0038354;C0496905;C0153943;C0154060|stomach
null|Stomach|Anatomy|false|false|C0872393;C0577027;C0038354;C0496905;C0153943;C0154060|stomachnull|Intraabdominal Route of Administration|Finding|false|false|C1285092|intra-abdominalnull|Intra-abdominal|Modifier|false|false||intra-abdominalnull|null|Device|false|false||loopsnull|Small|LabModifier|false|false||smallnull|Large Intestine|Anatomy|false|false|C5890938;C1416798|large bowelnull|LARGE1 wt Allele|Finding|false|false|C0021853;C0021851|large
null|LARGE1 gene|Finding|false|false|C0021853;C0021851|largenull|Large|LabModifier|false|false||largenull|Intestines|Anatomy|false|false|C5890938;C1416798|bowelnull|null|Modifier|false|false||unremarkablenull|Mesentery|Anatomy|false|false||mesentericnull|Lymphadenopathy|Disorder|false|false||lymphadenopathynull|Swollen Lymph Node|Finding|false|false||lymphadenopathynull|effusion|Finding|true|false||free fluidnull|Free of (attribute)|Finding|true|false||freenull|Empty (qualifier)|Modifier|false|false||freenull|fluid - substance|Drug|true|false||fluid
null|Liquid substance|Drug|true|false||fluidnull|Fluid Specimen Code|Finding|true|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Free of (attribute)|Finding|true|false||freenull|Empty (qualifier)|Modifier|false|false||freenull|Air (substance)|Drug|true|false||air
null|air|Drug|true|false||air
null|air|Drug|true|false||airnull|ACUTE INSULIN RESPONSE|Finding|true|false||air
null|AIRN gene|Finding|true|false||air
null|AI/RHEUM|Finding|true|false||airnull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|abdomennull|Abdomen problem|Finding|false|false|C0230168;C0000726|abdomennull|Abdomen|Anatomy|false|false|C0153662;C0941288|abdomen
null|Abdominal Cavity|Anatomy|false|false|C0153662;C0941288|abdomennull|Stat (do immediately)|Time|false|false||Immediatelynull|Adjacent|Modifier|false|false||adjacent tonull|Adjacent|Modifier|false|false||adjacentnull|To the left (qualifier value)|Modifier|false|false||to the leftnull|Structure of left common iliac artery|Anatomy|false|false|C1552822;C3245511;C1522138|left common iliac arterynull|Table Cell Horizontal Align - left|Finding|false|false|C1261084;C0226363;C0020887|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Common iliac artery structure|Anatomy|false|false|C1552822;C3245511;C1522138|common iliac arterynull|Common Specifications in HL7 V3 Publishing|Finding|false|false|C0020887;C0226363;C1261084|common
null|shared attribute|Finding|false|false|C0020887;C0226363;C1261084|commonnull|Common (qualifier value)|LabModifier|false|false||commonnull|Structure of iliac artery|Anatomy|false|false|C3245511;C1522138;C1552822|iliac arterynull|Bone structure of ilium|Anatomy|false|false||iliacnull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Linear|Modifier|false|false||linearnull|Has focus|Finding|false|false||focusnull|Focal|Modifier|false|false||focusnull|Hyperactive behavior|Disorder|false|false||hypernull|Materials|Drug|false|false||materialnull|patient appearance regarding mental status exam|Procedure|false|false|C0502420|appearancenull|null|Attribute|false|false||appearancenull|Personal appearance|Subject|false|false||appearancenull|Appearance|Modifier|false|false||appearancenull|Kind of quantity - Appearance|LabModifier|false|false||appearancenull|Suture Device|Device|false|false||suture material
null|Surgical sutures|Device|false|false||suture materialnull|Suture Dosage Form|Drug|false|false|C0502420|suturenull|null|Finding|false|false|C0502420|suturenull|Closure by suture|Procedure|false|false|C0502420|suturenull|Suture Joint|Anatomy|false|false|C0009068;C1546803;C2051406;C1706068|suturenull|Suture Device|Device|false|false||suture
null|Surgical sutures|Device|false|false||suturenull|Materials|Drug|false|false||materialnull|null|Finding|false|false||unchangednull|About The Same|Modifier|false|false||unchangednull|null|Time|false|false||priornull|Physical Examination|Procedure|false|false||examination
null|Medical Examination|Procedure|false|false||examinationnull|Examination|Event|false|false||examinationnull|Malignant neoplasm of pelvis|Disorder|true|false|C4266535;C0030797;C0559769|pelvisnull|Pelvis problem|Finding|true|false|C4266535;C0030797;C0559769|pelvisnull|Pelvis+|Anatomy|false|false|C0009068;C0153663;C0812455|pelvis
null|Pelvic cavity structure|Anatomy|false|false|C0009068;C0153663;C0812455|pelvis
null|Pelvis|Anatomy|false|false|C0009068;C0153663;C0812455|pelvisnull|Suture Device|Device|false|false||suture material
null|Surgical sutures|Device|false|false||suture materialnull|Suture Dosage Form|Drug|false|false|C0502420|suturenull|null|Finding|false|false|C0227391;C0502420|suturenull|Closure by suture|Procedure|false|false|C4266535;C0030797;C0559769;C0227391;C0502420|suturenull|Suture Joint|Anatomy|false|false|C1706068;C0009068;C1546803|suturenull|Suture Device|Device|false|false||suture
null|Surgical sutures|Device|false|false||suturenull|Materials|Drug|false|false|C0227391|materialnull|Distal Resection Margin|Attribute|false|false||distalnull|Distal (qualifier value)|Modifier|false|false||distalnull|Sigmoid colon|Anatomy|false|false|C0009068;C0520510;C1546803|sigmoidnull|Carcinoma in situ of colon|Disorder|false|false|C0009368;C4071907|colon
null|Neoplasm of uncertain or unknown behavior of colon|Disorder|false|false|C0009368;C4071907|colon
null|Colonic Diseases|Disorder|false|false|C0009368;C4071907|colonnull|COLON PROBLEM|Finding|false|false|C0009368;C4071907|colonnull|Colon structure (body structure)|Anatomy|false|false|C0750873;C2051406;C0154061;C0009373;C0496907;C0442739|colon
null|Abdomen+Pelvis>Colon|Anatomy|false|false|C0750873;C2051406;C0154061;C0009373;C0496907;C0442739|colonnull|TUBE,COLON,22FR,RADIOPAQUE RUBBER B#7370|Device|false|false||colonnull|Colon <Coloninae>|Entity|false|false||colonnull|null|Finding|false|false|C0009368;C4071907|unchangednull|About The Same|Modifier|false|false||unchangednull|patient appearance regarding mental status exam|Procedure|false|false|C0009368;C4071907|appearancenull|null|Attribute|false|false||appearancenull|Personal appearance|Subject|false|false||appearancenull|Appearance|Modifier|false|false||appearancenull|Kind of quantity - Appearance|LabModifier|false|false||appearancenull|null|Time|false|false||priornull|Physical Examination|Procedure|false|false||examination
null|Medical Examination|Procedure|false|false||examinationnull|Examination|Event|false|false||examinationnull|Consistent with|Finding|false|false|C0500470|consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|Large intestine anastomosis|Procedure|false|false|C0009368;C0500470|colonic anastomosisnull|Colon structure (body structure)|Anatomy|false|false|C0852681;C0332853;C0677554|colonicnull|Anastomosis|Disorder|false|false|C0009368;C0500470|anastomosisnull|null|Procedure|false|false|C0009368;C0500470|anastomosisnull|Anatomical anastomosis|Anatomy|false|false|C0332853;C0677554;C0852681;C0332290|anastomosisnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Stenosis|Finding|false|false|C1515974|stricturenull|Stenosis Morphology|Modifier|false|false||stricturenull|Obstruction|Finding|true|false|C1515974|obstructionnull|null|Finding|false|false|C1515974|sitenull|Anatomic Site|Anatomy|false|false|C1546778;C0028778;C1261287|sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Local Remote Control State - Local|Finding|true|false||localnull|Local|Modifier|false|false||localnull|fluid - substance|Drug|true|false||fluid
null|Liquid substance|Drug|true|false||fluidnull|Fluid Specimen Code|Finding|true|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Collection Object - UML Entity|Finding|false|false||collection
null|Item Collection|Finding|false|false||collection
null|Collections (publication)|Finding|false|false||collection
null|Collection (action)|Finding|false|false||collectionnull|Abscess|Disorder|false|false||abscessnull|null|Finding|false|false||abscessnull|Aspects of signs|Finding|true|false||signs
null|Physical findings|Finding|true|false||signsnull|Manufactured sign|Device|true|false||signsnull|Inflammation|Finding|false|false||inflammationnull|Pelvic cavity structure|Anatomy|false|false||intrapelvicnull|Intrapelvic|Modifier|false|false||intrapelvicnull|null|Device|false|false||loopsnull|Small|LabModifier|false|false||smallnull|Large Intestine|Anatomy|false|false|C5890938;C1416798|large bowelnull|LARGE1 wt Allele|Finding|false|false|C0021851|large
null|LARGE1 gene|Finding|false|false|C0021851|largenull|Large|LabModifier|false|false||largenull|Intestines|Anatomy|false|false||bowelnull|null|Modifier|false|false||unremarkablenull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false||air
null|AIRN gene|Finding|false|false||air
null|AI/RHEUM|Finding|false|false||airnull|Feces|Finding|false|false||stoolnull|Stool seat|Device|false|false||stoolnull|Patterns|Modifier|false|false||patternnull|Intestines|Anatomy|false|false|C0700124;C0012359;C1322279|bowelnull|Pathological Dilatation|Finding|true|false|C0021853|dilatation
null|Dilated|Finding|true|false|C0021853|dilatationnull|Dilate procedure|Procedure|true|false|C0021853|dilatationnull|Neoplasm of uncertain or unknown behavior of appendix|Disorder|false|false|C4037994;C0003617|appendix
null|Benign neoplasm of appendix|Disorder|false|false|C4037994;C0003617|appendix
null|Malignant neoplasm of appendix|Disorder|false|false|C4037994;C0003617|appendixnull|appendix - HTML link|Finding|false|false|C4037994;C0003617|appendixnull|Procedure on appendix|Procedure|false|false|C4037994;C0003617|appendixnull|Abdomen+Pelvis>Appendix|Anatomy|false|false|C0869813;C0348899;C0496779;C0496860;C1552860|appendix
null|Appendix|Anatomy|false|false|C0869813;C0348899;C0496779;C0496860;C1552860|appendixnull|Abdomen+Pelvis>Urinary bladder|Anatomy|false|false|C0872388;C0042131;C0496919;C0496930;C0154017;C0154091;C0869889|urinary bladder
null|Urinary Bladder|Anatomy|false|false|C0872388;C0042131;C0496919;C0496930;C0154017;C0154091;C0869889|urinary bladdernull|Urinary tract|Anatomy|false|false|C0872388;C0496930;C0154017;C0154091|urinarynull|urinary|Modifier|false|false||urinarynull|Neoplasm of uncertain or unknown behavior of bladder|Disorder|false|false|C0042027;C0005682;C0005682;C4037992|bladder
null|Benign neoplasm of bladder|Disorder|false|false|C0042027;C0005682;C0005682;C4037992|bladder
null|Carcinoma in situ of bladder|Disorder|false|false|C0042027;C0005682;C0005682;C4037992|bladdernull|Procedures on bladder|Procedure|false|false|C0005682;C4037992;C0042027;C0005682|bladdernull|Urinary Bladder|Anatomy|false|false|C0869889;C0042131;C0496919;C0496930;C0154017;C0154091;C0872388|bladdernull|Neoplasm of uncertain or unknown behavior of uterus|Disorder|false|false|C0005682;C4037992;C0005682;C4266525;C0042149;C1519876|uterus
null|Uterine Diseases|Disorder|false|false|C0005682;C4037992;C0005682;C4266525;C0042149;C1519876|uterusnull|examination of uterus|Procedure|false|false|C0005682;C4266525;C0042149;C1519876;C0005682;C4037992|uterusnull|Pelvis>Uterus|Anatomy|false|false|C0042131;C0496919;C0869889|uterus
null|Mouse Uterus|Anatomy|false|false|C0042131;C0496919;C0869889|uterus
null|Uterus|Anatomy|false|false|C0042131;C0496919;C0869889|uterusnull|Ocular adnexa structure|Anatomy|false|false||adnexa
null|Adnexa|Anatomy|false|false||adnexa
null|Uterine adnexae structure|Anatomy|false|false||adnexanull|null|Modifier|false|false||unremarkablenull|Lymphadenopathy|Disorder|true|false|C0024204|enlarged lymph nodesnull|Swollen Lymph Node|Finding|true|false|C0024204|enlarged lymph nodesnull|Enlargement procedure|Procedure|false|false|C0024204|enlargednull|Enlarged|Modifier|false|false||enlargednull|benign neoplasm of lymph nodes|Disorder|true|false|C0024204|lymph nodesnull|lymph nodes|Anatomy|false|false|C1293134;C0154054;C4282165;C0024202;C0497156|lymph nodesnull|Lymph|Finding|false|false|C0024204|lymphnull|Malignant neoplasm of pelvis|Disorder|false|false|C4266535;C0030797;C0559769|pelvisnull|Pelvis problem|Finding|false|false|C4266535;C0030797;C0559769|pelvisnull|Pelvis+|Anatomy|false|false|C0153663;C0812455|pelvis
null|Pelvic cavity structure|Anatomy|false|false|C0153663;C0812455|pelvis
null|Pelvis|Anatomy|false|false|C0153663;C0812455|pelvisnull|Platelet Glycoprotein 4, human|Drug|false|false|C0001527|fat
null|FAT1 protein, human|Drug|false|false|C0001527|fat
null|FAT1 protein, human|Drug|false|false|C0001527|fat
null|Fatty acid glycerol esters|Drug|false|false|C0001527|fat
null|Fatty acid glycerol esters|Drug|false|false|C0001527|fatnull|Platelet Glycoprotein 4, human|Finding|false|false|C0001527|fat
null|CD36 gene|Finding|false|false|C0001527|fat
null|FAT1 gene|Finding|false|false|C0001527|fat
null|CD36 wt Allele|Finding|false|false|C0001527|fat
null|FAT1 wt Allele|Finding|false|false|C0001527|fatnull|doxorubicin/fluorouracil/triazinate protocol|Procedure|false|false|C0001527|fatnull|Adipose tissue|Anatomy|false|false|C1435181;C0015677;C3887682;C0279453;C3887682;C0812278;C1705088;C1708004;C1366645;C0262537;C0019294;C0019270|fatnull|Obese build|Subject|false|false||fatnull|Fantse Language|Entity|false|false||fatnull|Left inguinal hernia|Disorder|false|false|C0001527;C0018246|left inguinal hernianull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Hernia, Inguinal|Disorder|false|false|C0001527;C0018246|inguinal hernianull|Inguinal region|Anatomy|false|false|C0019270;C0262537;C0019294|inguinalnull|Hernia|Disorder|false|false|C0018246;C0001527|hernianull|null|Finding|false|false||unchangednull|About The Same|Modifier|false|false||unchangednull|Physical Examination|Procedure|false|false|C0040300;C0225317|Examination
null|Medical Examination|Procedure|false|false|C0040300;C0225317|Examinationnull|Examination|Event|false|false|C0225317;C0040300|Examinationnull|soft tissue|Anatomy|false|false|C4321457;C3542022;C0582103;C0031809;C1522438|soft tissuesnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false|C0225317;C0040300|softnull|Soft|Modifier|false|false||softnull|Body tissue|Anatomy|false|false|C0582103;C0031809;C3542022;C4321457|tissuesnull|Subcutaneous Route of Administration|Finding|false|false|C0225317|subcutaneousnull|subcutaneous|Modifier|false|false||subcutaneousnull|Air (substance)|Drug|false|false|C0040300;C0225317|air
null|air|Drug|false|false|C0040300;C0225317|air
null|air|Drug|false|false|C0040300;C0225317|airnull|ACUTE INSULIN RESPONSE|Finding|false|false|C0225317;C0040300;C1548802|air
null|AIRN gene|Finding|false|false|C0225317;C0040300;C1548802|air
null|AI/RHEUM|Finding|false|false|C0225317;C0040300;C1548802|airnull|soft tissue|Anatomy|false|false|C2681903;C1140091;C1866503;C3542022;C0001861;C3536832|soft tissuesnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false|C1660780;C0040300;C0225317|softnull|Soft|Modifier|false|false||softnull|Body tissue|Anatomy|false|false|C3542022;C2681903;C1140091;C1866503;C0001861;C3536832|tissuesnull|midline cell component|Anatomy|false|false|C3542022|midlinenull|Midline (qualifier value)|Modifier|false|false||midlinenull|Lower anterior|Modifier|false|false||lower anteriornull|Body Site Modifier - Lower|Anatomy|false|false|C2003888;C2681903;C1140091;C1866503|lowernull|Lower (action)|Event|false|false|C1548802|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Adenohypophyseal Diseases|Disorder|false|false||anteriornull|Anterior|Modifier|false|false||anteriornull|Abdominal wall structure|Anatomy|false|false||abdominal wallnull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Walls of a building|Device|false|false||wallnull|Slightly (qualifier value)|Modifier|false|false||slightly
null|Slight (qualifier value)|Modifier|false|false||slightlynull|Greater|LabModifier|false|false||larger
null|Large|LabModifier|false|false||largernull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|null|Time|false|false||priornull|Physical Examination|Procedure|false|false||examination
null|Medical Examination|Procedure|false|false||examinationnull|Examination|Event|false|false||examinationnull|Approximate|Modifier|false|false||approximatelynull|2 Weeks|Time|false|false||2 weeksnull|week|Time|false|false||weeksnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|Small|LabModifier|false|false||smallnull|Has focus|Finding|false|false||focusnull|Focal|Modifier|false|false||focusnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Materials|Drug|false|false||materialnull|Abdominal wall structure|Anatomy|false|false||abdominal wallnull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Walls of a building|Device|false|false||wallnull|Set of muscles|Anatomy|false|false|C1522438|musculaturenull|Subcutaneous Tissue|Anatomy|false|false|C1522438|subcutaneous tissuesnull|Subcutaneous Route of Administration|Finding|false|false|C1995013;C0040300;C0278403|subcutaneousnull|subcutaneous|Modifier|false|false||subcutaneousnull|Body tissue|Anatomy|false|false|C1522438|tissuesnull|External route|Finding|false|false|C1548801|externalnull|Body Site Modifier - External|Anatomy|false|false|C1550509;C0424290;C1516698;C0521134|externalnull|Code System Type - External|Modifier|false|false||external
null|External|Modifier|false|false||externalnull|Compulsive hoarding|Disorder|false|false|C1548801|collectingnull|Collection (action)|Finding|false|false|C1548801|collectingnull|Participation Type - device|Finding|false|false|C1548801|devicenull|Medical Devices|Device|false|false||device
null|Devices|Device|false|false||devicenull|Kind of quantity - Device|LabModifier|false|false||devicenull|Separate|Modifier|false|false||discretenull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Collection Object - UML Entity|Finding|false|false||collection
null|Item Collection|Finding|false|false||collection
null|Collections (publication)|Finding|false|false||collection
null|Collection (action)|Finding|false|false||collectionnull|Abscess formation|Finding|false|false||abscess formationnull|Abscess|Disorder|false|false||abscessnull|null|Finding|false|false||abscessnull|Formation|Finding|false|false||formationnull|Anabolism|Phenomenon|false|false||formationnull|Formations|Modifier|false|false||formationnull|Amenable|Modifier|false|false||amenablenull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|patient appearance regarding mental status exam|Procedure|false|false||appearancenull|null|Attribute|false|false||appearancenull|Personal appearance|Subject|false|false||appearancenull|Appearance|Modifier|false|false||appearancenull|Kind of quantity - Appearance|LabModifier|false|false||appearancenull|Continuous|Finding|false|false||continuednull|Cellulitis|Disorder|false|false||cellulitisnull|cellulitis on exam (physical finding)|Finding|false|false||cellulitisnull|Physical Examination|Procedure|false|false|C4520924;C0262950|Examination
null|Medical Examination|Procedure|false|false|C4520924;C0262950|Examinationnull|Examination|Event|false|false|C4520924;C0262950|Examinationnull|Bone Tissue, Human|Anatomy|false|false|C4321457;C0582103;C0031809|osseous
null|Skeletal bone|Anatomy|false|false|C4321457;C0582103;C0031809|osseousnull|Structure|Modifier|false|false||structuresnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|biologic degeneration|Finding|false|false||degenerative
null|Abnormal degeneration|Finding|false|false||degenerativenull|Disease|Disorder|false|false||diseasenull|null|Modifier|false|false||unremarkablenull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Patient Condition Code - Stable|Finding|false|false||Stablenull|Stable status|Modifier|false|false||Stablenull|patient appearance regarding mental status exam|Procedure|false|false|C0227391;C0227391|appearancenull|null|Attribute|false|false||appearancenull|Personal appearance|Subject|false|false||appearancenull|Appearance|Modifier|false|false||appearancenull|Kind of quantity - Appearance|LabModifier|false|false||appearancenull|Malignant neoplasm of sigmoid colon|Disorder|false|false|C0009368;C4071907;C0500470;C0227391;C0227391|sigmoid colon
null|Benign neoplasm of sigmoid colon|Disorder|false|false|C0009368;C4071907;C0500470;C0227391;C0227391|sigmoid colonnull|Sigmoid colon|Anatomy|false|false|C0852681;C0009373;C0154061;C0496907;C0496864;C0153436;C2051406;C0750873;C0332853|sigmoid colonnull|Sigmoid colon|Anatomy|false|false|C0332853;C0852681;C0009373;C0154061;C0496907;C2051406;C0750873;C0496864;C0153436|sigmoidnull|Large intestine anastomosis|Procedure|false|false|C0009368;C4071907;C0227391;C0227391;C0500470|colon anastomosisnull|Neoplasm of uncertain or unknown behavior of colon|Disorder|false|false|C0227391;C0227391;C0500470;C0009368;C4071907|colon
null|Colonic Diseases|Disorder|false|false|C0227391;C0227391;C0500470;C0009368;C4071907|colon
null|Carcinoma in situ of colon|Disorder|false|false|C0227391;C0227391;C0500470;C0009368;C4071907|colonnull|COLON PROBLEM|Finding|false|false|C0500470;C0227391;C0009368;C4071907;C0227391|colonnull|Colon structure (body structure)|Anatomy|false|false|C0852681;C0496864;C0153436;C0750873;C0332853;C0009373;C0154061;C0496907|colon
null|Abdomen+Pelvis>Colon|Anatomy|false|false|C0852681;C0496864;C0153436;C0750873;C0332853;C0009373;C0154061;C0496907|colonnull|TUBE,COLON,22FR,RADIOPAQUE RUBBER B#7370|Device|false|false||colonnull|Colon <Coloninae>|Entity|false|false||colonnull|Anastomosis|Disorder|false|false|C0227391;C0500470;C0009368;C4071907;C0227391|anastomosisnull|null|Procedure|false|false|C0500470|anastomosisnull|Anatomical anastomosis|Anatomy|false|false|C0750873;C0496864;C0153436;C0852681;C0332853;C0009373;C0154061;C0496907;C0677554|anastomosisnull|Obstruction|Finding|false|false||obstructionnull|Abscess formation|Finding|false|false||abscess formationnull|Abscess|Disorder|false|false||abscessnull|null|Finding|false|false||abscessnull|Formation|Finding|false|false||formationnull|Anabolism|Phenomenon|false|false||formationnull|Formations|Modifier|false|false||formationnull|Subcutaneous air|Finding|false|false|C0836916|subcutaneous airnull|Subcutaneous Route of Administration|Finding|false|false||subcutaneousnull|subcutaneous|Modifier|false|false||subcutaneousnull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false|C0000726;C0836916|air
null|AIRN gene|Finding|false|false|C0000726;C0836916|air
null|AI/RHEUM|Finding|false|false|C0000726;C0836916|airnull|Body Site Modifier - Lower|Anatomy|false|false|C2003888|lowernull|Lower (action)|Event|false|false|C1548802;C0836916|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Abdominal wall structure|Anatomy|false|false|C3842127;C2003888;C2681903;C1140091;C1866503|abdominal wallnull|Abdomen|Anatomy|false|false|C2681903;C1140091;C1866503|abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Walls of a building|Device|false|false||wallnull|midline cell component|Anatomy|false|false|C0007642|midlinenull|Midline (qualifier value)|Modifier|false|false||midlinenull|Cellulitis|Disorder|false|false|C1660780|cellulitisnull|cellulitis on exam (physical finding)|Finding|false|false||cellulitisnull|Separate|Modifier|false|false||discretenull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Collection Object - UML Entity|Finding|false|false||collection
null|Item Collection|Finding|false|false||collection
null|Collections (publication)|Finding|false|false||collection
null|Collection (action)|Finding|false|false||collectionnull|Study Object|Finding|false|false||studynull|Scientific Study|Procedure|false|false||study
null|Study|Procedure|false|false||study
null|Clinical Research|Procedure|false|false||studynull|Room of building - Study|Device|false|false||studynull|Report (document)|Finding|false|false||reportnull|Reporting|Procedure|false|false||reportnull|null|Attribute|false|false||reportnull|Encounter Special Courtesy - staff|Finding|false|false||staffnull|Staff|Subject|false|false||staffnull|On Staff|Modifier|false|false||staffnull|Procedure Practitioner Identifier Code Type - Radiologist|Finding|false|false||radiologistnull|radiologist|Subject|false|false||radiologistnull|Sunlight|Phenomenon|false|false||SUNnull|The Sun|Entity|false|false||SUN
null|Sundanese language|Entity|false|false||SUNnull|Color of urine|Finding|false|false||URINE  COLORnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|color additive|Drug|false|false||COLOR
null|Coloring Excipient|Drug|false|false||COLORnull|color - solid dosage form|Modifier|false|false||COLOR
null|Color|Modifier|false|false||COLORnull|Color quantity|LabModifier|false|false||COLORnull|Cereal plant straw|Drug|false|false||Strawnull|Straw package type|Device|false|false||Strawnull|Straw Color|Modifier|false|false||Strawnull|Straw (unit of presentation)|LabModifier|false|false||Strawnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Hematuria|Disorder|false|false||URINE  BLOODnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|nitrite ion|Drug|false|false||NITRITE
null|Nitrites|Drug|false|false||NITRITE
null|Nitrites|Drug|false|false||NITRITE
null|Nitrites|Drug|false|false||NITRITE
null|nitrite ion|Drug|false|false||NITRITE
null|nitrite ion|Drug|false|false||NITRITEnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Proteins|Drug|false|false||PROTEIN
null|Proteins|Drug|false|false||PROTEINnull|Protein Info|Finding|false|false||PROTEINnull|Protein measurement|Procedure|false|false||PROTEINnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSEnull|Glucose measurement|Procedure|false|false||GLUCOSEnull|Glucose^1.5H post dose glucagon|Lab|false|false||GLUCOSEnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Ketones|Drug|false|false||KETONEnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|bilirubin preparation|Drug|false|false||BILIRUBIN
null|bilirubin preparation|Drug|false|false||BILIRUBIN
null|Bilirubin|Drug|false|false||BILIRUBIN
null|Bilirubin|Drug|false|false||BILIRUBINnull|Bilirubin, total measurement|Procedure|false|false||BILIRUBIN
null|blood bilirubin level test|Procedure|false|false||BILIRUBINnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSEnull|Glucose measurement|Procedure|false|false||GLUCOSEnull|Glucose^1.5H post dose glucagon|Lab|false|false||GLUCOSEnull|urea|Drug|false|false||UREA
null|urea|Drug|false|false||UREA
null|urea|Drug|false|false||UREAnull|Urea measurement|Procedure|false|false||UREAnull|Sodium supplements|Drug|false|false||SODIUM
null|sodium|Drug|false|false||SODIUM
null|sodium|Drug|false|false||SODIUM
null|Sodium Drug Class|Drug|false|false||SODIUMnull|Sodium metabolic function|Finding|false|false||SODIUMnull|Sodium measurement|Procedure|false|false||SODIUMnull|Potassium Drug Class|Drug|false|false||POTASSIUM
null|Dietary Potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|Potassium supplement|Drug|false|false||POTASSIUM
null|Potassium supplement|Drug|false|false||POTASSIUMnull|Potassium metabolic function|Finding|false|false||POTASSIUMnull|Potassium measurement|Procedure|false|false||POTASSIUMnull|chloride ion|Drug|false|false||CHLORIDE
null|Chlorides|Drug|false|false||CHLORIDEnull|Chloride metabolic function|Finding|false|false||CHLORIDEnull|Chloride measurement|Procedure|false|false||CHLORIDEnull|Total|Modifier|false|false||TOTALnull|carbon dioxide|Drug|false|false||CO2
null|carbon dioxide|Drug|false|false||CO2null|MT-CO2 gene|Finding|false|false||CO2
null|null|Finding|false|false||CO2
null|C2 wt Allele|Finding|false|false||CO2null|blood anion gap (lab test)|Procedure|false|false||ANION GAP
null|Anion gap measurement|Procedure|false|false||ANION GAPnull|Anion Gap|Attribute|false|false||ANION GAPnull|Anion gap result|Lab|false|false||ANION GAPnull|Anions|Drug|false|false||ANIONnull|Ras GTPase-Activating Protein 1, Human|Drug|false|false||GAP
null|Ras GTPase-Activating Protein 1, Human|Drug|false|false||GAP
null|GTPase-Activating Proteins|Drug|false|false||GAP
null|GTPase-Activating Proteins|Drug|false|false||GAPnull|RASA1 wt Allele|Finding|false|false||GAP
null|RASA1 gene|Finding|false|false||GAPnull|Gap (space)|Modifier|false|false||GAPnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGPT - Glutamate pyruvate transaminase|Drug|false|false||SGPT
null|SGPT - Glutamate pyruvate transaminase|Drug|false|false||SGPTnull|GPT gene|Finding|false|false||SGPTnull|Serum Alanine Transaminase Test|Procedure|false|false||SGPTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|ASTnull|Atypical Spitz Nevus|Disorder|false|false|C1185650|ASTnull|SLC17A5 wt Allele|Finding|false|false|C1185650|AST
null|SLC17A5 gene|Finding|false|false|C1185650|AST
null|GOT1 gene|Finding|false|false|C1185650|ASTnull|Asterion|Anatomy|false|false|C4522245;C0004002;C0242192;C1121182;C1415181;C1415181;C1420113;C5960784;C0201899|ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||SGOT
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||SGOTnull|GOT1 gene|Finding|false|false|C1185650|SGOTnull|Aspartate aminotransferase measurement|Procedure|false|false|C1185650|SGOTnull|Alkaline Phosphatase|Drug|false|false||ALK PHOS
null|Alkaline Phosphatase|Drug|false|false||ALK PHOSnull|Alkaline phosphatase measurement|Procedure|false|false||ALK PHOSnull|ALK protein, human|Drug|false|false||ALK
null|ALK protein, human|Drug|false|false||ALKnull|ALK protein, human|Finding|false|false||ALK
null|ALK gene|Finding|false|false||ALK
null|ALK wt Allele|Finding|false|false||ALKnull|Phos <Photinae>|Entity|false|false||PHOSnull|lipase|Drug|false|false||LIPASE
null|lipase|Drug|false|false||LIPASE
null|lipase|Drug|false|false||LIPASEnull|Lipase measurement|Procedure|false|false||LIPASEnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C0014792;C1114281|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||HGB
null|Hemoglobin|Drug|false|false||HGBnull|CYGB gene|Finding|false|false||HGBnull|Hemoglobin concentration|Lab|false|false||HGBnull|Hemopoietic stem cell transplant|Procedure|false|false||HCT
null|Hematocrit Measurement|Procedure|false|false||HCTnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Lymph|Finding|false|false||LYMPHSnull|Monos|Drug|false|false||MONOS
null|Mono-S|Drug|false|false||MONOS
null|Monos|Drug|false|false||MONOSnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||EOS
null|Familial eosinophilia|Disorder|false|false||EOSnull|PRSS33 gene|Finding|false|false||EOS
null|IKZF4 gene|Finding|false|false||EOSnull|Eos <Loriini>|Entity|false|false||EOSnull|Primed lymphocyte test|Procedure|false|false||PLTnull|Count Dosing Unit|LabModifier|false|false||COUNT
null|Count|LabModifier|false|false||COUNTnull|BRIEF Health Literacy Screening Tool|Finding|false|false||Brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||Briefnull|Brief|Time|false|false||Briefnull|Shortened|Modifier|false|false||Briefnull|Hospital course|Finding|false|false||Hospital Coursenull|null|Attribute|false|false||Hospital Coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||Coursenull|Admission activity|Procedure|false|false||Admitted
null|Hospital admission|Procedure|false|false||Admittednull|Early|Time|false|false||earlynull|Morning|Time|false|false||morningnull|NPO - Nothing by mouth|Procedure|false|false||NPOnull|null|Entity|false|false||NPOnull|Ventricular Fibrillation, Paroxysmal Familial, 1|Disorder|false|false|C0016520|IVFnull|SCN5A wt Allele|Finding|false|false|C0016520|IVF
null|SCN5A gene|Finding|false|false|C0016520|IVFnull|Assisted Reproductive Technologies|Procedure|false|false|C0016520|IVF
null|Fertilization in Vitro|Procedure|false|false|C0016520|IVFnull|Structure of interventricular foramen|Anatomy|false|false|C0872104;C0015915;C2751898;C1419864;C4321334;C0035273|IVFnull|Resuscitation (procedure)|Procedure|false|false|C0016520|resuscitationnull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Pelvis|Anatomy|false|false||pelvicnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Sigmoid colon|Anatomy|false|false|C0677554;C0332853|sigmoidnull|Anastomosis|Disorder|false|false|C0500470;C0227391|anastomosisnull|null|Procedure|false|false|C0500470;C0227391|anastomosisnull|Anatomical anastomosis|Anatomy|false|false|C0677554;C0332853|anastomosisnull|fluid - substance|Drug|true|false||fluid
null|Liquid substance|Drug|true|false||fluidnull|Fluid Specimen Code|Finding|true|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Free of (attribute)|Finding|false|false||freenull|Empty (qualifier)|Modifier|false|false||freenull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false||air
null|AIRN gene|Finding|false|false||air
null|AI/RHEUM|Finding|false|false||airnull|Firstly|Modifier|false|false||firstnull|First (number)|LabModifier|false|false||firstnull|Night time|Time|false|false||nightnull|monitoring of urine output for fluid balance|Procedure|false|false||urine outputnull|null|Attribute|false|false||urine output
null|null|Attribute|false|false||urine outputnull|Urine volume finding|LabModifier|false|false||urine outputnull|Portion of urine|Finding|false|false||urine
null|null|Finding|false|false||urine
null|Urine|Finding|false|false||urine
null|In Urine|Finding|false|false||urine
null|Urine specimen|Finding|false|false||urinenull|system output|Finding|false|false||outputnull|Measurement of fluid output|Procedure|false|false||outputnull|Constant - dosing instruction fragment|Finding|false|false||constantnull|Constant (qualifier)|Modifier|false|false||constantnull|Loose|Modifier|false|false||loosenull|Feces|Finding|false|false||stoolsnull|null|Attribute|false|false||stoolsnull|Stool seat|Device|false|false||stoolsnull|Toxin|Drug|false|false||toxin
null|Toxin|Drug|false|false||toxinnull|Toxin (disposition)|Modifier|false|false||toxinnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|HDAC2 protein, human|Drug|false|false||HD2
null|HDAC2 protein, human|Drug|false|false||HD2null|HDAC2 wt Allele|Finding|false|false||HD2null|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|GI CONSULT|Procedure|false|false||GI consultnull|Consultation|Procedure|false|false||consultnull|ActInformationPrivacyReason - service|Finding|false|false||servicenull|Software Service|Device|false|false||servicenull|Services|Event|false|false||servicenull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Relate - vinyl resin|Drug|false|false||relatednull|Role Link Type - related|Finding|false|false||related
null|Related (finding)|Finding|false|false||relatednull|Definitely Related to Intervention|Modifier|false|false||related
null|Relationships|Modifier|false|false||relatednull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Reflux|Finding|false|false||refluxnull|Postoperative Period|Time|false|false||postopnull|Course|Time|false|false||coursenull|Wound Infection|Finding|false|false||wound infectionnull|Traumatic Wound|Disorder|false|false||wound
null|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Recommendation|Finding|false|false||recommendationsnull|Anti-Ulcer Agent|Drug|false|false||antacid
null|Antacids|Drug|false|false||antacidnull|Antacid [PE]|Finding|false|false||antacidnull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Gastroenterologist|Subject|false|false||gastroenterologistnull|Helicobacter pylori|Entity|false|false||H.pylorinull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|null|Time|false|false||Prior tonull|null|Time|false|false||Priornull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Low residue diet|Procedure|false|false||low residue dietnull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Residue|Finding|false|false||residuenull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|escitalopram|Drug|false|false||Escitalopram
null|escitalopram|Drug|false|false||Escitalopramnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|pantoprazole|Drug|false|false||Pantoprazole
null|pantoprazole|Drug|false|false||Pantoprazolenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Delayed Release Dosage Form|Drug|false|false||Delayed Releasenull|Views delayed|Attribute|false|false||Delayednull|Deferred|Time|false|false||Delayednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Delayed Release Dosage Form|Drug|false|false||Delayed Releasenull|Views delayed|Attribute|false|false||Delayednull|Deferred|Time|false|false||Delayednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Every twelve hours|Time|false|false||Q12Hnull|12 hours (qualifier value)|Time|false|false||12 hoursnull|Hour|Time|false|false||hoursnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Delayed Release Dosage Form|Drug|false|false||Delayed Releasenull|Views delayed|Attribute|false|false||Delayednull|Deferred|Time|false|false||Delayednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|refill|Finding|false|false||Refillsnull|ranitidine hydrochloride|Drug|false|false||Ranitidine HCl
null|ranitidine hydrochloride|Drug|false|false||Ranitidine HClnull|ranitidine|Drug|false|false||Ranitidine
null|ranitidine|Drug|false|false||Ranitidinenull|Flinders medical centre-7 marker|Drug|false|false||HCl
null|hydrochloride|Drug|false|false||HCl
null|hydrochloride|Drug|false|false||HClnull|Hairy Cell Leukemia|Disorder|false|false||HClnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Bedtime (qualifier value)|Time|false|false||bedtime
null|Once a day, at bedtime|Time|false|false||bedtimenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|fluticasone|Drug|false|false||Fluticasone
null|fluticasone|Drug|false|false||Fluticasonenull|mcg/actuation|LabModifier|false|false||mcg/Actuationnull|microgram|LabModifier|false|false||mcgnull|Actuation (unit of presentation)|LabModifier|false|false||Actuationnull|SPRAY, SUSPENSION|Drug|false|false||Spray, Suspensionnull|Spray Dosage Form|Drug|false|false||Spraynull|Spray (administration method)|Finding|false|false||Spraynull|Spray (action)|Event|false|false||Spraynull|Spray Dosing Unit|LabModifier|false|false||Spraynull|Suspension substance|Drug|false|false||Suspension
null|Suspensions|Drug|false|false||Suspensionnull|Suspension (action)|Finding|false|false||Suspensionnull|Spray Dosage Form|Drug|false|false||Spraynull|Spray (administration method)|Finding|false|false|C0028429|Spraynull|Spray (action)|Event|false|false|C0028429|Spraynull|Spray Dosing Unit|LabModifier|false|false||Spraynull|Nasal brand of oxymetazoline|Drug|false|false|C0028429|Nasal
null|Nasal brand of oxymetazoline|Drug|false|false|C0028429|Nasal
null|Nasal dosage form|Drug|false|false|C0028429|Nasalnull|Nasal Route of Administration|Finding|false|false|C0028429|Nasal
null|Nasal (intended site)|Finding|false|false|C0028429|Nasalnull|null|Anatomy|false|false|C4520890;C1522019;C2003858;C1272939;C0721966;C4521772|Nasalnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|refill|Finding|false|false||Refillsnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Nausea and vomiting|Finding|false|false||nausea and vomitingnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Vomiting|Finding|false|false||vomitingnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Disease|Disorder|false|false||Conditionnull|Logical Condition|Finding|false|false||Conditionnull|null|Attribute|false|false||Conditionnull|Condition|Modifier|false|false||Conditionnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions