 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|25,29
No|30,32
:|32,33
_|36,37
_|37,38
_|38,39
<EOL>|39,40
<EOL>|41,42
Admission|42,51
Date|52,56
:|56,57
_|59,60
_|60,61
_|61,62
Discharge|76,85
Date|86,90
:|90,91
_|94,95
_|95,96
_|96,97
<EOL>|97,98
<EOL>|99,100
Date|100,104
of|105,107
Birth|108,113
:|113,114
_|116,117
_|117,118
_|118,119
Sex|132,135
:|135,136
F|139,140
<EOL>|140,141
<EOL>|142,143
Service|143,150
:|150,151
MEDICINE|152,160
<EOL>|160,161
<EOL>|162,163
IV|175,177
Dye|178,181
,|181,182
Iodine|183,189
Containing|190,200
Contrast|201,209
Media|210,215
/|216,217
Oxycodone|218,227
/|228,229
<EOL>|230,231
cilostazol|231,241
<EOL>|241,242
<EOL>|243,244
Attending|244,253
:|253,254
_|255,256
_|256,257
_|257,258
.|258,259
<EOL>|259,260
<EOL>|261,262
Pneumonia|279,288
identified|289,299
by|300,302
outpatient|303,313
CXR|314,317
<EOL>|317,318
<EOL>|318,319
<EOL>|320,321
Major|321,326
Surgical|327,335
or|336,338
Invasive|339,347
Procedure|348,357
:|357,358
<EOL>|358,359
None|359,363
<EOL>|363,364
<EOL>|364,365
<EOL>|366,367
_|395,396
_|396,397
_|397,398
PMH|399,402
of|403,405
Asthma|406,412
,|412,413
COPD|414,418
,|418,419
tobacco|420,427
use|428,431
,|431,432
p|434,435
/|435,436
w|436,437
4|438,439
days|440,444
of|445,447
"|448,449
cold|449,453
like|454,458
"|458,459
<EOL>|460,461
symptoms|461,469
.|469,470
Pt|471,473
noted|474,479
that|480,484
she|485,488
has|489,492
a|493,494
chronic|495,502
cough|503,508
at|509,511
baseline|512,520
,|520,521
<EOL>|522,523
worse|523,528
at|529,531
night|532,537
,|537,538
but|539,542
noted|543,548
that|549,553
her|554,557
cough|558,563
was|564,567
now|568,571
productive|572,582
of|583,585
<EOL>|586,587
_|587,588
_|588,589
_|589,590
sputum|591,597
and|598,601
was|602,605
a|606,607
/|607,608
w|608,609
wheezing|610,618
and|619,622
subjective|623,633
fevers|634,640
(|641,642
but|642,645
did|646,649
<EOL>|650,651
not|651,654
take|655,659
her|660,663
temperature|664,675
)|675,676
.|676,677
Pt|678,680
also|681,685
noted|686,691
that|692,696
baseline|697,705
DOE|706,709
<EOL>|710,711
increased|711,720
to|721,723
mild|724,728
shortness|729,738
of|739,741
breath|742,748
at|749,751
rest|752,756
during|757,763
the|764,767
same|768,772
<EOL>|773,774
time|774,778
period|779,785
.|785,786
Pt|787,789
took|790,794
tylenol|795,802
and|803,806
robitussin|807,817
to|818,820
good|821,825
effect|826,832
.|832,833
Pt|834,836
<EOL>|837,838
denied|838,844
any|845,848
CP|849,851
,|851,852
but|853,856
noted|857,862
that|863,867
she|868,871
felt|872,876
her|877,880
heart|881,886
"|887,888
flutter|888,895
"|895,896
<EOL>|897,898
during|898,904
this|905,909
time|910,914
period|915,921
.|921,922
No|923,925
changed|926,933
in|934,936
her|937,940
2|941,942
pillow|943,949
orthopnea|950,959
.|959,960
<EOL>|960,961
<EOL>|961,962
Pt|962,964
did|965,968
not|969,972
have|973,977
any|978,981
recent|982,988
sick|989,993
contacts|994,1002
and|1003,1006
denied|1007,1013
any|1014,1017
<EOL>|1018,1019
association|1019,1030
w|1031,1032
/|1032,1033
headache|1034,1042
,|1042,1043
sore|1044,1048
throat|1049,1055
,|1055,1056
sneezing|1057,1065
,|1065,1066
rhinorrhea|1067,1077
,|1077,1078
<EOL>|1079,1080
nausea|1080,1086
,|1086,1087
vomiting|1088,1096
,|1096,1097
diarrhea|1098,1106
,|1106,1107
abdominal|1108,1117
pain|1118,1122
.|1122,1123
<EOL>|1125,1126
<EOL>|1126,1127
In|1127,1129
ED|1130,1132
VS|1133,1135
were|1136,1140
T97|1141,1144
.8|1144,1146
P78|1147,1150
BP136|1151,1156
/|1156,1157
97|1157,1159
R18|1160,1163
O296|1164,1168
%|1168,1169
NC|1169,1171
.|1171,1172
WBC|1173,1176
was|1177,1180
normal|1181,1187
but|1188,1191
<EOL>|1192,1193
pt|1193,1195
noted|1196,1201
to|1202,1204
have|1205,1209
wheezing|1210,1218
on|1219,1221
exam|1222,1226
,|1226,1227
and|1228,1231
CXR|1232,1235
was|1236,1239
suggestive|1240,1250
of|1251,1253
RML|1254,1257
<EOL>|1258,1259
PNA|1259,1262
so|1263,1265
was|1266,1269
given|1270,1275
125mg|1276,1281
methylprednisone|1282,1298
,|1298,1299
750mg|1300,1305
levaquin|1306,1314
,|1314,1315
and|1316,1319
<EOL>|1320,1321
combo|1321,1326
nebs|1327,1331
(|1332,1333
albuterol|1333,1342
/|1342,1343
ipratropim|1343,1353
)|1353,1354
.|1354,1355
CHEM|1356,1360
/|1360,1361
Coags|1361,1366
/|1366,1367
UA|1367,1369
negative|1370,1378
.|1378,1379
<EOL>|1380,1381
<EOL>|1381,1382
Given|1382,1387
co-morbidities|1388,1402
,|1402,1403
decision|1404,1412
was|1413,1416
made|1417,1421
to|1422,1424
admit|1425,1430
pt|1431,1433
while|1434,1439
<EOL>|1440,1441
initiating|1441,1451
Abx|1452,1455
therapy|1456,1463
.|1463,1464
<EOL>|1465,1466
<EOL>|1466,1467
<EOL>|1468,1469
ASTHMA|1491,1497
/|1497,1498
COPD|1498,1502
/|1502,1503
Tobacco|1503,1510
use|1511,1514
<EOL>|1514,1515
Peripheral|1515,1525
Arterial|1526,1534
disease|1535,1542
s|1543,1544
/|1544,1545
p|1545,1546
recent|1547,1553
common|1554,1560
iliac|1561,1566
stenting|1567,1575
<EOL>|1575,1576
ATRIAL|1576,1582
TACHYCARDIA|1583,1594
<EOL>|1597,1598
ATYPICAL|1598,1606
CHEST|1607,1612
PAIN|1613,1617
<EOL>|1620,1621
CERVICAL|1621,1629
RADICULITIS|1630,1641
<EOL>|1644,1645
CERVICAL|1645,1653
SPONDYLOSIS|1654,1665
<EOL>|1668,1669
CORONARY|1669,1677
ARTERY|1678,1684
DISEASE|1685,1692
<EOL>|1695,1696
HEADACHE|1696,1704
<EOL>|1707,1708
HIP|1708,1711
REPLACEMENT|1712,1723
<EOL>|1726,1727
HYPERLIPIDEMIA|1727,1741
<EOL>|1744,1745
HYPERTENSION|1745,1757
<EOL>|1760,1761
OSTEOARTHRITIS|1761,1775
<EOL>|1778,1779
HERPES|1779,1785
ZOSTER|1786,1792
<EOL>|1795,1796
TOBACCO|1796,1803
ABUSE|1804,1809
<EOL>|1812,1813
ATRIAL|1813,1819
FIBRILLATION|1820,1832
<EOL>|1835,1836
ANXIETY|1836,1843
<EOL>|1847,1848
GASTROINTESTINAL|1848,1864
BLEEDING|1865,1873
<EOL>|1876,1877
OSTEOARTHRITIS|1877,1891
<EOL>|1894,1895
ATHEROSCLEROTIC|1895,1910
CARDIOVASCULAR|1911,1925
DISEASE|1926,1933
<EOL>|1936,1937
PERIPHERAL|1937,1947
VASCULAR|1948,1956
DISEASE|1957,1964
<EOL>|1967,1968
URINARY|1968,1975
TRACT|1976,1981
INFECTION|1982,1991
<EOL>|1994,1995
CATARACT|1995,2003
SURGERY|2004,2011
_|2012,2013
_|2013,2014
_|2014,2015
<EOL>|2016,2017
<EOL>|2017,2018
Surgery|2018,2025
:|2025,2026
<EOL>|2026,2027
BILATERAL|2027,2036
COMMON|2037,2043
ILIAC|2044,2049
ARTERY|2050,2056
STENTING|2057,2065
_|2066,2067
_|2067,2068
_|2068,2069
<EOL>|2070,2071
BUNIONECTOMY|2071,2083
<EOL>|2086,2087
HIP|2087,2090
REPLACEMENT|2091,2102
<EOL>|2105,2106
PRIOR|2106,2111
CESAREAN|2112,2120
SECTION|2121,2128
<EOL>|2131,2132
GANGLION|2132,2140
CYST|2141,2145
<EOL>|2146,2147
<EOL>|2148,2149
:|2163,2164
<EOL>|2164,2165
_|2165,2166
_|2166,2167
_|2167,2168
<EOL>|2168,2169
:|2183,2184
<EOL>|2184,2185
Mother|2185,2191
:|2191,2192
_|2193,2194
_|2194,2195
_|2195,2196
,|2196,2197
HTN|2198,2201
<EOL>|2203,2204
Father|2204,2210
:|2210,2211
_|2212,2213
_|2213,2214
_|2214,2215
CA|2216,2218
<EOL>|2220,2221
Brother|2221,2228
:|2228,2229
CA|2230,2232
?|2232,2233
<EOL>|2235,2236
Brother|2236,2243
:|2243,2244
_|2245,2246
_|2246,2247
_|2247,2248
<EOL>|2249,2250
<EOL>|2250,2251
<EOL>|2252,2253
Physical|2253,2261
_|2262,2263
_|2263,2264
_|2264,2265
:|2265,2266
<EOL>|2266,2267
ADMISSION|2267,2276
PHYSICAL|2277,2285
EXAM|2286,2290
:|2290,2291
<EOL>|2291,2292
=|2292,2293
=|2293,2294
=|2294,2295
=|2295,2296
=|2296,2297
=|2297,2298
=|2298,2299
=|2299,2300
=|2300,2301
=|2301,2302
=|2302,2303
=|2303,2304
=|2304,2305
=|2305,2306
=|2306,2307
=|2307,2308
=|2308,2309
=|2309,2310
=|2310,2311
=|2311,2312
=|2312,2313
=|2313,2314
=|2314,2315
=|2315,2316
=|2316,2317
=|2317,2318
=|2318,2319
=|2319,2320
<EOL>|2320,2321
Tm98|2321,2325
.4|2325,2327
,|2327,2328
BP141|2329,2334
/|2334,2335
82|2335,2337
,|2337,2338
P71|2339,2342
,|2342,2343
R20|2344,2347
,|2347,2348
O297|2349,2353
%|2353,2354
RA|2354,2356
<EOL>|2356,2357
GENERAL|2357,2364
:|2364,2365
AOx3|2366,2370
,|2370,2371
pleasant|2372,2380
affect|2381,2387
,|2387,2388
NAD|2389,2392
<EOL>|2392,2393
HEENT|2393,2398
:|2398,2399
MMM|2400,2403
.|2403,2404
no|2405,2407
LAD|2408,2411
.|2411,2412
no|2413,2415
JVD|2416,2419
<EOL>|2419,2420
HEART|2420,2425
:|2425,2426
RRR|2427,2430
,|2430,2431
S1|2432,2434
/|2434,2435
S2|2435,2437
normal|2438,2444
,|2444,2445
no|2446,2448
murmurs|2449,2456
/|2456,2457
gallops|2457,2464
/|2464,2465
rubs|2465,2469
.|2469,2470
<EOL>|2470,2471
LUNGS|2471,2476
:|2476,2477
Coarse|2478,2484
breath|2485,2491
sounds|2492,2498
b|2499,2500
/|2500,2501
l|2501,2502
with|2503,2507
expiratory|2508,2518
wheezing|2519,2527
<EOL>|2528,2529
diffusely|2529,2538
,|2538,2539
RML|2540,2543
/|2543,2544
RLL|2544,2547
crackles|2548,2556
,|2556,2557
no|2558,2560
incr|2561,2565
WOB|2566,2569
(|2570,2571
no|2571,2573
accessory|2574,2583
muscle|2584,2590
<EOL>|2591,2592
use|2592,2595
)|2595,2596
,|2596,2597
no|2598,2600
resp|2601,2605
distress|2606,2614
<EOL>|2614,2615
ABDOMEN|2615,2622
:|2622,2623
soft|2624,2628
,|2628,2629
nontender|2630,2639
,|2639,2640
nondistended|2641,2653
.|2653,2654
normoactive|2655,2666
BS|2667,2669
<EOL>|2671,2672
EXT|2672,2675
:|2675,2676
Warm|2677,2681
,|2681,2682
dry|2683,2686
,|2686,2687
well|2688,2692
perfused|2693,2701
,|2701,2702
1|2703,2704
+|2704,2705
peripheral|2706,2716
edema|2717,2722
to|2723,2725
mid|2726,2729
calves|2730,2736
<EOL>|2737,2738
b|2738,2739
/|2739,2740
l|2740,2741
<EOL>|2742,2743
SKIN|2743,2747
:|2747,2748
dry|2749,2752
,|2752,2753
warm|2754,2758
,|2758,2759
no|2760,2762
rashes|2763,2769
<EOL>|2769,2770
NEURO|2770,2775
/|2775,2776
PSYCH|2776,2781
:|2781,2782
AOx3|2783,2787
,|2787,2788
fluent|2789,2795
speech|2796,2802
,|2802,2803
MAE|2804,2807
spontaneously|2808,2821
<EOL>|2821,2822
<EOL>|2822,2823
DISCHARGE|2823,2832
PHYSICAL|2833,2841
EXAM|2842,2846
:|2846,2847
<EOL>|2847,2848
=|2848,2849
=|2849,2850
=|2850,2851
=|2851,2852
=|2852,2853
=|2853,2854
=|2854,2855
=|2855,2856
=|2856,2857
=|2857,2858
=|2858,2859
=|2859,2860
=|2860,2861
=|2861,2862
=|2862,2863
=|2863,2864
=|2864,2865
=|2865,2866
=|2866,2867
=|2867,2868
=|2868,2869
=|2869,2870
=|2870,2871
=|2871,2872
=|2872,2873
=|2873,2874
=|2874,2875
=|2875,2876
<EOL>|2876,2877
Tm|2877,2879
:|2879,2880
98.7|2880,2884
,|2884,2885
BP148|2886,2891
-|2891,2892
154|2892,2895
/|2895,2896
76|2896,2898
-|2898,2899
89|2899,2901
,|2901,2902
P72|2903,2906
-|2906,2907
81|2907,2909
,|2909,2910
R20|2911,2914
,|2914,2915
O29|2916,2919
_|2919,2920
_|2920,2921
_|2921,2922
-|2922,2923
99RA|2923,2927
<EOL>|2927,2928
GENERAL|2928,2935
:|2935,2936
AOx3|2937,2941
,|2941,2942
pleasant|2943,2951
affect|2952,2958
,|2958,2959
NAD|2960,2963
<EOL>|2963,2964
HEENT|2964,2969
:|2969,2970
MMM|2971,2974
.|2974,2975
no|2976,2978
LAD|2979,2982
.|2982,2983
no|2984,2986
JVD|2987,2990
<EOL>|2990,2991
HEART|2991,2996
:|2996,2997
RRR|2998,3001
,|3001,3002
S1|3003,3005
/|3005,3006
S2|3006,3008
normal|3009,3015
,|3015,3016
no|3017,3019
murmurs|3020,3027
/|3027,3028
gallops|3028,3035
/|3035,3036
rubs|3036,3040
.|3040,3041
<EOL>|3041,3042
LUNGS|3042,3047
:|3047,3048
Coarse|3049,3055
breath|3056,3062
sounds|3063,3069
b|3070,3071
/|3071,3072
l|3072,3073
with|3074,3078
scant|3079,3084
expiratory|3085,3095
wheeze|3096,3102
,|3102,3103
no|3104,3106
<EOL>|3107,3108
incr|3108,3112
WOB|3113,3116
(|3117,3118
no|3118,3120
accessory|3121,3130
muscle|3131,3137
use|3138,3141
)|3141,3142
,|3142,3143
no|3144,3146
resp|3147,3151
distress|3152,3160
<EOL>|3160,3161
ABDOMEN|3161,3168
:|3168,3169
soft|3170,3174
,|3174,3175
nontender|3176,3185
,|3185,3186
nondistended|3187,3199
.|3199,3200
normoactive|3201,3212
BS|3213,3215
<EOL>|3217,3218
EXT|3218,3221
:|3221,3222
Warm|3223,3227
,|3227,3228
dry|3229,3232
,|3232,3233
well|3234,3238
perfused|3239,3247
,|3247,3248
1|3249,3250
+|3250,3251
peripheral|3252,3262
edema|3263,3268
to|3269,3271
mid|3272,3275
calves|3276,3282
<EOL>|3283,3284
b|3284,3285
/|3285,3286
l|3286,3287
<EOL>|3288,3289
SKIN|3289,3293
:|3293,3294
dry|3295,3298
,|3298,3299
warm|3300,3304
,|3304,3305
no|3306,3308
rashes|3309,3315
<EOL>|3315,3316
NEURO|3316,3321
/|3321,3322
PSYCH|3322,3327
:|3327,3328
AOx3|3329,3333
,|3333,3334
fluent|3335,3341
speech|3342,3348
,|3348,3349
MAE|3350,3353
spontaneously|3354,3367
<EOL>|3367,3368
<EOL>|3368,3369
<EOL>|3370,3371
Pertinent|3371,3380
Results|3381,3388
:|3388,3389
<EOL>|3389,3390
PERTINENT|3390,3399
LABS|3400,3404
:|3404,3405
<EOL>|3405,3406
=|3406,3407
=|3407,3408
=|3408,3409
=|3409,3410
=|3410,3411
=|3411,3412
=|3412,3413
=|3413,3414
=|3414,3415
=|3415,3416
=|3416,3417
=|3417,3418
=|3418,3419
=|3419,3420
=|3420,3421
=|3421,3422
=|3422,3423
=|3423,3424
=|3424,3425
=|3425,3426
=|3426,3427
=|3427,3428
=|3428,3429
=|3429,3430
=|3430,3431
=|3431,3432
<EOL>|3432,3433
_|3433,3434
_|3434,3435
_|3435,3436
05|3437,3439
:|3439,3440
13PM|3440,3444
BLOOD|3445,3450
WBC|3451,3454
-|3454,3455
5.0|3455,3458
RBC|3459,3462
-|3462,3463
4|3463,3464
.|3464,3465
70|3465,3467
Hgb|3468,3471
-|3471,3472
13.8|3472,3476
Hct|3477,3480
-|3480,3481
42.7|3481,3485
MCV|3486,3489
-|3489,3490
91|3490,3492
<EOL>|3493,3494
MCH|3494,3497
-|3497,3498
29.3|3498,3502
MCHC|3503,3507
-|3507,3508
32.3|3508,3512
RDW|3513,3516
-|3516,3517
14.3|3517,3521
Plt|3522,3525
_|3526,3527
_|3527,3528
_|3528,3529
<EOL>|3529,3530
_|3530,3531
_|3531,3532
_|3532,3533
06|3534,3536
:|3536,3537
05AM|3537,3541
BLOOD|3542,3547
WBC|3548,3551
-|3551,3552
9|3552,3553
.|3553,3554
0|3554,3555
#|3555,3556
RBC|3557,3560
-|3560,3561
4.25|3561,3565
Hgb|3566,3569
-|3569,3570
12.6|3570,3574
Hct|3575,3578
-|3578,3579
38.6|3579,3583
<EOL>|3584,3585
MCV|3585,3588
-|3588,3589
91|3589,3591
MCH|3592,3595
-|3595,3596
29.7|3596,3600
MCHC|3601,3605
-|3605,3606
32.7|3606,3610
RDW|3611,3614
-|3614,3615
14.4|3615,3619
Plt|3620,3623
_|3624,3625
_|3625,3626
_|3626,3627
<EOL>|3627,3628
_|3628,3629
_|3629,3630
_|3630,3631
05|3632,3634
:|3634,3635
13PM|3635,3639
BLOOD|3640,3645
Neuts|3646,3651
-|3651,3652
53.9|3652,3656
_|3657,3658
_|3658,3659
_|3659,3660
Monos|3661,3666
-|3666,3667
6.6|3667,3670
Eos|3671,3674
-|3674,3675
0.5|3675,3678
<EOL>|3679,3680
Baso|3680,3684
-|3684,3685
0.8|3685,3688
<EOL>|3688,3689
_|3689,3690
_|3690,3691
_|3691,3692
05|3693,3695
:|3695,3696
13PM|3696,3700
BLOOD|3701,3706
_|3707,3708
_|3708,3709
_|3709,3710
PTT|3711,3714
-|3714,3715
31.7|3715,3719
_|3720,3721
_|3721,3722
_|3722,3723
<EOL>|3723,3724
_|3724,3725
_|3725,3726
_|3726,3727
12|3728,3730
:|3730,3731
39PM|3731,3735
BLOOD|3736,3741
UreaN|3742,3747
-|3747,3748
16|3748,3750
Creat|3751,3756
-|3756,3757
0.8|3757,3760
Na|3761,3763
-|3763,3764
138|3764,3767
K|3768,3769
-|3769,3770
3.5|3770,3773
Cl|3774,3776
-|3776,3777
98|3777,3779
<EOL>|3780,3781
HCO3|3781,3785
-|3785,3786
29|3786,3788
AnGap|3789,3794
-|3794,3795
15|3795,3797
<EOL>|3797,3798
_|3798,3799
_|3799,3800
_|3800,3801
06|3802,3804
:|3804,3805
05AM|3805,3809
BLOOD|3810,3815
Glucose|3816,3823
-|3823,3824
142|3824,3827
*|3827,3828
UreaN|3829,3834
-|3834,3835
15|3835,3837
Creat|3838,3843
-|3843,3844
0.7|3844,3847
Na|3848,3850
-|3850,3851
138|3851,3854
<EOL>|3855,3856
K|3856,3857
-|3857,3858
3.5|3858,3861
Cl|3862,3864
-|3864,3865
100|3865,3868
HCO3|3869,3873
-|3873,3874
29|3874,3876
AnGap|3877,3882
-|3882,3883
13|3883,3885
<EOL>|3885,3886
_|3886,3887
_|3887,3888
_|3888,3889
12|3890,3892
:|3892,3893
39PM|3893,3897
BLOOD|3898,3903
proBNP|3904,3910
-|3910,3911
233|3911,3914
<EOL>|3914,3915
_|3915,3916
_|3916,3917
_|3917,3918
05|3919,3921
:|3921,3922
13PM|3922,3926
BLOOD|3927,3932
Calcium|3933,3940
-|3940,3941
9.9|3941,3944
Phos|3945,3949
-|3949,3950
2|3950,3951
.|3951,3952
5|3952,3953
*|3953,3954
Mg|3955,3957
-|3957,3958
1.8|3958,3961
<EOL>|3961,3962
_|3962,3963
_|3963,3964
_|3964,3965
05|3966,3968
:|3968,3969
35PM|3969,3973
BLOOD|3974,3979
Lactate|3980,3987
-|3987,3988
1.5|3988,3991
<EOL>|3991,3992
<EOL>|3992,3993
PERTINENT|3993,4002
MICRO|4003,4008
:|4008,4009
<EOL>|4009,4010
=|4010,4011
=|4011,4012
=|4012,4013
=|4013,4014
=|4014,4015
=|4015,4016
=|4016,4017
=|4017,4018
=|4018,4019
=|4019,4020
=|4020,4021
=|4021,4022
=|4022,4023
=|4023,4024
=|4024,4025
=|4025,4026
=|4026,4027
=|4027,4028
=|4028,4029
=|4029,4030
=|4030,4031
=|4031,4032
=|4032,4033
=|4033,4034
=|4034,4035
=|4035,4036
<EOL>|4036,4037
Urinalysis|4037,4047
:|4047,4048
<EOL>|4048,4049
_|4049,4050
_|4050,4051
_|4051,4052
05|4053,4055
:|4055,4056
30PM|4056,4060
URINE|4061,4066
Blood|4067,4072
-|4072,4073
NEG|4073,4076
Nitrite|4077,4084
-|4084,4085
NEG|4085,4088
Protein|4089,4096
-|4096,4097
TR|4097,4099
<EOL>|4100,4101
Glucose|4101,4108
-|4108,4109
NEG|4109,4112
Ketone|4113,4119
-|4119,4120
NEG|4120,4123
Bilirub|4124,4131
-|4131,4132
NEG|4132,4135
Urobiln|4136,4143
-|4143,4144
NEG|4144,4147
pH|4148,4150
-|4150,4151
7.0|4151,4154
Leuks|4155,4160
-|4160,4161
NEG|4161,4164
<EOL>|4164,4165
_|4165,4166
_|4166,4167
_|4167,4168
05|4169,4171
:|4171,4172
30PM|4172,4176
URINE|4177,4182
RBC|4183,4186
-|4186,4187
0|4187,4188
WBC|4189,4192
-|4192,4193
<|4193,4194
1|4194,4195
Bacteri|4196,4203
-|4203,4204
NONE|4204,4208
Yeast|4209,4214
-|4214,4215
NONE|4215,4219
<EOL>|4220,4221
Epi|4221,4224
-|4224,4225
1|4225,4226
<EOL>|4226,4227
<EOL>|4227,4228
Blood|4228,4233
Cx|4234,4236
(|4237,4238
_|4238,4239
_|4239,4240
_|4240,4241
)|4241,4242
:|4242,4243
NGTD|4244,4248
(|4249,4250
preliminary|4250,4261
)|4261,4262
<EOL>|4262,4263
<EOL>|4263,4264
PERTINENT|4264,4273
STUDIES|4274,4281
:|4281,4282
<EOL>|4282,4283
=|4283,4284
=|4284,4285
=|4285,4286
=|4286,4287
=|4287,4288
=|4288,4289
=|4289,4290
=|4290,4291
=|4291,4292
=|4292,4293
=|4293,4294
=|4294,4295
=|4295,4296
=|4296,4297
=|4297,4298
=|4298,4299
=|4299,4300
=|4300,4301
=|4301,4302
=|4302,4303
=|4303,4304
=|4304,4305
=|4305,4306
=|4306,4307
=|4307,4308
=|4308,4309
<EOL>|4309,4310
<EOL>|4310,4311
EKG|4311,4314
:|4314,4315
Sinus|4316,4321
rhythm|4322,4328
with|4329,4333
frequent|4334,4342
atrial|4343,4349
premature|4350,4359
beats|4360,4365
.|4365,4366
Left|4367,4371
<EOL>|4372,4373
bundle|4373,4379
-|4379,4380
branch|4380,4386
block|4387,4392
with|4393,4397
extensive|4398,4407
repolarization|4408,4422
abnormalities|4423,4436
.|4436,4437
<EOL>|4438,4439
Compared|4439,4447
to|4448,4450
the|4451,4454
previous|4455,4463
tracing|4464,4471
of|4472,4474
_|4475,4476
_|4476,4477
_|4477,4478
the|4479,4482
rhythm|4483,4489
is|4490,4492
now|4493,4496
<EOL>|4497,4498
sinus|4498,4503
<EOL>|4504,4505
<EOL>|4505,4506
CXR|4506,4509
(|4510,4511
_|4511,4512
_|4512,4513
_|4513,4514
)|4514,4515
:|4515,4516
Right|4517,4522
middle|4523,4529
lobe|4530,4534
opacity|4535,4542
concerning|4543,4553
for|4554,4557
<EOL>|4558,4559
pneumonia|4559,4568
.|4568,4569
<EOL>|4569,4570
<EOL>|4571,4572
<EOL>|4594,4595
=|4618,4619
=|4619,4620
=|4620,4621
=|4621,4622
=|4622,4623
=|4623,4624
=|4624,4625
=|4625,4626
=|4626,4627
=|4627,4628
=|4628,4629
=|4629,4630
=|4630,4631
=|4631,4632
=|4632,4633
=|4633,4634
=|4634,4635
=|4635,4636
=|4636,4637
=|4637,4638
=|4638,4639
=|4639,4640
=|4640,4641
=|4641,4642
=|4642,4643
=|4643,4644
=|4644,4645
<EOL>|4645,4646
_|4646,4647
_|4647,4648
_|4648,4649
PMH|4650,4653
of|4654,4656
Asthma|4657,4663
,|4663,4664
COPD|4665,4669
,|4669,4670
CAD|4671,4674
,|4674,4675
tobacco|4676,4683
use|4684,4687
,|4687,4688
who|4689,4692
presented|4693,4702
w|4703,4704
/|4704,4705
4|4706,4707
<EOL>|4708,4709
days|4709,4713
of|4714,4716
shortness|4717,4726
of|4727,4729
breath|4730,4736
and|4737,4740
productive|4741,4751
cough|4752,4757
_|4758,4759
_|4759,4760
_|4760,4761
sputum|4762,4768
)|4768,4769
,|4769,4770
<EOL>|4771,4772
who|4772,4775
was|4776,4779
found|4780,4785
to|4786,4788
have|4789,4793
RML|4794,4797
opacity|4798,4805
on|4806,4808
CXR|4809,4812
at|4813,4815
outpatient|4816,4826
clinic|4827,4833
so|4834,4836
<EOL>|4837,4838
was|4838,4841
referred|4842,4850
to|4851,4853
the|4854,4857
ED|4858,4860
.|4860,4861
<EOL>|4861,4862
<EOL>|4862,4863
ACTIVE|4863,4869
ISSUES|4870,4876
:|4876,4877
<EOL>|4877,4878
=|4878,4879
=|4879,4880
=|4880,4881
=|4881,4882
=|4882,4883
=|4883,4884
=|4884,4885
=|4885,4886
=|4886,4887
=|4887,4888
=|4888,4889
=|4889,4890
=|4890,4891
=|4891,4892
=|4892,4893
=|4893,4894
=|4894,4895
=|4895,4896
=|4896,4897
=|4897,4898
=|4898,4899
=|4899,4900
=|4900,4901
=|4901,4902
=|4902,4903
=|4903,4904
=|4904,4905
<EOL>|4905,4906
#|4906,4907
Community|4907,4916
Acquired|4917,4925
Pneumonia|4926,4935
<EOL>|4935,4936
Pt|4936,4938
presented|4939,4948
to|4949,4951
outpatient|4952,4962
cardiology|4963,4973
appointment|4974,4985
w|4986,4987
/|4987,4988
4|4989,4990
days|4991,4995
of|4996,4998
<EOL>|4999,5000
shortness|5000,5009
of|5010,5012
breath|5013,5019
and|5020,5023
productive|5024,5034
cough|5035,5040
_|5041,5042
_|5042,5043
_|5043,5044
sputum|5045,5051
)|5051,5052
,|5052,5053
and|5054,5057
was|5058,5061
<EOL>|5062,5063
referred|5063,5071
to|5072,5074
primary|5075,5082
care|5083,5087
clinic|5088,5094
(|5095,5096
Dr|5096,5098
.|5098,5099
_|5100,5101
_|5101,5102
_|5102,5103
.|5103,5104
Dr|5105,5107
_|5108,5109
_|5109,5110
_|5110,5111
<EOL>|5112,5113
_|5113,5114
_|5114,5115
_|5115,5116
a|5117,5118
CXR|5119,5122
which|5123,5128
showed|5129,5135
RML|5136,5139
opacity|5140,5147
on|5148,5150
CXR|5151,5154
.|5154,5155
Given|5156,5161
pt|5162,5164
's|5164,5166
<EOL>|5167,5168
underlying|5168,5178
lung|5179,5183
pathology|5184,5193
(|5194,5195
COPD|5195,5199
_|5200,5201
_|5201,5202
_|5202,5203
longstanding|5204,5216
tobacco|5217,5224
use|5225,5228
)|5228,5229
,|5229,5230
<EOL>|5231,5232
and|5232,5235
multiple|5236,5244
co-morbidities|5245,5259
,|5259,5260
she|5261,5264
was|5265,5268
admitted|5269,5277
briefly|5278,5285
to|5286,5288
<EOL>|5289,5290
initiate|5290,5298
antibiotics|5299,5310
/|5310,5311
steroids|5311,5319
and|5320,5323
ensure|5324,5330
that|5331,5335
she|5336,5339
remained|5340,5348
<EOL>|5349,5350
clinically|5350,5360
stable|5361,5367
.|5367,5368
<EOL>|5368,5369
<EOL>|5369,5370
While|5370,5375
RML|5376,5379
opacification|5380,5393
was|5394,5397
suggestive|5398,5408
of|5409,5411
CAP|5412,5415
,|5415,5416
COPD|5417,5421
flare|5422,5427
was|5428,5431
<EOL>|5432,5433
also|5433,5437
consideration|5438,5451
given|5452,5457
afebrile|5458,5466
status|5467,5473
and|5474,5477
normal|5478,5484
WBC|5485,5488
.|5488,5489
Exam|5490,5494
<EOL>|5495,5496
significant|5496,5507
for|5508,5511
afebrile|5512,5520
status|5521,5527
,|5527,5528
saturation|5529,5539
of|5540,5542
97|5543,5545
%|5545,5546
on|5547,5549
RA|5550,5552
<EOL>|5553,5554
(|5554,5555
baseline|5555,5563
95|5564,5566
%|5566,5567
RA|5568,5570
)|5570,5571
,|5571,5572
and|5573,5576
coarse|5577,5583
breath|5584,5590
sounds|5591,5597
w|5598,5599
/|5599,5600
diffuse|5601,5608
<EOL>|5609,5610
expiratory|5610,5620
wheezing|5621,5629
.|5629,5630
<EOL>|5630,5631
<EOL>|5631,5632
Pt|5632,5634
was|5635,5638
treated|5639,5646
w|5647,5648
/|5648,5649
Levaquin|5650,5658
750mg|5659,5664
daily|5665,5670
(|5671,5672
planned|5672,5679
5d|5680,5682
course|5683,5689
)|5689,5690
,|5690,5691
<EOL>|5692,5693
steroids|5693,5701
(|5702,5703
recieved|5703,5711
125|5712,5715
methylprednisone|5716,5732
then|5733,5737
4d|5738,5740
course|5741,5747
of|5748,5750
PO|5751,5753
<EOL>|5754,5755
prednisone|5755,5765
)|5765,5766
,|5766,5767
and|5768,5771
had|5772,5775
nebulizer|5776,5785
treatments|5786,5796
for|5797,5800
symptom|5801,5808
relief|5809,5815
.|5815,5816
<EOL>|5817,5818
<EOL>|5818,5819
Given|5819,5824
her|5825,5828
clinical|5829,5837
stability|5838,5847
,|5847,5848
she|5849,5852
was|5853,5856
discharged|5857,5867
home|5868,5872
with|5873,5877
an|5878,5880
<EOL>|5881,5882
outpatient|5882,5892
f|5893,5894
/|5894,5895
u|5895,5896
w|5897,5898
/|5898,5899
PCP|5900,5903
(|5904,5905
Dr|5905,5907
.|5907,5908
_|5909,5910
_|5910,5911
_|5911,5912
on|5913,5915
_|5916,5917
_|5917,5918
_|5918,5919
.|5919,5920
Until|5921,5926
then|5927,5931
,|5931,5932
<EOL>|5933,5934
pt|5934,5936
will|5937,5941
need|5942,5946
to|5947,5949
complete|5950,5958
course|5959,5965
of|5966,5968
Antibiotics|5969,5980
and|5981,5984
Steroids|5985,5993
.|5993,5994
Pt|5995,5997
<EOL>|5998,5999
was|5999,6002
instructed|6003,6013
to|6014,6016
continue|6017,6025
her|6026,6029
outpatient|6030,6040
COPD|6041,6045
treatment|6046,6055
regimen|6056,6063
<EOL>|6064,6065
on|6065,6067
discharge|6068,6077
.|6077,6078
<EOL>|6078,6079
<EOL>|6079,6080
CHRONIC|6080,6087
ISSUES|6088,6094
:|6094,6095
<EOL>|6095,6096
=|6096,6097
=|6097,6098
=|6098,6099
=|6099,6100
=|6100,6101
=|6101,6102
=|6102,6103
=|6103,6104
=|6104,6105
=|6105,6106
=|6106,6107
=|6107,6108
=|6108,6109
=|6109,6110
=|6110,6111
=|6111,6112
=|6112,6113
=|6113,6114
=|6114,6115
=|6115,6116
=|6116,6117
=|6117,6118
=|6118,6119
=|6119,6120
=|6120,6121
=|6121,6122
<EOL>|6122,6123
#|6123,6124
Coronary|6124,6132
Artery|6133,6139
Disease|6140,6147
<EOL>|6147,6148
Pt|6148,6150
has|6151,6154
a|6155,6156
known|6157,6162
history|6163,6170
of|6171,6173
CAD|6174,6177
,|6177,6178
but|6179,6182
did|6183,6186
not|6187,6190
have|6191,6195
any|6196,6199
chest|6200,6205
pain|6206,6210
<EOL>|6211,6212
during|6212,6218
this|6219,6223
hospitalization|6224,6239
and|6240,6243
EKG|6244,6247
was|6248,6251
unchanged|6252,6261
from|6262,6266
prior|6267,6272
.|6272,6273
<EOL>|6274,6275
Accordingly|6275,6286
,|6286,6287
she|6288,6291
was|6292,6295
continued|6296,6305
on|6306,6308
home|6309,6313
dosages|6314,6321
of|6322,6324
plavix|6325,6331
,|6331,6332
<EOL>|6333,6334
aspirin|6334,6341
,|6341,6342
isosorbid|6343,6352
mononitrate|6353,6364
and|6365,6368
diltiazem|6369,6378
<EOL>|6378,6379
<EOL>|6379,6380
#|6380,6381
Hypertension|6381,6393
<EOL>|6393,6394
Pt|6394,6396
has|6397,6400
a|6401,6402
known|6403,6408
history|6409,6416
of|6417,6419
hypertension|6420,6432
and|6433,6436
was|6437,6440
continued|6441,6450
on|6451,6453
her|6454,6457
<EOL>|6458,6459
home|6459,6463
dose|6464,6468
hydrochlorothiazide|6469,6488
.|6488,6489
<EOL>|6489,6490
<EOL>|6490,6491
#|6491,6492
Glaucoma|6492,6500
<EOL>|6500,6501
Pt|6501,6503
was|6504,6507
continued|6508,6517
on|6518,6520
latanoprost|6521,6532
drops|6533,6538
before|6539,6545
bed|6546,6549
.|6549,6550
<EOL>|6550,6551
<EOL>|6551,6552
#|6552,6553
Hyperlipidemia|6553,6567
<EOL>|6567,6568
Pt|6568,6570
was|6571,6574
continued|6575,6584
on|6585,6587
home|6588,6592
dose|6593,6597
simvastatin|6598,6609
.|6609,6610
<EOL>|6610,6611
<EOL>|6611,6612
Transitional|6612,6624
Issues|6625,6631
:|6631,6632
<EOL>|6632,6633
=|6633,6634
=|6634,6635
=|6635,6636
=|6636,6637
=|6637,6638
=|6638,6639
=|6639,6640
=|6640,6641
=|6641,6642
=|6642,6643
=|6643,6644
=|6644,6645
=|6645,6646
=|6646,6647
=|6647,6648
=|6648,6649
=|6649,6650
=|6650,6651
=|6651,6652
=|6652,6653
=|6653,6654
<EOL>|6654,6655
1.|6655,6657
Pt|6658,6660
will|6661,6665
need|6666,6670
to|6671,6673
continue|6674,6682
Levaquin|6683,6691
750mg|6692,6697
daily|6698,6703
to|6704,6706
complete|6707,6715
5|6716,6717
<EOL>|6718,6719
day|6719,6722
course|6723,6729
(|6730,6731
Day|6731,6734
1|6735,6736
-|6737,6738
_|6739,6740
_|6740,6741
_|6741,6742
<EOL>|6742,6743
2.|6743,6745
Pt|6746,6748
will|6749,6753
need|6754,6758
to|6759,6761
continue|6762,6770
Prednisone|6771,6781
40mg|6782,6786
daily|6787,6792
to|6793,6795
complete|6796,6804
4|6805,6806
<EOL>|6807,6808
day|6808,6811
course|6812,6818
(|6819,6820
Day|6820,6823
1|6824,6825
-|6826,6827
_|6828,6829
_|6829,6830
_|6830,6831
<EOL>|6831,6832
3.|6832,6834
Pt|6835,6837
will|6838,6842
need|6843,6847
to|6848,6850
f|6851,6852
/|6852,6853
u|6853,6854
w|6855,6856
/|6856,6857
PCP|6858,6861
_|6862,6863
_|6863,6864
_|6864,6865
_|6866,6867
_|6867,6868
_|6868,6869
to|6870,6872
assess|6873,6879
response|6880,6888
to|6889,6891
<EOL>|6892,6893
tx|6893,6895
and|6896,6899
for|6900,6903
general|6904,6911
health|6912,6918
care|6919,6923
maintenance|6924,6935
<EOL>|6935,6936
4.|6936,6938
Pt|6939,6941
will|6942,6946
need|6947,6951
to|6952,6954
use|6955,6958
Nebulizer|6959,6968
treatments|6969,6979
at|6980,6982
home|6983,6987
for|6988,6991
<EOL>|6992,6993
symptomatic|6993,7004
relief|7005,7011
for|7012,7015
the|7016,7019
next|7020,7024
wk|7025,7027
until|7028,7033
pneumonia|7034,7043
clears|7044,7050
<EOL>|7050,7051
<EOL>|7051,7052
Code|7052,7056
Status|7057,7063
:|7063,7064
FULL|7065,7069
(|7070,7071
confirmed|7071,7080
w|7081,7082
/|7082,7083
pt|7084,7086
)|7086,7087
<EOL>|7087,7088
Contact|7088,7095
:|7095,7096
_|7097,7098
_|7098,7099
_|7099,7100
(|7101,7102
husband|7102,7109
_|7110,7111
_|7111,7112
_|7112,7113
,|7113,7114
_|7115,7116
_|7116,7117
_|7117,7118
(|7119,7120
_|7120,7121
_|7121,7122
_|7122,7123
)|7123,7124
<EOL>|7124,7125
<EOL>|7126,7127
Medications|7127,7138
on|7139,7141
Admission|7142,7151
:|7151,7152
<EOL>|7152,7153
The|7153,7156
Preadmission|7157,7169
Medication|7170,7180
list|7181,7185
is|7186,7188
accurate|7189,7197
and|7198,7201
complete|7202,7210
.|7210,7211
<EOL>|7211,7212
1.|7212,7214
Albuterol|7215,7224
0.083|7225,7230
%|7230,7231
Neb|7232,7235
Soln|7236,7240
1|7241,7242
NEB|7243,7246
IH|7247,7249
Q6H|7250,7253
:|7253,7254
PRN|7254,7257
shortness|7258,7267
of|7268,7270
<EOL>|7271,7272
breath|7272,7278
<EOL>|7279,7280
2.|7280,7282
Albuterol|7283,7292
Inhaler|7293,7300
2|7301,7302
PUFF|7303,7307
IH|7308,7310
Q4H|7311,7314
:|7314,7315
PRN|7315,7318
shortness|7319,7328
of|7329,7331
breath|7332,7338
<EOL>|7339,7340
3.|7340,7342
Symbicort|7343,7352
(|7353,7354
budesonide|7354,7364
-|7364,7365
formoterol|7365,7375
)|7375,7376
160|7377,7380
-|7380,7381
4.5|7381,7384
mcg|7385,7388
/|7388,7389
actuation|7389,7398
<EOL>|7399,7400
inhalation|7400,7410
BID|7411,7414
<EOL>|7415,7416
4.|7416,7418
Clopidogrel|7419,7430
75|7431,7433
mg|7434,7436
PO|7437,7439
DAILY|7440,7445
<EOL>|7446,7447
5.|7447,7449
Diltiazem|7450,7459
Extended|7460,7468
-|7468,7469
Release|7469,7476
180|7477,7480
mg|7481,7483
PO|7484,7486
DAILY|7487,7492
<EOL>|7493,7494
6.|7494,7496
Fluticasone|7497,7508
Propionate|7509,7519
NASAL|7520,7525
2|7526,7527
SPRY|7528,7532
NU|7533,7535
DAILY|7536,7541
:|7541,7542
PRN|7542,7545
nasal|7546,7551
<EOL>|7552,7553
congestion|7553,7563
<EOL>|7564,7565
7.|7565,7567
Hydrochlorothiazide|7568,7587
50|7588,7590
mg|7591,7593
PO|7594,7596
DAILY|7597,7602
<EOL>|7603,7604
8.|7604,7606
Isosorbide|7607,7617
Mononitrate|7618,7629
(|7630,7631
Extended|7631,7639
Release|7640,7647
)|7647,7648
240|7649,7652
mg|7653,7655
PO|7656,7658
DAILY|7659,7664
<EOL>|7665,7666
9.|7666,7668
Latanoprost|7669,7680
0.005|7681,7686
%|7686,7687
Ophth|7688,7693
.|7693,7694
Soln.|7695,7700
1|7701,7702
DROP|7703,7707
LEFT|7708,7712
EYE|7713,7716
HS|7717,7719
<EOL>|7720,7721
10.|7721,7724
Simvastatin|7725,7736
20|7737,7739
mg|7740,7742
PO|7743,7745
DAILY|7746,7751
<EOL>|7752,7753
11.|7753,7756
Theophylline|7757,7769
ER|7770,7772
300|7773,7776
mg|7777,7779
PO|7780,7782
BID|7783,7786
<EOL>|7787,7788
12.|7788,7791
Tiotropium|7792,7802
Bromide|7803,7810
1|7811,7812
CAP|7813,7816
IH|7817,7819
DAILY|7820,7825
<EOL>|7826,7827
13.|7827,7830
Acetaminophen|7831,7844
325|7845,7848
mg|7849,7851
PO|7852,7854
Q4H|7855,7858
:|7858,7859
PRN|7859,7862
pain|7863,7867
<EOL>|7868,7869
14.|7869,7872
Aspirin|7873,7880
81|7881,7883
mg|7884,7886
PO|7887,7889
DAILY|7890,7895
<EOL>|7896,7897
15.|7897,7900
Calcarb|7901,7908
600|7909,7912
With|7913,7917
Vitamin|7918,7925
D|7926,7927
(|7928,7929
calcium|7929,7936
carbonate|7937,7946
-|7946,7947
vitamin|7947,7954
D3|7955,7957
)|7957,7958
<EOL>|7959,7960
315|7960,7963
/|7963,7964
200|7964,7967
mg|7968,7970
oral|7971,7975
daily|7976,7981
<EOL>|7982,7983
16.|7983,7986
cod|7987,7990
liver|7991,7996
oil|7997,8000
1,250|8001,8006
-|8006,8007
135|8007,8010
unit|8011,8015
oral|8016,8020
BID|8021,8024
<EOL>|8025,8026
17.|8026,8029
Multivitamins|8030,8043
W|8044,8045
/|8045,8046
minerals|8046,8054
1|8055,8056
TAB|8057,8060
PO|8061,8063
DAILY|8064,8069
<EOL>|8070,8071
<EOL>|8071,8072
<EOL>|8073,8074
Discharge|8074,8083
Medications|8084,8095
:|8095,8096
<EOL>|8096,8097
1.|8097,8099
Acetaminophen|8100,8113
325|8114,8117
mg|8118,8120
PO|8121,8123
Q4H|8124,8127
:|8127,8128
PRN|8128,8131
pain|8132,8136
<EOL>|8137,8138
2.|8138,8140
Albuterol|8141,8150
0.083|8151,8156
%|8156,8157
Neb|8158,8161
Soln|8162,8166
1|8167,8168
NEB|8169,8172
IH|8173,8175
Q6H|8176,8179
:|8179,8180
PRN|8180,8183
shortness|8184,8193
of|8194,8196
<EOL>|8197,8198
breath|8198,8204
<EOL>|8205,8206
3.|8206,8208
Aspirin|8209,8216
81|8217,8219
mg|8220,8222
PO|8223,8225
DAILY|8226,8231
<EOL>|8232,8233
4.|8233,8235
Clopidogrel|8236,8247
75|8248,8250
mg|8251,8253
PO|8254,8256
DAILY|8257,8262
<EOL>|8263,8264
5.|8264,8266
Diltiazem|8267,8276
Extended|8277,8285
-|8285,8286
Release|8286,8293
180|8294,8297
mg|8298,8300
PO|8301,8303
DAILY|8304,8309
<EOL>|8310,8311
6.|8311,8313
Fluticasone|8314,8325
Propionate|8326,8336
NASAL|8337,8342
2|8343,8344
SPRY|8345,8349
NU|8350,8352
DAILY|8353,8358
:|8358,8359
PRN|8359,8362
nasal|8363,8368
<EOL>|8369,8370
congestion|8370,8380
<EOL>|8381,8382
7.|8382,8384
Hydrochlorothiazide|8385,8404
50|8405,8407
mg|8408,8410
PO|8411,8413
DAILY|8414,8419
<EOL>|8420,8421
8.|8421,8423
Isosorbide|8424,8434
Mononitrate|8435,8446
(|8447,8448
Extended|8448,8456
Release|8457,8464
)|8464,8465
240|8466,8469
mg|8470,8472
PO|8473,8475
DAILY|8476,8481
<EOL>|8482,8483
9.|8483,8485
Latanoprost|8486,8497
0.005|8498,8503
%|8503,8504
Ophth|8505,8510
.|8510,8511
Soln.|8512,8517
1|8518,8519
DROP|8520,8524
LEFT|8525,8529
EYE|8530,8533
HS|8534,8536
<EOL>|8537,8538
10.|8538,8541
Multivitamins|8542,8555
W|8556,8557
/|8557,8558
minerals|8558,8566
1|8567,8568
TAB|8569,8572
PO|8573,8575
DAILY|8576,8581
<EOL>|8582,8583
11.|8583,8586
Simvastatin|8587,8598
20|8599,8601
mg|8602,8604
PO|8605,8607
DAILY|8608,8613
<EOL>|8614,8615
12.|8615,8618
Theophylline|8619,8631
ER|8632,8634
300|8635,8638
mg|8639,8641
PO|8642,8644
BID|8645,8648
<EOL>|8649,8650
13.|8650,8653
Tiotropium|8654,8664
Bromide|8665,8672
1|8673,8674
CAP|8675,8678
IH|8679,8681
DAILY|8682,8687
<EOL>|8688,8689
14.|8689,8692
Albuterol|8693,8702
Inhaler|8703,8710
2|8711,8712
PUFF|8713,8717
IH|8718,8720
Q4H|8721,8724
:|8724,8725
PRN|8725,8728
shortness|8729,8738
of|8739,8741
breath|8742,8748
<EOL>|8749,8750
15.|8750,8753
Calcarb|8754,8761
600|8762,8765
With|8766,8770
Vitamin|8771,8778
D|8779,8780
(|8781,8782
calcium|8782,8789
carbonate|8790,8799
-|8799,8800
vitamin|8800,8807
D3|8808,8810
)|8810,8811
<EOL>|8812,8813
315|8813,8816
/|8816,8817
200|8817,8820
mg|8821,8823
oral|8824,8828
daily|8829,8834
<EOL>|8835,8836
16.|8836,8839
cod|8840,8843
liver|8844,8849
oil|8850,8853
1,250|8854,8859
-|8859,8860
135|8860,8863
unit|8864,8868
oral|8869,8873
BID|8874,8877
<EOL>|8878,8879
17.|8879,8882
Symbicort|8883,8892
(|8893,8894
budesonide|8894,8904
-|8904,8905
formoterol|8905,8915
)|8915,8916
160|8917,8920
-|8920,8921
4.5|8921,8924
mcg|8925,8928
/|8928,8929
actuation|8929,8938
<EOL>|8939,8940
INHALATION|8940,8950
BID|8951,8954
<EOL>|8955,8956
18.|8956,8959
Cepastat|8960,8968
(|8969,8970
Phenol|8970,8976
)|8976,8977
Lozenge|8978,8985
2|8986,8987
LOZ|8988,8991
PO|8992,8994
Q2H|8995,8998
:|8998,8999
PRN|8999,9002
sore|9003,9007
throat|9008,9014
<EOL>|9015,9016
RX|9016,9018
*|9019,9020
phenol|9020,9026
[|9027,9028
Cepastat|9028,9036
]|9036,9037
14.5|9038,9042
mg|9043,9045
2|9046,9047
lozenges|9048,9056
every|9057,9062
_|9063,9064
_|9064,9065
_|9065,9066
as|9067,9069
needed|9070,9076
<EOL>|9077,9078
for|9078,9081
sore|9082,9086
throat|9087,9093
Disp|9094,9098
#|9099,9100
*|9100,9101
36|9101,9103
Lozenge|9104,9111
Refills|9112,9119
:|9119,9120
*|9120,9121
0|9121,9122
<EOL>|9122,9123
19|9123,9125
.|9125,9126
Levofloxacin|9127,9139
750|9140,9143
mg|9144,9146
PO|9147,9149
Q24H|9150,9154
Duration|9155,9163
:|9163,9164
2|9165,9166
Days|9167,9171
<EOL>|9172,9173
RX|9173,9175
*|9176,9177
levofloxacin|9177,9189
750|9190,9193
mg|9194,9196
1|9197,9198
tablet|9199,9205
(|9205,9206
s|9206,9207
)|9207,9208
by|9209,9211
mouth|9212,9217
daily|9218,9223
Disp|9224,9228
#|9229,9230
*|9230,9231
2|9231,9232
<EOL>|9233,9234
Tablet|9234,9240
Refills|9241,9248
:|9248,9249
*|9249,9250
0|9250,9251
<EOL>|9251,9252
20|9252,9254
.|9254,9255
PredniSONE|9256,9266
40|9267,9269
mg|9270,9272
PO|9273,9275
DAILY|9276,9281
Duration|9282,9290
:|9290,9291
2|9292,9293
Days|9294,9298
<EOL>|9299,9300
RX|9300,9302
*|9303,9304
prednisone|9304,9314
20|9315,9317
mg|9318,9320
2|9321,9322
tablet|9323,9329
(|9329,9330
s|9330,9331
)|9331,9332
by|9333,9335
mouth|9336,9341
daily|9342,9347
Disp|9348,9352
#|9353,9354
*|9354,9355
4|9355,9356
Tablet|9357,9363
<EOL>|9364,9365
Refills|9365,9372
:|9372,9373
*|9373,9374
0|9374,9375
<EOL>|9375,9376
<EOL>|9376,9377
<EOL>|9378,9379
Discharge|9379,9388
Disposition|9389,9400
:|9400,9401
<EOL>|9401,9402
Home|9402,9406
<EOL>|9406,9407
<EOL>|9408,9409
Discharge|9409,9418
Diagnosis|9419,9428
:|9428,9429
<EOL>|9429,9430
Community|9430,9439
Acquired|9440,9448
Pneumonia|9449,9458
<EOL>|9458,9459
COPD|9459,9463
<EOL>|9463,9464
Asthma|9464,9470
<EOL>|9470,9471
<EOL>|9471,9472
<EOL>|9473,9474
Discharge|9495,9504
Condition|9505,9514
:|9514,9515
Stable|9516,9522
<EOL>|9522,9523
Mental|9523,9529
Status|9530,9536
:|9536,9537
AOx3|9538,9542
(|9543,9544
Baseline|9544,9552
)|9552,9553
<EOL>|9553,9554
Ambulatory|9554,9564
Status|9565,9571
:|9571,9572
Baseline|9573,9581
<EOL>|9581,9582
<EOL>|9582,9583
<EOL>|9584,9585
Ms.|9609,9612
_|9613,9614
_|9614,9615
_|9615,9616
,|9616,9617
<EOL>|9617,9618
<EOL>|9618,9619
It|9619,9621
was|9622,9625
a|9626,9627
pleasure|9628,9636
taking|9637,9643
care|9644,9648
of|9649,9651
you|9652,9655
while|9656,9661
you|9662,9665
were|9666,9670
hospitalized|9671,9683
<EOL>|9684,9685
at|9685,9687
_|9688,9689
_|9689,9690
_|9690,9691
.|9691,9692
As|9693,9695
you|9696,9699
know|9700,9704
,|9704,9705
you|9706,9709
were|9710,9714
<EOL>|9715,9716
admitted|9716,9724
for|9725,9728
initial|9729,9736
treatment|9737,9746
of|9747,9749
pneumonia|9750,9759
,|9759,9760
to|9761,9763
ensure|9764,9770
that|9771,9775
you|9776,9779
<EOL>|9780,9781
were|9781,9785
responding|9786,9796
well|9797,9801
to|9802,9804
the|9805,9808
antibiotics|9809,9820
,|9820,9821
given|9822,9827
your|9828,9832
history|9833,9840
of|9841,9843
<EOL>|9844,9845
COPD|9845,9849
/|9849,9850
Asthma|9850,9856
.|9856,9857
Fortunately|9858,9869
,|9869,9870
you|9871,9874
responded|9875,9884
quite|9885,9890
well|9891,9895
to|9896,9898
the|9899,9902
<EOL>|9903,9904
Antiobiotics|9904,9916
,|9916,9917
Steroids|9918,9926
,|9926,9927
and|9928,9931
Nebulizer|9932,9941
treatments|9942,9952
that|9953,9957
were|9958,9962
<EOL>|9963,9964
administered|9964,9976
.|9976,9977
Since|9978,9983
your|9984,9988
breathing|9989,9998
was|9999,10002
stable|10003,10009
and|10010,10013
you|10014,10017
were|10018,10022
<EOL>|10023,10024
responding|10024,10034
appropriately|10035,10048
to|10049,10051
treatments|10052,10062
,|10062,10063
you|10064,10067
were|10068,10072
discharged|10073,10083
to|10084,10086
<EOL>|10087,10088
home|10088,10092
.|10092,10093
However|10094,10101
,|10101,10102
you|10103,10106
should|10107,10113
be|10114,10116
vigilant|10117,10125
in|10126,10128
making|10129,10135
sure|10136,10140
that|10141,10145
you|10146,10149
<EOL>|10150,10151
continue|10151,10159
the|10160,10163
antibiotics|10164,10175
&|10176,10177
steroids|10178,10186
for|10187,10190
the|10191,10194
short|10195,10200
course|10201,10207
listed|10208,10214
<EOL>|10215,10216
on|10216,10218
the|10219,10222
medication|10223,10233
page|10234,10238
.|10238,10239
You|10240,10243
should|10244,10250
also|10251,10255
be|10256,10258
sure|10259,10263
to|10264,10266
see|10267,10270
Dr.|10271,10274
_|10275,10276
_|10276,10277
_|10277,10278
<EOL>|10279,10280
at|10280,10282
your|10283,10287
next|10288,10292
appointment|10293,10304
to|10305,10307
ensure|10308,10314
that|10315,10319
your|10320,10324
pneumonia|10325,10334
has|10335,10338
<EOL>|10339,10340
resolved|10340,10348
.|10348,10349
<EOL>|10349,10350
<EOL>|10351,10352
Followup|10352,10360
Instructions|10361,10373
:|10373,10374
<EOL>|10374,10375
_|10375,10376
_|10376,10377
_|10377,10378
<EOL>|10378,10379

