CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Known|Modifier|false|false||Knownnull|Hypersensitivity|Finding|true|false||Allergiesnull|null|Attribute|true|false||Allergiesnull|Pharmaceutical Preparations|Drug|false|false||Drugsnull|Drugs - dental services|Procedure|false|false||Drugsnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Chief complaint (finding)|Finding|false|false||Chief Complaintnull|Complaint (finding)|Finding|false|false||Complaintnull|null|Attribute|false|false||Complaintnull|Abdomen distended|Finding|false|false|C0000726|Abdominal distentionnull|Abdomen|Anatomy|false|false|C0424755;C0015967;C0000731;C3714614;C0012359;C1549543;C0030193|Abdominalnull|Abdominal (qualifier value)|Modifier|false|false||Abdominalnull|Distention|Finding|false|false|C0000726|distention
null|Pathological Dilatation|Finding|false|false|C0000726|distentionnull|Pain and Fever|Drug|false|false||pain and fever
null|Pain and Fever|Drug|false|false||pain and fevernull|Administration Method - Pain|Finding|false|false|C0000726|pain
null|Pain|Finding|false|false|C0000726|painnull|null|Attribute|false|false||painnull|Fever symptoms (finding)|Finding|false|false|C0000726|fever
null|Fever|Finding|false|false|C0000726|fevernull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Paracentesis|Procedure|false|false||Paracentesisnull|Diagnostic agents|Drug|false|false||diagnosticnull|Location Service Code - Diagnostic|Finding|false|false||diagnostic
null|Diagnostic|Finding|false|false||diagnosticnull|Diagnostic dental procedure|Procedure|false|false||diagnostic
null|Diagnosis|Procedure|false|false||diagnosticnull|Therapeutic brand of coal tar|Drug|false|false||therapeutic
null|Therapeutic brand of coal tar|Drug|false|false||therapeuticnull|Therapeutic - Location Service Code|Finding|false|false||therapeutic
null|Therapeutic|Finding|false|false||therapeuticnull|Therapeutic procedure|Procedure|false|false||therapeuticnull|History of present illness (finding)|Finding|false|false||History of Present Illnessnull|null|Attribute|false|false||History of Present Illnessnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Present illness|Finding|false|false||Present Illnessnull|Present|Finding|false|false||Present
null|Presentation|Finding|false|false||Presentnull|Illness (finding)|Finding|false|false||Illnessnull|Recent|Time|false|false||recentlynull|Hepatitis, Alcoholic|Disorder|false|false||alcoholic hepatitisnull|Alcoholics|Subject|false|false||alcoholicnull|Hepatitis A|Disorder|false|false||hepatitis
null|Hepatitis|Disorder|false|false||hepatitisnull|Persistent|Time|false|false||persistentnull|Ascites|Disorder|false|false||ascitesnull|Peritoneal Effusion|Finding|false|false||ascitesnull|Persistent|Time|false|false||persistentnull|Fever|Finding|false|false||feversnull|Leukocytosis|Disorder|false|false||leukocytosisnull|Blood leukocyte number above reference range|Finding|false|false||leukocytosisnull|Hepatitis A|Disorder|false|false||hepatitis
null|Hepatitis|Disorder|false|false||hepatitisnull|Patient Outcome - Worsening|Finding|false|false||worseningnull|Worsening (qualifier value)|Modifier|false|false||worseningnull|Abdomen distended|Finding|false|false|C0000726|abdominal distentionnull|Abdomen|Anatomy|false|false|C3714614;C0012359;C0000731|abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Distention|Finding|false|false|C0000726|distention
null|Pathological Dilatation|Finding|false|false|C0000726|distentionnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Persistent fever|Finding|false|false||persistent fevernull|Persistent|Time|false|false||persistentnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Chills|Finding|true|false||chillsnull|Have Sweats|Finding|false|false||have sweatsnull|Sweating|Finding|false|false||sweats
null|Sweat|Finding|false|false||sweatsnull|Night time|Time|false|false||nightnull|null|Time|false|false||prior tonull|null|Time|false|false||priornull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Compliance behavior|Finding|false|false||compliantnull|Compliant (qualifier value)|Modifier|false|false||compliantnull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Fluid restriction|Procedure|false|false||fluid restrictionnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Restricted|Finding|false|false||restrictionnull|Increased (finding)|Finding|false|false||increased
null|Increase|Finding|false|false||increasednull|Increased|LabModifier|false|false||increasednull|fluid - substance|Drug|true|false||fluid
null|Liquid substance|Drug|true|false||fluidnull|Fluid Specimen Code|Finding|true|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Sodium supplements|Drug|true|false||sodium
null|sodium|Drug|true|false||sodium
null|sodium|Drug|true|false||sodium
null|Sodium Drug Class|Drug|true|false||sodiumnull|Sodium metabolic function|Finding|true|false||sodiumnull|Sodium measurement|Procedure|true|false||sodiumnull|Intake|Finding|false|false||intakenull|Measurement of fluid intake|Procedure|false|false||intake
null|Intake (treatment)|Procedure|false|false||intakenull|sobriety|Finding|false|false||sobrietynull|Alcohols|Drug|false|false||alcohol
null|Alcohols|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcoholnull|Alcohol - Recreational Drug Use Code|Finding|false|false||alcoholnull|Fever|Finding|false|false||febrilenull|Tender|Modifier|false|false||tendernull|Palpation|Procedure|false|false||palpationnull|Initial (abbreviation)|Finding|false|false||initialnull|Initially|Time|false|false||initialnull|Firstly|Modifier|false|false||initialnull|Taking vital signs|Procedure|false|false||vital signsnull|null|Attribute|false|false||vital signs
null|Vital signs|Attribute|false|false||vital signsnull|Vital High Nitrogen Enteral Nutrition|Drug|false|false||vitalnull|Vital (qualifier value)|Modifier|false|false||vitalnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|C1orf210 gene|Finding|false|false||tempnull|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Procedure|false|false||tempnull|Temperature|LabModifier|false|false||tempnull|Physiologic pulse|Finding|false|false||pulsenull|Pulse taking|Procedure|false|false||pulsenull|Pulse Rate|Attribute|false|false||pulsenull|Pulse phenomenon|Phenomenon|false|false||pulsenull|Ativan|Drug|false|false||Ativan
null|Ativan|Drug|false|false||Ativannull|morphine|Drug|false|false||morphine
null|morphine|Drug|false|false||morphinenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Tylenol|Drug|false|false||tylenol
null|Tylenol|Drug|false|false||tylenolnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|ondansetron|Drug|false|false||ondansetron
null|ondansetron|Drug|false|false||ondansetronnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Anxiety Disorders|Disorder|false|false||anxiety
null|Anxiety|Disorder|false|false||anxietynull|Anxiety symptoms|Finding|false|false||anxietynull|Diagnostic agents|Drug|false|false||diagnosticnull|Location Service Code - Diagnostic|Finding|false|false||diagnostic
null|Diagnostic|Finding|false|false||diagnosticnull|Diagnostic dental procedure|Procedure|false|false||diagnostic
null|Diagnosis|Procedure|false|false||diagnosticnull|Paracentesis|Procedure|false|false||paracentesisnull|Initially|Time|false|false||initiallynull|ceftriaxone|Drug|false|false||ceftriaxone
null|ceftriaxone|Drug|false|false||ceftriaxonenull|Possible|Finding|false|false||possiblenull|Possible diagnosis|Modifier|false|false||possible
null|Possibly Related to Intervention|Modifier|false|false||possiblenull|Androgen Binding Protein|Drug|false|false||SBP
null|Androgen Binding Protein|Drug|false|false||SBPnull|CCHCR1 wt Allele|Finding|false|false||SBP
null|SHBG wt Allele|Finding|false|false||SBPnull|Systolic blood pressure measurement|Procedure|false|false||SBPnull|Systolic Pressure|Attribute|false|false||SBPnull|Pharmaceutical Preparations|Drug|false|false||Medicinenull|Medicine|Title|false|false||Medicinenull|Further|Modifier|false|false||furthernull|Disease Management|Procedure|false|false||managementnull|Management Occupations|Subject|false|false||managementnull|Management procedure|Event|false|false||management
null|Administration occupational activities|Event|false|false||managementnull|Floor (anatomic)|Anatomy|false|false||floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Floor (anatomic)|Anatomy|false|false|C3889585;C0026516;C5444612|floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Mood (psychological function)|Finding|false|false|C3714591|mood
null|mood (physical finding)|Finding|false|false|C3714591|mood
null|Mood (attribute)|Finding|false|false|C3714591|moodnull|null|Attribute|false|false||moodnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Weepiness|Finding|false|false||tearfulnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Pleasant|Finding|false|false||pleasantnull|Confusion|Disorder|true|false||confusednull|Precaution Code - Confused|Finding|true|false||confused
null|Clouded consciousness|Finding|true|false||confusednull|Cough (guaifenesin)|Drug|true|false||cough
null|Cough (guaifenesin)|Drug|true|false||coughnull|Coughing|Finding|true|false||coughnull|Dysuria|Finding|true|false||dysurianull|rectal discharge diarrhea (physical finding)|Finding|false|false||diarrhea
null|Diarrhea|Finding|false|false||diarrheanull|Eruption of skin (disorder)|Disorder|false|false||rashnull|Skin rash|Finding|false|false||rash
null|Eruptions|Finding|false|false||rash
null|Exanthema|Finding|false|false||rashnull|Decreasing|Finding|false|false||decreased
null|Reduced|Finding|false|false||decreasednull|Decreased|LabModifier|false|false||decreasednull|day|Time|false|false||daysnull|Review of systems (procedure)|Procedure|false|false||Review of Systemsnull|null|Attribute|false|false||Review of Systems
null|null|Attribute|false|false||Review of Systemsnull|Review of|Finding|false|false||Review ofnull|Review (Publication Type)|Finding|false|false||Review
null|Act Class - review|Finding|false|false||Reviewnull|System|Finding|false|false||Systemsnull|Proline dehydrogenase deficiency|Disorder|false|false||HPInull|History of present illness (finding)|Finding|false|false||HPI
null|allene oxide synthase activity|Finding|false|false||HPInull|Chills|Finding|true|false||chillsnull|Headache|Finding|true|false||headachenull|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false|C1305231;C0030471|sinus
null|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false|C1305231;C0030471|sinusnull|pathologic fistula|Disorder|false|false|C1305231;C0030471|sinusnull|Sinus - general anatomical term|Anatomy|false|false|C0684239;C0234233;C0723346;C0016169|sinus
null|Nasal sinus|Anatomy|false|false|C0684239;C0234233;C0723346;C0016169|sinusnull|Emotional tenderness|Finding|false|false|C1305231;C0030471|tenderness
null|Sore to touch|Finding|false|false|C1305231;C0030471|tendernessnull|Rhinorrhea|Finding|false|false||rhinorrheanull|Congestion|Finding|false|false||congestionnull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C2926613;C1549543;C0030193;C0741025;C0008031|chest
null|Anterior thoracic region|Anatomy|false|false|C2926613;C1549543;C0030193;C0741025;C0008031|chestnull|Administration Method - Pain|Finding|false|false|C1527391;C0817096|pain
null|Pain|Finding|false|false|C1527391;C0817096|painnull|null|Attribute|false|false||painnull|Tightness sensation quality|Modifier|false|false||tightnessnull|Palpitations|Finding|false|false||palpitationsnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Dyspnea|Finding|true|false||shortness of breathnull|null|Attribute|true|false||shortness of breathnull|Breath|Finding|false|false||breathnull|Wheezing|Finding|true|false||wheezesnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Vomiting|Finding|false|false||vomitingnull|rectal discharge diarrhea (physical finding)|Finding|false|false||diarrhea
null|Diarrhea|Finding|false|false||diarrheanull|Constipation|Finding|false|false||constipationnull|Recent|Time|false|false||recentnull|Changing|Finding|true|false|C0021853|change innull|Changed status|LabModifier|false|false||change innull|Changing|Finding|true|false|C0021853|changenull|Change - procedure|Procedure|true|false|C0021853|changenull|Delta (difference)|LabModifier|false|false||change
null|Changed status|LabModifier|false|false||changenull|Intestines|Anatomy|false|false|C0392747;C0392747;C4319952|bowelnull|Neoplasm of uncertain or unknown behavior of bladder|Disorder|false|false|C0005682|bladder
null|Benign neoplasm of bladder|Disorder|false|false|C0005682|bladder
null|Carcinoma in situ of bladder|Disorder|false|false|C0005682|bladdernull|Procedures on bladder|Procedure|false|false|C0005682|bladdernull|Urinary Bladder|Anatomy|false|false|C0018464;C2242848;C0496930;C0154017;C0154091;C0872388|bladdernull|Behaviorial Habits|Finding|false|false|C0005682|habits
null|habits (history)|Finding|false|false|C0005682|habitsnull|Dysuria|Finding|true|false||dysurianull|Arthralgia|Finding|true|false||arthralgiasnull|Myalgia|Finding|true|false||myalgiasnull|Skin rash|Finding|true|false||rashes
null|Exanthema|Finding|true|false||rashesnull|Impaired skin integrity|Finding|true|false|C1123023;C4520765|skin breakdown
null|Broken skin|Finding|true|false|C1123023;C4520765|skin breakdownnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765|skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765|skinnull|Skin Specimen Source Code|Finding|false|false|C1123023;C4520765|skin
null|Skin Specimen|Finding|false|false|C1123023;C4520765|skinnull|Skin, Human|Anatomy|false|false|C0699900;C4048181;C0150077;C1265875;C1546781;C0444099;C0178298;C0496955|skin
null|Skin|Anatomy|false|false|C0699900;C4048181;C0150077;C1265875;C1546781;C0444099;C0178298;C0496955|skinnull|Disintegration (morphologic abnormality)|Disorder|false|false|C1123023;C4520765|breakdownnull|Catabolism|Finding|false|false|C1123023;C4520765|breakdownnull|Numbness|Finding|true|false||numbness
null|Hypesthesia|Finding|true|false||numbnessnull|Paresthesia|Disorder|true|false||tinglingnull|Has tingling sensation|Finding|true|false||tinglingnull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|Subject's Feelings|Finding|true|false||feelings
null|Feelings|Finding|true|false||feelingsnull|Cancer patients and suicide and depression|Disorder|true|false||depression
null|Mental Depression|Disorder|true|false||depression
null|Depressive disorder|Disorder|true|false||depression
null|Depressed mood|Disorder|true|false||depressionnull|Depression - motion|Finding|true|false||depression
null|null|Finding|true|false||depressionnull|Depression - recess|Modifier|false|false||depressionnull|Anxiety Disorders|Disorder|false|false||anxiety
null|Anxiety|Disorder|false|false||anxietynull|Anxiety symptoms|Finding|false|false||anxietynull|All other|Finding|false|false||All othernull|Review of systems (procedure)|Procedure|false|false||review of systemsnull|null|Attribute|false|false||review of systems
null|null|Attribute|false|false||review of systemsnull|Review of|Finding|false|false||review ofnull|Review (Publication Type)|Finding|false|false||review
null|Act Class - review|Finding|false|false||reviewnull|System|Finding|false|false||systemsnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Alcohol abuse|Disorder|false|false||Alcohol abusenull|Alcohols|Drug|false|false||Alcohol
null|Alcohols|Drug|false|false||Alcohol
null|ethanol|Drug|false|false||Alcohol
null|ethanol|Drug|false|false||Alcoholnull|Alcohol - Recreational Drug Use Code|Finding|false|false||Alcoholnull|Drug abuse|Disorder|false|false||abusenull|Victim of abuse (finding)|Finding|false|false||abusenull|Abuse|Event|false|false||abusenull|Hepatitis, Alcoholic|Disorder|false|false||Alcoholic hepatitisnull|Alcoholics|Subject|false|false||Alcoholicnull|Hepatitis A|Disorder|false|false||hepatitis
null|Hepatitis|Disorder|false|false||hepatitisnull|Persistent fever|Finding|false|false||persistent fevernull|Persistent|Time|false|false||persistentnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Leukocytosis|Disorder|false|false||leukocytosisnull|Blood leukocyte number above reference range|Finding|false|false||leukocytosisnull|Ascites|Disorder|false|false||Ascitesnull|Peritoneal Effusion|Finding|false|false||Ascitesnull|Chronic back pain|Finding|false|false||Chronic back painnull|Chronic - Admission Level of Care Code|Finding|false|false||Chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||Chronicnull|chronic|Time|false|false||Chronicnull|Back Pain|Finding|false|false||back painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Social and personal history|Finding|false|false||Social History
null|Social History|Finding|false|false||Social Historynull|Social|Finding|false|false||Socialnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Family Medical History|Finding|false|false||Family Historynull|Entity Name Part Type - family|Finding|false|false||Family
null|Last Name|Finding|false|false||Family
null|Living Arrangement - Family|Finding|false|false||Family
null|Family (taxonomic)|Finding|false|false||Family
null|Family Collection|Finding|false|false||Familynull|Family|Subject|false|false||Familynull|History of present illness (finding)|Finding|false|true||History
null|History of previous events|Finding|false|true||History
null|Historical aspects qualifier|Finding|false|true||History
null|Medical History|Finding|false|true||History
null|Concept History|Finding|false|true||Historynull|History|Subject|false|false||Historynull|Relationship - Mother|Finding|false|false||Mothernull|Mother (person)|Subject|false|false||Mothernull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|Family Medical History|Finding|true|false|C4037986;C1278929;C0023884|family history ofnull|Family Medical History|Finding|true|false|C4037986;C1278929;C0023884|family historynull|Entity Name Part Type - family|Finding|false|false||family
null|Last Name|Finding|false|false||family
null|Living Arrangement - Family|Finding|false|false||family
null|Family (taxonomic)|Finding|false|false||family
null|Family Collection|Finding|false|false||familynull|Family|Subject|false|false||familynull|null|Finding|true|true|C4037986;C1278929;C0023884|history of liver diseasenull|Medical History|Finding|true|true|C4037986;C1278929;C0023884|history ofnull|History of present illness (finding)|Finding|true|false|C4037986;C1278929;C0023884|history
null|History of previous events|Finding|true|false|C4037986;C1278929;C0023884|history
null|Historical aspects qualifier|Finding|true|false|C4037986;C1278929;C0023884|history
null|Medical History|Finding|true|false|C4037986;C1278929;C0023884|history
null|Concept History|Finding|true|false|C4037986;C1278929;C0023884|historynull|History|Subject|false|false||historynull|Liver diseases|Disorder|true|true|C4037986;C1278929;C0023884|liver disease
null|Hepatobiliary Disorder|Disorder|true|true|C4037986;C1278929;C0023884|liver diseasenull|Liver brand of Vitamin B 12|Drug|true|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|true|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|true|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|true|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|true|false|C4037986;C1278929;C0023884|livernull|Benign neoplasm of liver|Disorder|true|false|C4037986;C1278929;C0023884|liver
null|Liver diseases|Disorder|true|false|C4037986;C1278929;C0023884|livernull|Liver problem|Finding|true|false|C4037986;C1278929;C0023884|livernull|Procedures on liver|Procedure|true|false|C4037986;C1278929;C0023884|livernull|Abdomen>Liver|Anatomy|false|false|C0721399;C0023899;C0872387;C0012634;C0241889;C0023895;C0496870;C0577060;C0241889;C0262926;C1705255;C0019665;C0262512;C2004062;C0267792;C0023895;C0455550;C0262926|liver
null|null|Anatomy|false|false|C0721399;C0023899;C0872387;C0012634;C0241889;C0023895;C0496870;C0577060;C0241889;C0262926;C1705255;C0019665;C0262512;C2004062;C0267792;C0023895;C0455550;C0262926|liver
null|Liver|Anatomy|false|false|C0721399;C0023899;C0872387;C0012634;C0241889;C0023895;C0496870;C0577060;C0241889;C0262926;C1705255;C0019665;C0262512;C2004062;C0267792;C0023895;C0455550;C0262926|livernull|Disease|Disorder|true|true|C4037986;C1278929;C0023884|diseasenull|Numerous|LabModifier|false|false||Multiplenull|Relative (related person)|Subject|false|false||relativesnull|Alcoholic Intoxication, Chronic|Disorder|false|false||alcoholismnull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GEN
null|GEN1 wt Allele|Finding|false|false||GEN
null|GEN1 gene|Finding|false|false||GENnull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|Labile affect|Disorder|false|false||labile affectnull|Affect (mental function)|Finding|false|false||affectnull|assessment of affect|Procedure|false|false||affectnull|Pleasant|Finding|false|false||pleasantnull|Weepiness|Finding|false|false||tearfulnull|HEENT|Anatomy|false|false||HEENTnull|Lesion|Finding|true|false||lesionsnull|Mild Severity of Illness Code|Finding|false|false|C0036410|mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Scleral icterus|Finding|false|false|C0036410|scleral icterusnull|Sclera|Anatomy|false|false|C1547225;C0240962;C0022346|scleralnull|Icterus|Finding|false|false|C0036410|icterusnull|Icterus <Icteridae>|Entity|false|false||icterusnull|null|LabModifier|false|false||icterusnull|MAS1L gene|Finding|true|false||MRGnull|Pulmonary ventilator management|Procedure|false|false||PULMnull|Basilar Rales|Finding|false|false||crackles
null|Rales|Finding|false|false||cracklesnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false|C0449202;C0000726|ABDnull|ABD (body structure)|Anatomy|false|false|C3811055|ABD
null|Abdomen|Anatomy|false|false|C3811055|ABDnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|Dilated|Finding|false|false||distendednull|Distended|Modifier|false|false||distendednull|Tender|Modifier|false|false||tendernull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Obvious|Modifier|false|false||obviousnull|Collateral branch of vessel|Anatomy|false|false|C0398102|collateralnull|Collateral|Modifier|false|false||collateralnull|Procedure on vein|Procedure|false|false|C1275670;C0042449|veinsnull|Veins|Anatomy|false|false|C0398102|veinsnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Limb structure|Anatomy|false|false||LIMBSnull|Sequence Chromatogram|Finding|false|false||Tracenull|Trace Dosing Unit|LabModifier|false|false||Trace
null|trace amount|LabModifier|false|false||Trace
null|unknown - trace|LabModifier|false|false||Tracenull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Tremor|Finding|true|false||tremorsnull|Asterixis|Finding|true|false||asterixisnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765|SKIN
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765|SKINnull|Skin Specimen Source Code|Finding|false|false|C1123023;C4520765|SKIN
null|Skin Specimen|Finding|false|false|C1123023;C4520765|SKINnull|Skin, Human|Anatomy|false|false|C0178298;C0496955;C1546781;C0444099|SKIN
null|Skin|Anatomy|false|false|C0178298;C0496955;C1546781;C0444099|SKINnull|Skin rash|Finding|true|false||rashes
null|Exanthema|Finding|true|false||rashesnull|Impaired skin integrity|Finding|true|false|C1123023;C4520765|skin breakdown
null|Broken skin|Finding|true|false|C1123023;C4520765|skin breakdownnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765|skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765|skinnull|Skin Specimen Source Code|Finding|false|false|C1123023;C4520765|skin
null|Skin Specimen|Finding|false|false|C1123023;C4520765|skinnull|Skin, Human|Anatomy|false|false|C1546781;C0444099;C4048181;C0150077;C1265875;C0699900;C0178298;C0496955|skin
null|Skin|Anatomy|false|false|C1546781;C0444099;C4048181;C0150077;C1265875;C0699900;C0178298;C0496955|skinnull|Disintegration (morphologic abnormality)|Disorder|true|false|C1123023;C4520765|breakdownnull|Catabolism|Finding|true|false|C1123023;C4520765|breakdownnull|Scattered|Modifier|false|false||scatterednull|Ecchymosis|Finding|true|false||ecchymosesnull|Puncture wound|Disorder|false|false||puncturenull|Puncture procedure|Procedure|false|false||puncturenull|Site|Modifier|false|false||sitesnull|Neurology speciality|Title|false|false||NEUROnull|Neurologic (qualifier value)|Modifier|false|false||NEUROnull|Pronator drift|Finding|true|false||pronator driftnull|Observation of reflex|Finding|true|false||reflexes
null|Reflex action|Finding|true|false||reflexesnull|Examination of reflexes|Procedure|true|false||reflexesnull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Lower Extremity|Anatomy|false|false|C2003888|lower extremitiesnull|Body Site Modifier - Lower|Anatomy|false|false|C2003888|lowernull|Lower (action)|Event|false|false|C0023216;C0278454;C0015385;C1548802|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|All extremities|Anatomy|false|false|C2003888|extremities
null|Limb structure|Anatomy|false|false|C2003888|extremitiesnull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false||Bloodnull|peripheral blood|Finding|false|false||Blood
null|Blood|Finding|false|false||Blood
null|In Blood|Finding|false|false||Bloodnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||HGB
null|Hemoglobin|Drug|false|false||HGBnull|CYGB gene|Finding|false|false||HGBnull|Hemoglobin concentration|Lab|false|false||HGBnull|Hemopoietic stem cell transplant|Procedure|false|false||HCT
null|Hematocrit Measurement|Procedure|false|false||HCTnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||PLTnull|Count Dosing Unit|LabModifier|false|false||COUNT
null|Count|LabModifier|false|false||COUNTnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Albumin|Drug|false|false||ALBUMIN
null|Albumins|Drug|false|false||ALBUMIN
null|Albumins|Drug|false|false||ALBUMIN
null|Albumin|Drug|false|false||ALBUMINnull|Albumin metabolic function|Finding|false|false||ALBUMIN
null|ALB gene|Finding|false|false||ALBUMINnull|Albumin measurement|Procedure|false|false||ALBUMINnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGPT - Glutamate pyruvate transaminase|Drug|false|false||SGPT
null|SGPT - Glutamate pyruvate transaminase|Drug|false|false||SGPTnull|GPT gene|Finding|false|false||SGPTnull|Serum Alanine Transaminase Test|Procedure|false|false||SGPTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|ASTnull|Atypical Spitz Nevus|Disorder|false|false|C1185650|ASTnull|SLC17A5 wt Allele|Finding|false|false|C1185650|AST
null|SLC17A5 gene|Finding|false|false|C1185650|AST
null|GOT1 gene|Finding|false|false|C1185650|ASTnull|Asterion|Anatomy|false|false|C1415181;C4522245;C1415181;C1420113;C5960784;C0201899;C0004002;C0242192;C1121182|ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||SGOT
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||SGOTnull|GOT1 gene|Finding|false|false|C1185650|SGOTnull|Aspartate aminotransferase measurement|Procedure|false|false|C1185650|SGOTnull|Alkaline Phosphatase|Drug|false|false||ALK PHOS
null|Alkaline Phosphatase|Drug|false|false||ALK PHOSnull|Alkaline phosphatase measurement|Procedure|false|false||ALK PHOSnull|ALK protein, human|Drug|false|false||ALK
null|ALK protein, human|Drug|false|false||ALKnull|ALK protein, human|Finding|false|false||ALK
null|ALK gene|Finding|false|false||ALK
null|ALK wt Allele|Finding|false|false||ALKnull|Phos <Photinae>|Entity|false|false||PHOSnull|Ascitic Fluid|Finding|false|false||Ascitic Fluidnull|Ascitic|Modifier|false|false||Asciticnull|fluid - substance|Drug|false|false||Fluid
null|Liquid substance|Drug|false|false||Fluidnull|Fluid Specimen Code|Finding|false|false||Fluidnull|Fluid behavior|Modifier|false|false||Fluidnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|5'-Inosinic acid, 2'-deoxy-2'-fluoro-, homopolymer|Drug|false|false||POLYS
null|Poly A|Drug|false|false||POLYSnull|Lymph|Finding|false|false||LYMPHSnull|Monos|Drug|false|false||MONOS
null|Mono-S|Drug|false|false||MONOS
null|Monos|Drug|false|false||MONOSnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||EOS
null|Familial eosinophilia|Disorder|false|false||EOSnull|PRSS33 gene|Finding|false|false||EOS
null|IKZF4 gene|Finding|false|false||EOSnull|Eos <Loriini>|Entity|false|false||EOSnull|SLC6A7 gene|Finding|false|false||PROTnull|Lactate Dehydrogenase|Drug|false|false||LDH
null|Lactate Dehydrogenase|Drug|false|false||LDHnull|Lifetime Drinking History|Finding|false|false||LDHnull|Lactate dehydrogenase measurement|Procedure|false|false||LDHnull|Albumin|Drug|false|false||ALBUMIN
null|Albumins|Drug|false|false||ALBUMIN
null|Albumins|Drug|false|false||ALBUMIN
null|Albumin|Drug|false|false||ALBUMINnull|Albumin metabolic function|Finding|false|false||ALBUMIN
null|ALB gene|Finding|false|false||ALBUMINnull|Albumin measurement|Procedure|false|false||ALBUMINnull|Ascitic Fluid|Finding|false|false||Ascitic Fluidnull|Ascitic|Modifier|false|false||Asciticnull|fluid - substance|Drug|false|false||Fluid
null|Liquid substance|Drug|false|false||Fluidnull|Fluid Specimen Code|Finding|false|false||Fluidnull|Fluid behavior|Modifier|false|false||Fluidnull|Leukocytes|Anatomy|false|false||WBCnull|NACC2 wt Allele|Finding|false|false||RBB
null|NACC2 gene|Finding|false|false||RBBnull|5'-Inosinic acid, 2'-deoxy-2'-fluoro-, homopolymer|Drug|false|false||POLYS
null|Poly A|Drug|false|false||POLYSnull|Lymph|Finding|false|false||LYMPHSnull|Monos|Drug|false|false||MONOS
null|Mono-S|Drug|false|false||MONOS
null|Monos|Drug|false|false||MONOSnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||EOS
null|Familial eosinophilia|Disorder|false|false||EOSnull|PRSS33 gene|Finding|false|false||EOS
null|IKZF4 gene|Finding|false|false||EOSnull|Eos <Loriini>|Entity|false|false||EOSnull|Blood and lymphatic system disorders|Disorder|false|false||Bloodnull|peripheral blood|Finding|false|false||Blood
null|Blood|Finding|false|false||Blood
null|In Blood|Finding|false|false||Bloodnull|Leukocytes|Anatomy|false|false|C0472699;C0018935|WBCnull|Hemopoietic stem cell transplant|Procedure|false|false|C0023516|HCT
null|Hematocrit Measurement|Procedure|false|false|C0023516|HCTnull|radiology referral type|Finding|false|false||RADIOLOGY
null|Radiology Section ID|Finding|false|false||RADIOLOGY
null|Encounter due to radiological examination|Finding|false|false||RADIOLOGYnull|Radiology studies|Procedure|false|false||RADIOLOGY
null|Diagnostic radiologic examination|Procedure|false|false||RADIOLOGY
null|Radiographic imaging procedure|Procedure|false|false||RADIOLOGYnull|Radiology Specialty|Title|false|false||RADIOLOGYnull|Lumbo-sacral|Anatomy|false|false||Lumbo-sacralnull|Sacral Region|Anatomy|false|false||sacral
null|Bone structure of sacrum|Anatomy|false|false||sacralnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false|C0549207|evidencenull|Osteomyelitis|Disorder|true|false|C0549207|osteomyelitisnull|Bone structure of spine|Anatomy|false|false|C0029443;C3887511|vertebralnull|Compression fracture|Finding|false|false||compression fracturenull|null|Finding|false|false||compression
null|Compressed structure|Finding|false|false||compressionnull|Compression Therapy|Procedure|false|false||compression
null|Data Compression|Procedure|false|false||compressionnull|Compression|Phenomenon|false|false||compressionnull|Fracture|Disorder|false|false||fracturenull|BRIEF Health Literacy Screening Tool|Finding|false|false||Brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||Briefnull|Brief|Time|false|false||Briefnull|Shortened|Modifier|false|false||Briefnull|Hospital course|Finding|false|false||Hospital Coursenull|null|Attribute|false|false||Hospital Coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||Coursenull|Abdomen distended|Finding|false|false|C0000726|Abdominal distentionnull|Abdomen|Anatomy|false|false|C1549543;C0030193;C3714614;C0012359;C0000731|Abdominalnull|Abdominal (qualifier value)|Modifier|false|false||Abdominalnull|Distention|Finding|false|false|C0000726|distention
null|Pathological Dilatation|Finding|false|false|C0000726|distentionnull|Administration Method - Pain|Finding|false|false|C0000726|pain
null|Pain|Finding|false|false|C0000726|painnull|null|Attribute|false|false||painnull|Concern|Finding|false|false||concernnull|Spontaneous|Finding|false|false||spontaneousnull|Acute bacterial peritonitis|Disorder|false|false||bacterial peritonitis
null|Bacterial peritonitis|Disorder|false|false||bacterial peritonitisnull|Bacterial|Modifier|false|false||bacterialnull|Peritonitis|Finding|false|false||peritonitisnull|ceftriaxone|Drug|false|false||ceftriaxone
null|ceftriaxone|Drug|false|false||ceftriaxonenull|Diagnostic agents|Drug|false|false||diagnosticnull|Location Service Code - Diagnostic|Finding|false|false||diagnostic
null|Diagnostic|Finding|false|false||diagnosticnull|Diagnostic dental procedure|Procedure|false|false||diagnostic
null|Diagnosis|Procedure|false|false||diagnosticnull|Paracentesis|Procedure|false|false||paracentesisnull|Ascitic Fluid|Finding|false|false||Ascitic fluidnull|Ascitic|Modifier|false|false||Asciticnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|analysis aspect|Finding|false|false||analysisnull|Analysis of substances|Procedure|false|false||analysis
null|Analysis|Procedure|false|false||analysisnull|acute spontaneous bacterial peritonitis|Disorder|false|false||Spontaneous bacterial peritonitis
null|Primary bacterial peritonitis|Disorder|false|false||Spontaneous bacterial peritonitisnull|Spontaneous|Finding|false|false||Spontaneousnull|Acute bacterial peritonitis|Disorder|false|false||bacterial peritonitis
null|Bacterial peritonitis|Disorder|false|false||bacterial peritonitisnull|Bacterial|Modifier|false|false||bacterialnull|Peritonitis|Finding|false|false||peritonitisnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Cell Count|Procedure|false|false|C0007634|cell countnull|CELP gene|Finding|false|false|C0007634|cell
null|CEL gene|Finding|false|false|C0007634|cellnull|Cells|Anatomy|false|false|C0007584;C1413336;C1413337|cellnull|Cell Device|Device|false|false||cell
null|Cellular Phone|Device|false|false||cellnull|Cell (compartment)|Modifier|false|false||cellnull|Count Dosing Unit|LabModifier|false|false||count
null|Count|LabModifier|false|false||countnull|Leukocytes|Anatomy|false|false||WBCnull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|Volume (publication)|Finding|false|false||volumenull|Volume|LabModifier|false|false||volumenull|Paracentesis|Procedure|false|false||paracentesisnull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|Procedure (set of actions)|Finding|false|false||procedurenull|Interventional procedure|Procedure|false|false||procedurenull|null|Attribute|false|false||procedurenull|Act Class - procedure|Event|false|false||procedurenull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|abdomennull|Abdomen problem|Finding|false|false|C0230168;C0000726|abdomennull|Abdomen|Anatomy|false|false|C0153662;C0941288|abdomen
null|Abdominal Cavity|Anatomy|false|false|C0153662;C0941288|abdomennull|Smaller|Modifier|false|false||lessnull|Less Than|LabModifier|false|false||lessnull|Dilated|Finding|false|false||distendednull|Distended|Modifier|false|false||distendednull|Smaller|Modifier|false|false||lessnull|Less Than|LabModifier|false|false||lessnull|Pain|Finding|false|false||painfulnull|fluid - substance|Drug|false|false||Fluid
null|Liquid substance|Drug|false|false||Fluidnull|Fluid Specimen Code|Finding|false|false||Fluidnull|Fluid behavior|Modifier|false|false||Fluidnull|analysis aspect|Finding|false|false||analysisnull|Analysis of substances|Procedure|false|false||analysis
null|Analysis|Procedure|false|false||analysisnull|Androgen Binding Protein|Drug|true|false||SBP
null|Androgen Binding Protein|Drug|true|false||SBPnull|CCHCR1 wt Allele|Finding|true|false||SBP
null|SHBG wt Allele|Finding|true|false||SBPnull|Systolic blood pressure measurement|Procedure|true|false||SBPnull|Systolic Pressure|Attribute|true|false||SBPnull|Hepatitis, Alcoholic|Disorder|false|false||Alcoholic hepatitisnull|Alcoholics|Subject|false|false||Alcoholicnull|Hepatitis A|Disorder|false|false||hepatitis
null|Hepatitis|Disorder|false|false||hepatitisnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|false|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|false|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|livernull|Benign neoplasm of liver|Disorder|false|false|C4037986;C1278929;C0023884|liver
null|Liver diseases|Disorder|false|false|C4037986;C1278929;C0023884|livernull|Liver problem|Finding|false|false|C4037986;C1278929;C0023884|livernull|Procedures on liver|Procedure|false|false|C4037986;C1278929;C0023884|livernull|Abdomen>Liver|Anatomy|false|false|C0023895;C0496870;C0721399;C0023899;C0577060;C0872387;C0598463;C0542341;C1705273;C0031843|liver
null|null|Anatomy|false|false|C0023895;C0496870;C0721399;C0023899;C0577060;C0872387;C0598463;C0542341;C1705273;C0031843|liver
null|Liver|Anatomy|false|false|C0023895;C0496870;C0721399;C0023899;C0577060;C0872387;C0598463;C0542341;C1705273;C0031843|livernull|Synthesis|Event|false|false||syntheticnull|Function (attribute)|Finding|false|false|C4037986;C1278929;C0023884|function
null|physiological aspects|Finding|false|false|C4037986;C1278929;C0023884|function
null|Mathematical Operator|Finding|false|false|C4037986;C1278929;C0023884|function
null|Functional Status|Finding|false|false|C4037986;C1278929;C0023884|functionnull|Function Axis|Subject|false|false||functionnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|GDC Regimen Terminology|Finding|false|false||regimennull|Treatment Protocols|Procedure|false|false||regimennull|lactulose|Drug|false|false||lactulose
null|lactulose|Drug|false|false||lactulosenull|Urine Specimen Collection|Procedure|false|false||urine collectionnull|Portion of urine|Finding|false|false||urine
null|null|Finding|false|false||urine
null|Urine|Finding|false|false||urine
null|In Urine|Finding|false|false||urine
null|Urine specimen|Finding|false|false||urinenull|Collection Object - UML Entity|Finding|false|false||collection
null|Item Collection|Finding|false|false||collection
null|Collections (publication)|Finding|false|false||collection
null|Collection (action)|Finding|false|false||collectionnull|copper|Drug|false|false||copper
null|copper|Drug|false|false||copper
null|copper|Drug|false|false||coppernull|Copper measurement|Procedure|false|false||coppernull|Disease|Disorder|false|false||diseasenull|Leukocytosis|Disorder|false|false||Leukocytosisnull|Blood leukocyte number above reference range|Finding|false|false||Leukocytosisnull|Low grade fever|Finding|false|false||mild fevernull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Presentation|Finding|false|false||presentationnull|Aspects of signs|Finding|true|false||signs
null|Physical findings|Finding|true|false||signsnull|Manufactured sign|Device|true|false||signsnull|Symptoms aspect|Finding|true|false||symptoms
null|Symptoms|Finding|true|false||symptomsnull|Communicable Diseases|Disorder|true|false||infectionnull|Infection|Finding|true|false||infectionnull|Urine culture|Procedure|false|false||Urine culturenull|Portion of urine|Finding|false|false||Urine
null|null|Finding|false|false||Urine
null|Urine|Finding|false|false||Urine
null|In Urine|Finding|false|false||Urine
null|Urine specimen|Finding|false|false||Urinenull|Culture Dose Form|Drug|false|false||culturenull|Culture (Anthropological)|Finding|false|false||culture
null|Cultural aspects|Finding|false|false||culturenull|Microbial culture (procedure)|Procedure|false|false||culture
null|Laboratory culture|Procedure|false|false||culturenull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|Contamination|Finding|false|false||contaminationnull|adulteration|Phenomenon|false|false||contaminationnull|Specimen Reject Reason - Contamination|Modifier|false|false||contaminationnull|arrival - ActRelationshipType|Finding|false|false||arrivalnull|null|Event|false|false||arrivalnull|Floor (anatomic)|Anatomy|false|false|C1547311;C0886414|floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Body temperature measurement|Procedure|false|false|C3714591|temperaturenull|Body Temperature|Subject|false|false||temperaturenull|Temperature|LabModifier|false|false||temperaturenull|Patient Condition Code - Stable|Finding|false|false|C3714591|stablenull|Stable status|Modifier|false|false||stablenull|Leukocytes|Anatomy|false|false||WBCnull|Hospitalization|Procedure|false|false||hospitalizationnull|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Tachycardia by ECG Finding|Finding|false|false||Tachycardia
null|Tachycardia|Finding|false|false||Tachycardianull|null|Finding|false|false|C4037974;C0018787|heart ratenull|examination of heart rate|Procedure|false|false|C4037974;C0018787|heart ratenull|heart rate|Attribute|false|false|C4037974;C0018787|heart rate
null|null|Attribute|false|false|C4037974;C0018787|heart ratenull|Mean Heart Rate|LabModifier|false|false||heart ratenull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C0018810;C0488794;C2041121;C0795691;C1549480;C0153957;C0153500;C0871208;C2197023|heart
null|Heart|Anatomy|false|false|C0018810;C0488794;C2041121;C0795691;C1549480;C0153957;C0153500;C0871208;C2197023|heartnull|Amount type - Rate|Finding|false|false|C4037974;C0018787|ratenull|Rating (action)|Event|false|false|C4037974;C0018787|ratenull|Rate|LabModifier|false|false||ratenull|Hospitalization|Procedure|false|false||hospitalizationnull|Language Ability Proficiency - Good|Finding|false|false||good
null|Language Proficiency - Good|Finding|false|false||goodnull|Specimen Quality - Good|Modifier|false|false||good
null|Good|Modifier|false|false||goodnull|Alveolar ventilation function|Finding|false|false||oxygenation
null|Cell Respiration|Finding|false|false||oxygenationnull|Complaint (finding)|Finding|true|false||complaintsnull|Dyspnea|Finding|false|false||SOBnull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C2926613;C0008031;C0741025;C1549543;C0030193|chest
null|Anterior thoracic region|Anatomy|false|false|C2926613;C0008031;C0741025;C1549543;C0030193|chestnull|Administration Method - Pain|Finding|false|false|C1527391;C0817096|pain
null|Pain|Finding|false|false|C1527391;C0817096|painnull|null|Attribute|false|false||painnull|Palpitations|Finding|false|false||palpitationsnull|most likely|Finding|false|false||most likelynull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Science of Etiology|Finding|false|false||etiology
null|Etiology aspects|Finding|false|false||etiology
null|Etiology|Finding|false|false||etiologynull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Anxiety Disorders|Disorder|false|false||anxiety
null|Anxiety|Disorder|false|false||anxietynull|Anxiety symptoms|Finding|false|false||anxietynull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Intravascular Route of Administration|Finding|false|false||intravascularnull|Intravascular|Modifier|false|false||intravascularnull|Volume (publication)|Finding|false|false||volumenull|Volume|LabModifier|false|false||volumenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Back Pain|Finding|false|false||Back painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Lumbosacral spine|Anatomy|false|false|C4019020;C0150920|Lumbosacral spinenull|Lumbosacral|Modifier|false|false||Lumbosacralnull|Spine Problem|Finding|false|false|C0223603;C2752558;C0037949|spinenull|Neuron spine|Anatomy|false|false|C4019020;C0150920|spine
null|Vertebral column|Anatomy|false|false|C4019020;C0150920|spinenull|Film Dosage Form|Drug|false|false||film
null|film - layer|Drug|false|false||filmnull|null|Finding|false|false|C2752558;C0037949;C0223603|filmnull|film (photographic)|Device|false|false||film
null|Film Device|Device|false|false||film
null|Film Container Cap|Device|false|false||filmnull|Film (unit of presentation)|LabModifier|false|false||film
null|Film Dosing Unit|LabModifier|false|false||filmnull|Abnormality of the skeletal system|Disorder|true|false||skeletal abnormalitiesnull|Skeletal|Modifier|false|false||skeletalnull|Congenital Abnormality|Disorder|true|false||abnormalitiesnull|teratologic|Finding|true|false||abnormalitiesnull|Compression fracture of vertebral column|Finding|false|false|C0549207|vertebral compression fracturenull|Compression fracture of vertebral column|Finding|false|false|C0549207|vertebral compressionnull|Bone structure of spine|Anatomy|false|false|C0728907;C1257972;C0565514;C0016658;C0029443;C0262431;C0332459;C4551657;C0521169;C0262431|vertebralnull|Compression fracture|Finding|false|false|C0549207|compression fracturenull|null|Finding|false|false|C0549207|compression
null|Compressed structure|Finding|false|false|C0549207|compressionnull|Compression Therapy|Procedure|false|false|C0549207|compression
null|Data Compression|Procedure|false|false|C0549207|compressionnull|Compression|Phenomenon|false|false|C0549207|compressionnull|Fracture|Disorder|false|false|C0549207|fracturenull|Osteomyelitis|Disorder|false|false|C0549207|osteomyelitisnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Hospitalization|Procedure|false|false||hospitalizationnull|oxycodone|Drug|false|false||oxycodone
null|oxycodone|Drug|false|false||oxycodonenull|Oxycodone measurement|Procedure|false|false||oxycodonenull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Primary Care Provider - Provider role|Finding|false|false||primary care providernull|null|Attribute|false|false||primary care providernull|Primary care provider|Subject|false|false||primary care providernull|Location Service Code - Primary Care|Finding|false|false||primary carenull|Primary Health Care|Procedure|false|false||primary carenull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Transaction counts and value totals - provider|Finding|false|false||provider
null|Provider|Finding|false|false||providernull|Disease Management|Procedure|false|false||managementnull|Management Occupations|Subject|false|false||managementnull|Management procedure|Event|false|false||management
null|Administration occupational activities|Event|false|false||managementnull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Diet (animal life circumstance)|Drug|false|false||Diet
null|Diet|Drug|false|false||Dietnull|diet - supply|Finding|false|false||Dietnull|Diet therapy|Procedure|false|false||Dietnull|Sodium decreased|Finding|false|false||Low sodiumnull|Low sodium diet|Procedure|false|false||Low sodiumnull|IPSS-R Risk Category Low|Finding|false|false||Low
null|IPSS Risk Category Low|Finding|false|false||Low
null|low confidentiality|Finding|false|false||Lownull|Low - MessageWaitingPriority|Modifier|false|false||Low
null|low|Modifier|false|false||Low
null|low exposure|Modifier|false|false||Lownull|null|LabModifier|false|false||Lownull|Sodium supplements|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|Sodium Drug Class|Drug|false|false||sodiumnull|Sodium metabolic function|Finding|false|false||sodiumnull|Sodium measurement|Procedure|false|false||sodiumnull|per day|Time|false|false||/daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Fluid restriction|Procedure|false|false||fluid restrictionnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Restricted|Finding|false|false||restrictionnull|per day|Time|false|false||/daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|MDF Attribute Type - Code|Finding|false|false||Code
null|A Codes|Finding|false|false||Code
null|Code|Finding|false|false||Codenull|Coding|Event|false|false||Codenull|Full|Modifier|false|false||Fullnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|amitriptyline|Drug|false|false||AMITRIPTYLINE
null|amitriptyline|Drug|false|false||AMITRIPTYLINEnull|oxycodone|Drug|false|false||OXYCODONE
null|oxycodone|Drug|false|false||OXYCODONEnull|Oxycodone measurement|Procedure|false|false||OXYCODONEnull|Every eight hours|Time|false|false||Q8Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Thiamine Drug Class|Drug|false|false||Thiamine
null|thiamine|Drug|false|false||Thiamine
null|thiamine|Drug|false|false||Thiamine
null|thiamine|Drug|false|false||Thiamine
null|Thiamine Drug Class|Drug|false|false||Thiaminenull|Thiamine measurement|Procedure|false|false||Thiaminenull|Daily|Time|false|false||dailynull|folic acid|Drug|false|false||Folic acid
null|folic acid|Drug|false|false||Folic acid
null|folic acid|Drug|false|false||Folic acidnull|Folic acid measurement|Procedure|false|false||Folic acidnull|Daily|Time|false|false||dailynull|MVI Regimen|Procedure|false|false||MVInull|Daily|Time|false|false||dailynull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|thiamine hydrochloride|Drug|false|false||Thiamine HCl
null|thiamine hydrochloride|Drug|false|false||Thiamine HCl
null|thiamine hydrochloride|Drug|false|false||Thiamine HClnull|Thiamine Drug Class|Drug|false|false||Thiamine
null|thiamine|Drug|false|false||Thiamine
null|thiamine|Drug|false|false||Thiamine
null|thiamine|Drug|false|false||Thiamine
null|Thiamine Drug Class|Drug|false|false||Thiaminenull|Thiamine measurement|Procedure|false|false||Thiaminenull|Flinders medical centre-7 marker|Drug|false|false||HCl
null|hydrochloride|Drug|false|false||HCl
null|hydrochloride|Drug|false|false||HClnull|Hairy Cell Leukemia|Disorder|false|false||HClnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|folic acid|Drug|false|false||Folic Acid
null|folic acid|Drug|false|false||Folic Acid
null|folic acid|Drug|false|false||Folic Acidnull|Folic acid measurement|Procedure|false|false||Folic Acidnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|amitriptyline|Drug|false|false||Amitriptyline
null|amitriptyline|Drug|false|false||Amitriptylinenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Bedtime (qualifier value)|Time|false|false||bedtime
null|Once a day, at bedtime|Time|false|false||bedtimenull|Multivitamin tablet|Drug|false|false||Multivitamin     Tabletnull|Multivitamin preparation|Drug|false|false||Multivitamin
null|Multivitamin preparation|Drug|false|false||Multivitamin
null|Multivitamin preparation|Drug|false|false||Multivitaminnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|lactulose|Drug|true|false||Lactulose
null|lactulose|Drug|true|false||Lactulosenull|gram|LabModifier|false|false||gramnull|Syrup Drug Form|Drug|true|false||Syrup
null|Syrup (dietary)|Drug|true|false||Syrupnull|Receptors, Antigen, B-Cell|Drug|false|false|C0262329|Sig
null|Receptors, Antigen, B-Cell|Drug|false|false|C0262329|Signull|Receptors, Antigen, B-Cell|Finding|false|false|C0262329|Signull|Short insular gyrus|Anatomy|false|false|C0034789;C0034789|Signull|Surveillance Implementation Group|Entity|false|false||Sig
null|Staphylococcus intermedius group|Entity|false|false||Signull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|oxycodone|Drug|false|false||Oxycodone
null|oxycodone|Drug|false|false||Oxycodonenull|Oxycodone measurement|Procedure|false|false||Oxycodonenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Hour|Time|false|false||hoursnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|True primary (qualifier value)|Time|false|false||Primarynull|Primary|Modifier|false|false||Primarynull|Ascites|Disorder|false|false||Ascitesnull|Peritoneal Effusion|Finding|false|false||Ascitesnull|Portal Hypertension|Disorder|false|false|C0205054|Portal hypertensionnull|Hepatic|Anatomy|false|false|C0020538;C0020541|Portalnull|Hypertensive disease|Disorder|false|false|C0205054|hypertensionnull|Hepatitis, Alcoholic|Disorder|false|false||Alcoholic hepatitisnull|Alcoholics|Subject|false|false||Alcoholicnull|Hepatitis A|Disorder|false|false||hepatitis
null|Hepatitis|Disorder|false|false||hepatitisnull|Neoplasm Metastasis|Disorder|false|false||Secondarynull|metastatic qualifier|Finding|false|false||Secondarynull|Secondary to|Modifier|false|false||Secondarynull|second (number)|LabModifier|false|false||Secondarynull|Chronic back pain|Finding|false|false||Chronic back painnull|Chronic - Admission Level of Care Code|Finding|false|false||Chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||Chronicnull|chronic|Time|false|false||Chronicnull|Back Pain|Finding|false|false||back painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Disease|Disorder|false|false||Conditionnull|Logical Condition|Finding|false|false||Conditionnull|null|Attribute|false|false||Conditionnull|Condition|Modifier|false|false||Conditionnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Oriented to place|Finding|false|false||Orientednull|Orientation, Spatial|Modifier|false|false||Orientednull|Without Help|Finding|false|false||without helpnull|Help document|Finding|true|false||helpnull|Assisted (qualifier value)|Modifier|false|false||helpnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Apyrexial|Finding|false|false||afebrilenull|Discharge instructions|Finding|false|false||Discharge Instructionsnull|hospital discharge instructions (treatment)|Procedure|false|false||Discharge Instructionsnull|null|Attribute|false|false||Discharge Instructionsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|Complaint (finding)|Finding|false|false|C0000726|complaintsnull|Increasing (qualifier value)|Finding|false|false||increasingnull|Abdominal distention and pain|Finding|false|false|C0000726|abdominal distention and painnull|Abdomen distended|Finding|false|false|C0000726|abdominal distentionnull|Abdomen|Anatomy|false|false|C2749840;C3714614;C0012359;C5441521;C0000731;C1549543;C0030193|abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Distention|Finding|false|false|C0000726|distention
null|Pathological Dilatation|Finding|false|false|C0000726|distentionnull|Administration Method - Pain|Finding|false|false|C0000726|pain
null|Pain|Finding|false|false|C0000726|painnull|null|Attribute|false|false||painnull|Clinic|Device|false|false||clinic
null|Ambulatory Care Facilities|Device|false|false||clinicnull|Clinic|Entity|false|false||clinic
null|Ambulatory Care Facilities|Entity|false|false||clinicnull|Patient location type - Clinic|Modifier|false|false||clinic
null|Person location type - Clinic|Modifier|false|false||clinicnull|Low grade fever|Finding|false|false||mild fevernull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Tachycardia|Finding|false|false|C4037974;C0018787|fast heart ratenull|Fas-activated serine/threonine kinase activity|Finding|false|false||fast
null|FASTK Gene|Finding|false|false||fast
null|FOXD3-AS1 gene|Finding|false|false||fast
null|FASTK wt Allele|Finding|false|false||fast
null|Fasting|Finding|false|false||fastnull|Rapid|Modifier|false|false||fastnull|null|Finding|false|false|C4037974;C0018787|heart ratenull|examination of heart rate|Procedure|false|false|C4037974;C0018787|heart ratenull|heart rate|Attribute|false|false|C4037974;C0018787|heart rate
null|null|Attribute|false|false|C4037974;C0018787|heart ratenull|Mean Heart Rate|LabModifier|false|false||heart ratenull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C2041121;C0153957;C0153500;C0795691;C2197023;C0039231;C0018810;C0488794|heart
null|Heart|Anatomy|false|false|C2041121;C0153957;C0153500;C0795691;C2197023;C0039231;C0018810;C0488794|heartnull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|White blood count|Finding|false|false||white blood countnull|White (population group)|Subject|false|false||white
null|Caucasian|Subject|false|false||white
null|Caucasians|Subject|false|false||whitenull|White color|Modifier|false|false||whitenull|Blood Cell Count|Procedure|false|false||blood countnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Count Dosing Unit|LabModifier|false|false||count
null|Count|LabModifier|false|false||countnull|Consent Non-Disclosure Reason - Emergency|Finding|false|false||emergency
null|Admission Type - Emergency|Finding|false|false||emergency
null|Referral category - Emergency|Finding|false|false||emergency
null|Emergencies [Disease/Finding]|Finding|false|false||emergency
null|Consent Bypass Reason - Emergency|Finding|false|false||emergency
null|Level of Care - Emergency|Finding|false|false||emergency
null|Certification patient type - Emergency|Finding|false|false||emergency
null|Encounter Admission Source - emergency|Finding|false|false||emergency
null|Patient Class - Emergency|Finding|false|false||emergency
null|Visit Priority Code - Emergency|Finding|false|false||emergencynull|emergency encounter|Procedure|false|false||emergencynull|Emergency Situation|Phenomenon|false|false||emergencynull|Specialty Type - Emergency|Title|false|false||emergencynull|Bale out|Time|false|false||emergencynull|Department - No suggested values defined|Finding|false|false||department
null|Organization Unit Type - Department|Finding|false|false||department
null|Department - Charge type|Finding|false|false||departmentnull|Department|Entity|false|false||departmentnull|Patient location type - Department|Modifier|false|false||department
null|Department - Person location type|Modifier|false|false||departmentnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Further|Modifier|false|false||furthernull|Hospitalization|Procedure|false|false||hospitalizationnull|Ascitic Fluid|Finding|false|false||ascitic fluidnull|Ascitic|Modifier|false|false||asciticnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|What subject filter - Result|Finding|false|false||result
null|Result|Finding|false|false||result
null|Experimental Result|Finding|false|false||resultnull|Communicable Diseases|Disorder|true|false||infectionnull|Infection|Finding|true|false||infectionnull|Ascitic Fluid|Finding|false|false||ascitic fluidnull|Ascitic|Modifier|false|false||asciticnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|abdomennull|Abdomen problem|Finding|false|false|C0230168;C0000726|abdomennull|Abdomen|Anatomy|false|false|C0153662;C0034115;C0941288|abdomen
null|Abdominal Cavity|Anatomy|false|false|C0153662;C0034115;C0941288|abdomennull|Paracentesis|Procedure|false|false|C0230168;C0000726|paracentesisnull|Portion of urine|Finding|false|false||urine
null|null|Finding|false|false||urine
null|Urine|Finding|false|false||urine
null|In Urine|Finding|false|false||urine
null|Urine specimen|Finding|false|false||urinenull|Collection Object - UML Entity|Finding|false|false||collection
null|Item Collection|Finding|false|false||collection
null|Collections (publication)|Finding|false|false||collection
null|Collection (action)|Finding|false|false||collectionnull|copper|Drug|false|false||copper
null|copper|Drug|false|false||copper
null|copper|Drug|false|false||coppernull|Copper measurement|Procedure|false|false||coppernull|Potential|Modifier|false|false||potentialnull|Etiology aspects|Finding|false|false||causes
null|Etiology|Finding|false|false||causesnull|Liver diseases|Disorder|false|false|C4037986;C1278929;C0023884|liver disease
null|Hepatobiliary Disorder|Disorder|false|false|C4037986;C1278929;C0023884|liver diseasenull|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|false|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|false|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|livernull|Benign neoplasm of liver|Disorder|false|false|C4037986;C1278929;C0023884|liver
null|Liver diseases|Disorder|false|false|C4037986;C1278929;C0023884|livernull|Liver problem|Finding|false|false|C4037986;C1278929;C0023884|livernull|Procedures on liver|Procedure|false|false|C4037986;C1278929;C0023884|livernull|Abdomen>Liver|Anatomy|false|false|C0872387;C0267792;C0023895;C0012634;C0577060;C0721399;C0023899;C0023895;C0496870|liver
null|null|Anatomy|false|false|C0872387;C0267792;C0023895;C0012634;C0577060;C0721399;C0023899;C0023895;C0496870|liver
null|Liver|Anatomy|false|false|C0872387;C0267792;C0023895;C0012634;C0577060;C0721399;C0023899;C0023895;C0496870|livernull|Disease|Disorder|false|false|C4037986;C1278929;C0023884|diseasenull|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|false|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|false|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|livernull|Benign neoplasm of liver|Disorder|false|false|C4037986;C1278929;C0023884|liver
null|Liver diseases|Disorder|false|false|C4037986;C1278929;C0023884|livernull|Liver problem|Finding|false|false|C4037986;C1278929;C0023884|livernull|Procedures on liver|Procedure|false|false|C4037986;C1278929;C0023884|livernull|Abdomen>Liver|Anatomy|false|false|C0577060;C0023895;C0496870;C0721399;C0023899;C0872387|liver
null|null|Anatomy|false|false|C0577060;C0023895;C0496870;C0721399;C0023899;C0872387|liver
null|Liver|Anatomy|false|false|C0577060;C0023895;C0496870;C0721399;C0023899;C0872387|livernull|Clinic|Device|false|false||clinic
null|Ambulatory Care Facilities|Device|false|false||clinicnull|Clinic|Entity|false|false||clinic
null|Ambulatory Care Facilities|Entity|false|false||clinicnull|Patient location type - Clinic|Modifier|false|false||clinic
null|Person location type - Clinic|Modifier|false|false||clinicnull|Tests (qualifier value)|Finding|false|false||testsnull|Laboratory Procedures|Procedure|false|false||testsnull|Back Pain|Finding|false|false||back painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Hospitalization|Procedure|false|false||hospitalizationnull|X-rays, Homeopathic Preparations|Drug|false|false||x-raysnull|Plain x-ray|Procedure|false|false||x-rays
null|Diagnostic radiologic examination|Procedure|false|false||x-raysnull|Roentgen Rays|Phenomenon|false|false||x-raysnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Fracture|Disorder|true|false||fracturenull|Specimen Type - Bone|Finding|true|false|C1442209;C0262950|bone
null|null|Finding|true|false|C1442209;C0262950|bonenull|Skeletal bone|Anatomy|false|false|C1546560;C1550616|bone
null|XXX bone|Anatomy|false|false|C1546560;C1550616|bonenull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|GDC Regimen Terminology|Finding|false|false||regimennull|Treatment Protocols|Procedure|false|false||regimennull|Primary Care Provider - Provider role|Finding|false|false||primary care providernull|null|Attribute|false|false||primary care providernull|Primary care provider|Subject|false|false||primary care providernull|Location Service Code - Primary Care|Finding|false|false||primary carenull|Primary Health Care|Procedure|false|false||primary carenull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Transaction counts and value totals - provider|Finding|false|false||provider
null|Provider|Finding|false|false||providernull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|lactulose|Drug|false|false||lactulose
null|lactulose|Drug|false|false||lactulosenull|Constipation|Finding|false|false||constipationnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Herbals (publications)|Finding|false|false||herbalnull|Herbal|Modifier|false|false||herbalnull|TONICS|Drug|false|false||tonicnull|Homeopathic Remedies|Drug|false|false||remediesnull|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|false|false|C4037986;C1278929;C0023884|liver
null|liver extract|Drug|false|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|liver
null|Liver brand of Vitamin B 12|Drug|false|false|C4037986;C1278929;C0023884|livernull|Benign neoplasm of liver|Disorder|false|false|C4037986;C1278929;C0023884|liver
null|Liver diseases|Disorder|false|false|C4037986;C1278929;C0023884|livernull|Liver problem|Finding|false|false|C4037986;C1278929;C0023884|livernull|Procedures on liver|Procedure|false|false|C4037986;C1278929;C0023884|livernull|Abdomen>Liver|Anatomy|false|false|C0023895;C0496870;C0577060;C0872387;C0721399;C0023899|liver
null|null|Anatomy|false|false|C0023895;C0496870;C0577060;C0872387;C0721399;C0023899|liver
null|Liver|Anatomy|false|false|C0023895;C0496870;C0577060;C0872387;C0721399;C0023899|livernull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|Therapeutic procedure|Procedure|false|false||therapiesnull|Electrical Current|Phenomenon|false|false||currentnull|Current (present time)|Time|false|false||currentnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Difficult (qualifier value)|Finding|false|false||difficultnull|Laboratory Results|Lab|false|false||laboratory resultsnull|Diagnostic Service Section ID - Laboratory|Finding|false|false||laboratory
null|Laboratory domain|Finding|false|false||laboratory
null|Referral type - Laboratory|Finding|false|false||laboratorynull|null|Attribute|false|false||laboratorynull|Laboratory|Device|false|false||laboratorynull|Laboratory observation|Lab|false|false||laboratorynull|Laboratory|Entity|false|false||laboratorynull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions