 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Procedure|Health Care Activity|SIMPLE_SEGMENT|39,48|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|39,53|false|false|false|C2598112||Admission Date
Finding|Body Substance|SIMPLE_SEGMENT|73,82|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|73,82|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|73,82|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|73,82|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|73,87|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|105,110|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|105,110|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|105,110|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|129,132|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|140,147|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|140,147|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|149,157|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|Allergies|181,190|false|false|false|C1717415||Allergies
Finding|Pathologic Function|Allergies|181,190|false|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|Allergies|193,215|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|Allergies|201,205|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|Allergies|201,205|false|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|Allergies|201,215|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Finding|Functional Concept|Allergies|218,227|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|Chief Complaint|253,260|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|Chief Complaint|253,260|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|Chief Complaint|253,272|false|false|false|C0231807|Dyspnea on exertion|dyspnea on exertion
Finding|Organism Function|Chief Complaint|264,272|false|false|false|C0015264|Exertion|exertion
Finding|Classification|Chief Complaint|275,280|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|281,289|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|281,289|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|293,311|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|302,311|false|false|false|C0945766||Procedure
Event|Occupational Activity|Chief Complaint|302,311|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|302,311|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|302,311|false|false|false|C0184661|Interventional procedure|Procedure
Finding|Conceptual Entity|History of Present Illness|360,367|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|360,367|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|360,367|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|360,370|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|History of Present Illness|374,377|false|false|false|C0020538|Hypertensive disease|HTN
Disorder|Disease or Syndrome|History of Present Illness|379,382|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|379,382|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|History of Present Illness|379,382|false|false|false|C1504769|DFFB protein, human|CAD
Finding|Gene or Genome|History of Present Illness|379,382|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|History of Present Illness|379,382|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|History of Present Illness|379,382|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|379,382|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|History of Present Illness|387,390|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|387,390|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|History of Present Illness|387,390|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|History of Present Illness|387,390|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|History of Present Illness|387,390|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|History of Present Illness|387,390|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Finding|Gene or Genome|History of Present Illness|387,390|false|false|false|C1413980|DES gene|DES
Finding|Functional Concept|History of Present Illness|396,404|false|false|false|C0475224|Ischemic|ischemic
Finding|Organ or Tissue Function|History of Present Illness|413,421|false|false|false|C0039155|Systole|systolic
Finding|Pathologic Function|History of Present Illness|413,433|false|false|false|C0749225|Systolic dysfunction|systolic dysfunction
Disorder|Disease or Syndrome|History of Present Illness|422,433|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Finding|Conceptual Entity|History of Present Illness|422,433|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|History of Present Illness|422,433|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|History of Present Illness|422,433|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Drug|Organic Chemical|History of Present Illness|442,451|false|false|false|C0076840|torsemide|torsemide
Drug|Pharmacologic Substance|History of Present Illness|442,451|false|false|false|C0076840|torsemide|torsemide
Anatomy|Body Location or Region|History of Present Illness|459,462|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|History of Present Illness|459,462|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|History of Present Illness|459,462|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Finding|Finding|History of Present Illness|493,500|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|History of Present Illness|493,500|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|History of Present Illness|493,512|false|false|false|C0231807|Dyspnea on exertion|dyspnea on exertion
Finding|Organism Function|History of Present Illness|504,512|false|false|false|C0015264|Exertion|exertion
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|514,517|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Pathologic Function|History of Present Illness|514,526|false|false|false|C0581394|Swelling of lower limb|leg swelling
Finding|Finding|History of Present Illness|518,526|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|History of Present Illness|518,526|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Attribute|Clinical Attribute|History of Present Illness|535,541|false|false|false|C0944911||weight
Finding|Finding|History of Present Illness|535,541|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|History of Present Illness|535,541|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|History of Present Illness|535,541|false|false|false|C1305866|Weighing patient|weight
Finding|Body Substance|History of Present Illness|559,566|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|559,566|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|559,566|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|583,588|false|false|false|C0018787;C4037974|Chest>Heart;Heart|Heart
Disorder|Neoplastic Process|History of Present Illness|583,588|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|Heart
Finding|Sign or Symptom|History of Present Illness|583,588|false|false|false|C0795691|HEART PROBLEM|Heart
Disorder|Disease or Syndrome|History of Present Illness|583,596|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|Heart Failure
Finding|Functional Concept|History of Present Illness|589,596|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|Failure
Finding|Idea or Concept|History of Present Illness|589,596|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|Failure
Finding|Individual Behavior|History of Present Illness|589,596|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|Failure
Finding|Finding|History of Present Illness|670,677|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|History of Present Illness|670,677|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|History of Present Illness|670,689|false|false|false|C0231807|Dyspnea on exertion|dyspnea on exertion
Finding|Organism Function|History of Present Illness|681,689|false|false|false|C0015264|Exertion|exertion
Disorder|Disease or Syndrome|History of Present Illness|694,697|false|false|false|C1956415|Paroxysmal nocturnal dyspnea|PND
Finding|Gene or Genome|History of Present Illness|694,697|false|false|false|C1417807;C4552608|NPPA gene;NPPA wt Allele|PND
Procedure|Health Care Activity|History of Present Illness|721,736|false|false|false|C0019993|Hospitalization|hospitalization
Anatomy|Body Location or Region|History of Present Illness|741,744|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|History of Present Illness|741,744|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|History of Present Illness|741,744|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Finding|Finding|History of Present Illness|758,762|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|History of Present Illness|758,762|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|History of Present Illness|758,762|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Drug|Organic Chemical|History of Present Illness|791,800|false|false|false|C0076840|torsemide|torsemide
Drug|Pharmacologic Substance|History of Present Illness|791,800|false|false|false|C0076840|torsemide|torsemide
Finding|Functional Concept|History of Present Illness|830,838|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|History of Present Illness|830,838|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|History of Present Illness|851,858|false|false|false|C0019843|Holidays|holiday
Finding|Finding|History of Present Illness|877,881|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|History of Present Illness|877,881|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|History of Present Illness|877,881|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Drug|Chemical Viewed Structurally|History of Present Illness|882,886|false|false|false|C0036140;C0037494;C0206136|Salts;Sodium Chloride, Dietary;sodium chloride|salt
Drug|Food|History of Present Illness|882,886|false|false|false|C0036140;C0037494;C0206136|Salts;Sodium Chloride, Dietary;sodium chloride|salt
Drug|Inorganic Chemical|History of Present Illness|882,886|false|false|false|C0036140;C0037494;C0206136|Salts;Sodium Chloride, Dietary;sodium chloride|salt
Drug|Food|History of Present Illness|887,891|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Finding|Functional Concept|History of Present Illness|887,891|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|History of Present Illness|887,891|false|false|false|C0012159|Diet therapy|diet
Finding|Finding|History of Present Illness|918,925|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|History of Present Illness|918,925|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|History of Present Illness|918,937|false|false|false|C0231807|Dyspnea on exertion|dyspnea on exertion
Finding|Organism Function|History of Present Illness|929,937|false|false|false|C0015264|Exertion|exertion
Drug|Pharmacologic Substance|History of Present Illness|950,960|true|false|false|C0013227|Pharmaceutical Preparations|medication
Finding|Intellectual Product|History of Present Illness|950,960|true|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Anatomy|Body Location or Region|History of Present Illness|977,982|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|977,982|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|977,987|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|977,987|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|983,987|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|983,987|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|983,987|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|History of Present Illness|989,1001|false|false|false|C0030252|Palpitations|palpitations
Finding|Finding|History of Present Illness|1003,1015|false|false|false|C0030252|Palpitations|palpitations
Disorder|Disease or Syndrome|History of Present Illness|1028,1031|false|false|false|C1956415|Paroxysmal nocturnal dyspnea|PND
Finding|Gene or Genome|History of Present Illness|1028,1031|false|false|false|C1417807;C4552608|NPPA gene;NPPA wt Allele|PND
Finding|Daily or Recreational Activity|History of Present Illness|1043,1051|false|false|false|C0015259|Exercise|exercise
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1043,1051|false|false|false|C1522704|Exercise Pain Management|exercise
Attribute|Clinical Attribute|History of Present Illness|1043,1061|false|false|false|C0162521;C2709256|Exercise Tolerance|exercise tolerance
Finding|Finding|History of Present Illness|1043,1061|false|false|false|C2024889||exercise tolerance
Finding|Finding|History of Present Illness|1052,1061|false|false|false|C0013220;C0020963;C0220929;C0231197|Drug Tolerance;Immune Tolerance;Mental tolerance;Physiologic tolerance|tolerance
Finding|Mental Process|History of Present Illness|1052,1061|false|false|false|C0013220;C0020963;C0220929;C0231197|Drug Tolerance;Immune Tolerance;Mental tolerance;Physiologic tolerance|tolerance
Finding|Pathologic Function|History of Present Illness|1052,1061|false|false|false|C0013220;C0020963;C0220929;C0231197|Drug Tolerance;Immune Tolerance;Mental tolerance;Physiologic tolerance|tolerance
Finding|Physiologic Function|History of Present Illness|1052,1061|false|false|false|C0013220;C0020963;C0220929;C0231197|Drug Tolerance;Immune Tolerance;Mental tolerance;Physiologic tolerance|tolerance
Finding|Finding|History of Present Illness|1063,1069|false|false|false|C1299582|Unable|unable
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1082,1086|false|false|false|C0016504|Foot|feet
Finding|Finding|History of Present Illness|1093,1102|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Finding|Sign or Symptom|History of Present Illness|1093,1102|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Finding|Body Substance|History of Present Illness|1117,1124|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1117,1124|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1117,1124|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Anatomy|Body Location or Region|History of Present Illness|1156,1161|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|History of Present Illness|1156,1161|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1163,1172|false|false|false|C0015385|Limb structure|extremity
Finding|Pathologic Function|History of Present Illness|1163,1178|false|false|false|C0085649|Peripheral edema|extremity edema
Attribute|Clinical Attribute|History of Present Illness|1173,1178|false|false|false|C1717255||edema
Finding|Pathologic Function|History of Present Illness|1173,1178|false|false|false|C0013604|Edema|edema
Finding|Finding|History of Present Illness|1199,1207|false|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Finding|Functional Concept|History of Present Illness|1211,1215|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|History of Present Illness|1211,1215|false|false|false|C0582103|Medical Examination|exam
Finding|Body Substance|History of Present Illness|1217,1224|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|1217,1224|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|1217,1224|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Procedure|Diagnostic Procedure|History of Present Illness|1236,1239|false|false|false|C0039985|Plain chest X-ray|CXR
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1241,1244|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Hormone|History of Present Illness|1241,1244|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Pharmacologic Substance|History of Present Illness|1241,1244|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Finding|Gene or Genome|History of Present Illness|1241,1244|false|false|false|C1417808;C2982014|NPPB gene;NPPB wt Allele|BNP
Procedure|Laboratory Procedure|History of Present Illness|1241,1244|false|false|false|C1095989|Brain natriuretic peptide measurement|BNP
Drug|Organic Chemical|History of Present Illness|1280,1285|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|History of Present Illness|1280,1285|false|false|false|C0699992|Lasix|Lasix
Finding|Idea or Concept|History of Present Illness|1298,1305|false|false|false|C1555582|Initial (abbreviation)|initial
Finding|Functional Concept|History of Present Illness|1356,1364|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|History of Present Illness|1356,1364|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|History of Present Illness|1356,1364|false|false|false|C4706767|Transfer (immobility management)|transfer
Finding|Body Substance|History of Present Illness|1400,1407|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|1400,1407|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|1400,1407|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Lab|Laboratory or Test Result|History of Present Illness|1410,1414|false|false|false|C0587081|Laboratory test finding|labs
Drug|Biologically Active Substance|History of Present Illness|1436,1442|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|History of Present Illness|1436,1442|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|History of Present Illness|1436,1442|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Finding|Physiologic Function|History of Present Illness|1436,1442|false|false|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|History of Present Illness|1436,1442|false|false|false|C0337443|Sodium measurement|sodium
Drug|Element, Ion, or Isotope|History of Present Illness|1448,1456|false|false|false|C0008203;C0596019|Chlorides;chloride ion|Chloride
Finding|Physiologic Function|History of Present Illness|1448,1456|false|false|false|C4553021|Chloride metabolic function|Chloride
Procedure|Laboratory Procedure|History of Present Illness|1448,1456|false|false|false|C0201952|Chloride measurement|Chloride
Drug|Organic Chemical|History of Present Illness|1469,1475|false|false|false|C0074722|sodium bicarbonate|Bicarb
Drug|Pharmacologic Substance|History of Present Illness|1469,1475|false|false|false|C0074722|sodium bicarbonate|Bicarb
Drug|Biologically Active Substance|History of Present Illness|1480,1483|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Drug|Inorganic Chemical|History of Present Illness|1480,1483|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Procedure|Laboratory Procedure|History of Present Illness|1480,1483|false|false|false|C0005845|Blood urea nitrogen measurement|BUN
Drug|Biologically Active Substance|History of Present Illness|1489,1499|false|false|false|C0010294|creatinine|Creatinine
Drug|Organic Chemical|History of Present Illness|1489,1499|false|false|false|C0010294|creatinine|Creatinine
Finding|Physiologic Function|History of Present Illness|1489,1499|false|false|false|C4551889|Creatinine metabolic function|Creatinine
Procedure|Laboratory Procedure|History of Present Illness|1489,1499|false|false|false|C0201975|Creatinine measurement|Creatinine
Finding|Body Substance|History of Present Illness|1505,1512|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|1505,1512|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|1505,1512|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Body Substance|History of Present Illness|1550,1557|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|1550,1557|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|1550,1557|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1562,1565|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Hormone|History of Present Illness|1562,1565|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Pharmacologic Substance|History of Present Illness|1562,1565|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Finding|Gene or Genome|History of Present Illness|1562,1565|false|false|false|C1417808;C2982014|NPPB gene;NPPB wt Allele|BNP
Procedure|Laboratory Procedure|History of Present Illness|1562,1565|false|false|false|C1095989|Brain natriuretic peptide measurement|BNP
Finding|Body Substance|History of Present Illness|1577,1584|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|1577,1584|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|1577,1584|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1594,1597|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|History of Present Illness|1594,1597|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|History of Present Illness|1594,1597|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|History of Present Illness|1594,1597|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|History of Present Illness|1603,1606|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1603,1606|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Anatomy|Cell|History of Present Illness|1614,1622|false|false|false|C0005821|Blood Platelets|Platelet
Anatomy|Cell|History of Present Illness|1628,1631|false|false|false|C0023516|Leukocytes|WBC
Procedure|Laboratory Procedure|History of Present Illness|1637,1647|false|false|false|C0042014;C0373521|Urinalysis;Urinalysis; qualitative or semiquantitative, except immunoassays|Urinalysis
Disorder|Disease or Syndrome|History of Present Illness|1648,1653|false|false|false|C1410088|Still|still
Finding|Idea or Concept|History of Present Illness|1654,1661|false|false|false|C1691786;C1704475|Pending - Allergy Clinical Status;Pending - referral status|pending
Finding|Body Substance|History of Present Illness|1667,1676|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|History of Present Illness|1667,1676|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|History of Present Illness|1667,1676|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|History of Present Illness|1667,1676|false|false|false|C0030685|Patient Discharge|discharge
Finding|Intellectual Product|History of Present Illness|1680,1683|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|History of Present Illness|1680,1683|false|false|false|C1623258|Electrocardiography|EKG
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1709,1712|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|History of Present Illness|1709,1712|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|History of Present Illness|1709,1712|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Finding|Social Behavior|History of Present Illness|1725,1733|false|false|false|C0678975|inferiority|inferior
Finding|Finding|History of Present Illness|1755,1764|false|true|false|C0442739||unchanged
Anatomy|Anatomical Structure|History of Present Illness|1791,1796|false|false|false|C3714591|Floor (anatomic)|floor
Disorder|Disease or Syndrome|Past Medical History|1881,1893|false|false|false|C0020538|Hypertensive disease|hypertension
Disorder|Disease or Syndrome|Past Medical History|1898,1906|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|diabetes
Disorder|Disease or Syndrome|Past Medical History|1914,1917|false|false|false|C0001365;C0038454|Acute ill-defined cerebrovascular disease;Cerebrovascular accident|CVA
Drug|Pharmacologic Substance|Past Medical History|1914,1917|false|false|false|C5779650|Cyclophosphamide/Doxorubicin/Vincristine|CVA
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1919,1929|false|false|false|C0007765|Cerebellum|cerebellar
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1930,1939|false|false|false|C0001629;C0025148;C1550278|Adrenal Medulla;Medulla Oblongata;Medullary - body parts|medullary
Disorder|Disease or Syndrome|Past Medical History|1940,1946|false|false|false|C0038454|Cerebrovascular accident|stroke
Finding|Finding|Past Medical History|1940,1946|false|false|false|C5977286|Stroke (heart beat)|stroke
Disorder|Disease or Syndrome|Past Medical History|1958,1961|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Past Medical History|1958,1961|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Past Medical History|1958,1961|false|false|false|C1504769|DFFB protein, human|CAD
Finding|Gene or Genome|Past Medical History|1958,1961|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Past Medical History|1958,1961|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Past Medical History|1958,1961|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1958,1961|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|Past Medical History|1979,1982|false|false|false|C0006430|Burning Mouth Syndrome|BMS
Disorder|Disease or Syndrome|Past Medical History|2014,2041|false|false|false|C0085096;C1704436|Peripheral Arterial Diseases;Peripheral Vascular Diseases|peripheral arterial disease
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2025,2033|false|false|false|C0003842|Arteries|arterial
Disorder|Disease or Syndrome|Past Medical History|2025,2041|false|false|false|C0852949|Arteriopathic disease|arterial disease
Disorder|Disease or Syndrome|Past Medical History|2034,2041|false|false|false|C0012634|Disease|disease
Disorder|Disease or Syndrome|Past Medical History|2043,2055|false|true|false|C0021775|Intermittent Claudication|claudication
Finding|Finding|Past Medical History|2043,2055|false|true|false|C0311395;C1456822|Claudication (finding);Lameness|claudication
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2070,2078|false|false|false|C0005847|Blood Vessel|vascular
Attribute|Clinical Attribute|Past Medical History|2105,2110|false|false|false|C1300072|Tumor stage|stage
Finding|Intellectual Product|Past Medical History|2105,2113|false|false|false|C0441772|Stage level 4|stage IV
Disorder|Disease or Syndrome|Past Medical History|2114,2117|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Drug|Biomedical or Dental Material|Past Medical History|2119,2127|false|false|false|C0168634|BaseLine dental cement|baseline
Finding|Idea or Concept|Past Medical History|2119,2127|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Disorder|Disease or Syndrome|Past Medical History|2141,2145|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Disorder|Disease or Syndrome|Past Medical History|2146,2156|false|false|false|C0014852|Esophageal Diseases|esophageal
Disorder|Disease or Syndrome|Past Medical History|2146,2162|false|false|false|C0267081|Terminal esophageal web|esophageal rings
Finding|Conceptual Entity|Family Medical History|2201,2207|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|Family Medical History|2201,2207|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Anatomy|Body Location or Region|Family Medical History|2231,2235|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2231,2235|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Family Medical History|2231,2235|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Family Medical History|2231,2235|false|false|false|C0740941|Lung Problem|lung
Disorder|Disease or Syndrome|Family Medical History|2231,2243|false|false|false|C0024115|Lung diseases|lung disease
Disorder|Disease or Syndrome|Family Medical History|2236,2243|false|false|false|C0012634|Disease|disease
Finding|Idea or Concept|Family Medical History|2246,2252|false|false|false|C1546508|Relationship - Mother|Mother
Drug|Amino Acid, Peptide, or Protein|Family Medical History|2280,2287|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Immunologic Factor|Family Medical History|2280,2287|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Pharmacologic Substance|Family Medical History|2280,2287|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Finding|Finding|Family Medical History|2280,2287|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Functional Concept|Family Medical History|2280,2287|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Idea or Concept|Family Medical History|2280,2287|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Intellectual Product|Family Medical History|2280,2287|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Conceptual Entity|Family Medical History|2288,2293|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Finding|Functional Concept|Family Medical History|2288,2293|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Disorder|Disease or Syndrome|Family Medical History|2305,2308|true|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Family Medical History|2305,2308|true|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Family Medical History|2305,2308|true|false|false|C1504769|DFFB protein, human|CAD
Finding|Gene or Genome|Family Medical History|2305,2308|true|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Family Medical History|2305,2308|true|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Family Medical History|2305,2308|true|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2305,2308|true|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2319,2326|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|Family Medical History|2319,2326|true|false|false|C1314974|Cardiac attachment|cardiac
Finding|Finding|Family Medical History|2328,2333|false|false|false|C0011065;C1306577;C1546949|Cessation of life;Death (finding);Event Consequence - Death|death
Finding|Idea or Concept|Family Medical History|2328,2333|false|false|false|C0011065;C1306577;C1546949|Cessation of life;Death (finding);Event Consequence - Death|death
Finding|Organism Function|Family Medical History|2328,2333|false|false|false|C0011065;C1306577;C1546949|Cessation of life;Death (finding);Event Consequence - Death|death
Finding|Conceptual Entity|Family Medical History|2350,2357|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|2350,2357|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Family Medical History|2350,2357|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|2350,2360|false|false|false|C0262926|Medical History|history of
Finding|Finding|Family Medical History|2350,2367|true|false|false|C0455471|History of malignant neoplasm|history of cancer
Disorder|Neoplastic Process|Family Medical History|2361,2367|true|false|false|C0006826|Malignant Neoplasms|cancer
Procedure|Health Care Activity|General Exam|2386,2395|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Finding|Finding|General Exam|2396,2404|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|General Exam|2396,2404|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|General Exam|2396,2404|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|General Exam|2396,2416|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAMINATION
Procedure|Health Care Activity|General Exam|2396,2416|false|false|false|C0031809|Physical Examination|PHYSICAL EXAMINATION
Event|Activity|General Exam|2405,2416|false|false|false|C4321457|Examination|EXAMINATION
Procedure|Health Care Activity|General Exam|2405,2416|false|false|false|C0031809;C0582103|Medical Examination;Physical Examination|EXAMINATION
Procedure|Health Care Activity|General Exam|2477,2486|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|General Exam|2487,2493|false|false|false|C0944911||weight
Finding|Finding|General Exam|2487,2493|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|General Exam|2487,2493|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|General Exam|2487,2493|false|false|false|C1305866|Weighing patient|weight
Finding|Classification|General Exam|2501,2508|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|General Exam|2501,2508|false|false|false|C3812897|General medical service|GENERAL
Disorder|Disease or Syndrome|General Exam|2516,2521|false|false|false|C0028754|Obesity|obese
Finding|Finding|General Exam|2523,2538|false|false|false|C1280451|Sitting upright|sitting upright
Finding|Intellectual Product|General Exam|2531,2538|false|false|false|C1550127|Special Handling Code - Upright|upright
Phenomenon|Human-caused Phenomenon or Process|General Exam|2531,2538|false|false|false|C1550585|Entity Handling - upright|upright
Disorder|Disease or Syndrome|General Exam|2542,2545|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Finding|Intellectual Product|General Exam|2542,2545|false|false|false|C2346952|Bachelor of Education|bed
Disorder|Disease or Syndrome|General Exam|2550,2553|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|2550,2553|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|2550,2553|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|2550,2553|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|2550,2553|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Finding|Finding|General Exam|2550,2553|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Attribute|Clinical Attribute|General Exam|2562,2566|false|false|false|C2713234||Mood
Finding|Conceptual Entity|General Exam|2562,2566|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Finding|Finding|General Exam|2562,2566|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Finding|Mental Process|General Exam|2562,2566|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Anatomy|Body Location or Region|General Exam|2590,2595|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|General Exam|2603,2609|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|General Exam|2603,2609|false|false|false|C0036412|Scleral Diseases|Sclera
Procedure|Health Care Activity|General Exam|2603,2609|false|false|false|C2228481|examination of sclera|Sclera
Finding|Finding|General Exam|2610,2619|false|false|false|C0205180|Anicteric|anicteric
Finding|Finding|General Exam|2621,2626|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Anatomy|Body Part, Organ, or Organ Component|General Exam|2634,2645|false|false|false|C0009758;C0229274|Structure of palpebral conjunctiva;conjunctiva|Conjunctiva
Disorder|Disease or Syndrome|General Exam|2634,2645|false|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|Conjunctiva
Disorder|Neoplastic Process|General Exam|2634,2645|false|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|Conjunctiva
Finding|Body Substance|General Exam|2634,2645|false|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|Conjunctiva
Finding|Intellectual Product|General Exam|2634,2645|false|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|Conjunctiva
Procedure|Health Care Activity|General Exam|2634,2645|false|false|false|C0872390;C2228431|Procedure on conjunctiva;examination of conjunctiva|Conjunctiva
Finding|Finding|General Exam|2661,2667|true|false|false|C0241137|Pallor of skin|pallor
Finding|Sign or Symptom|General Exam|2671,2679|true|false|false|C0010520|Cyanosis|cyanosis
Anatomy|Body Space or Junction|General Exam|2687,2691|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|General Exam|2687,2691|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|General Exam|2687,2691|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|General Exam|2687,2691|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Anatomy|Body Part, Organ, or Organ Component|General Exam|2687,2698|false|false|false|C0026639|Oral mucous membrane structure|oral mucosa
Anatomy|Tissue|General Exam|2692,2698|false|false|false|C0026724|Mucous Membrane|mucosa
Finding|Intellectual Product|General Exam|2692,2698|false|false|false|C1561514||mucosa
Anatomy|Body Location or Region|General Exam|2700,2704|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|General Exam|2700,2704|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|General Exam|2700,2704|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Finding|Functional Concept|General Exam|2706,2712|false|false|false|C0332254|Supple|Supple
Finding|Finding|General Exam|2718,2721|false|false|false|C0428897|Jugular venous pressure|JVP
Anatomy|Body Part, Organ, or Organ Component|General Exam|2732,2739|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|General Exam|2732,2739|false|false|false|C1314974|Cardiac attachment|CARDIAC
Finding|Finding|General Exam|2741,2744|false|false|false|C1417244;C1418674;C1823304;C5238618;C5780972|MPI gene;PMM2 gene;PMM2 wt Allele;Point of Maximum Impulse;TMEM11 gene|PMI
Finding|Gene or Genome|General Exam|2741,2744|false|false|false|C1417244;C1418674;C1823304;C5238618;C5780972|MPI gene;PMM2 gene;PMM2 wt Allele;Point of Maximum Impulse;TMEM11 gene|PMI
Anatomy|Body Space or Junction|General Exam|2760,2777|false|false|false|C0230136;C4085247|Space of intercostal compartment;Structure of intercostal space|intercostal space
Phenomenon|Natural Phenomenon or Process|General Exam|2772,2777|false|false|false|C0282173|Space (Astronomy)|space
Drug|Biologically Active Substance|General Exam|2794,2798|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|2794,2798|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Substance|General Exam|2794,2798|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Finding|Intellectual Product|General Exam|2794,2798|false|false|false|C1546701|line source specimen code|line
Finding|Finding|General Exam|2827,2834|true|false|false|C0018808|Heart murmur|murmurs
Finding|Finding|General Exam|2835,2839|true|false|false|C0232267|Pericardial friction rub|rubs
Finding|Finding|General Exam|2853,2860|false|false|false|C0232269|Cardiac thrill (finding)|thrills
Anatomy|Body Part, Organ, or Organ Component|General Exam|2870,2875|false|false|false|C0024109|Lung|LUNGS
Attribute|Clinical Attribute|General Exam|2877,2881|false|false|false|C0231832|Respiratory rate|Resp
Disorder|Disease or Syndrome|General Exam|2877,2881|false|false|false|C0851355|Respiratory, thoracic and mediastinal disorders|Resp
Finding|Functional Concept|General Exam|2887,2896|false|false|false|C2983702|Unlabored|unlabored
Disorder|Congenital Abnormality|General Exam|2901,2917|true|false|false|C0158784|Accessory skeletal muscle|accessory muscle
Finding|Finding|General Exam|2901,2921|true|false|false|C1821466|Use of accessory muscles|accessory muscle use
Anatomy|Body Part, Organ, or Organ Component|General Exam|2911,2917|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|General Exam|2911,2917|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Finding|Functional Concept|General Exam|2918,2921|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|General Exam|2918,2921|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Finding|General Exam|2923,2931|false|false|false|C0277854|dyspneic|dyspneic
Drug|Amino Acid, Peptide, or Protein|General Exam|2940,2943|false|false|false|C0082420|Endoglin, human|end
Drug|Immunologic Factor|General Exam|2940,2943|false|false|false|C0082420|Endoglin, human|end
Finding|Functional Concept|General Exam|2940,2943|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Finding|Gene or Genome|General Exam|2940,2943|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Finding|Intellectual Product|General Exam|2954,2962|false|false|false|C0876929|Sentence|sentence
Finding|Finding|General Exam|2974,2982|false|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Anatomy|Body Location or Region|General Exam|2990,2996|false|false|false|C0817096|Chest|thorax
Disorder|Neoplastic Process|General Exam|2990,2996|false|false|false|C0153661|Malignant neoplasm of thorax|thorax
Finding|Finding|General Exam|2999,3015|false|false|false|C2089439|diffuse wheezing|diffuse wheezing
Finding|Sign or Symptom|General Exam|3007,3015|false|false|false|C0043144|Wheezing|wheezing
Anatomy|Body Location or Region|General Exam|3019,3026|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|General Exam|3019,3026|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Finding|Finding|General Exam|3019,3026|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|General Exam|3028,3032|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Finding|Gene or Genome|General Exam|3043,3046|true|false|false|C1537594|LRRC4B gene|HSM
Finding|Mental Process|General Exam|3050,3060|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|General Exam|3050,3060|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Anatomy|Body Part, Organ, or Organ Component|General Exam|3064,3075|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Attribute|Clinical Attribute|General Exam|3080,3085|false|false|false|C1717255||edema
Finding|Pathologic Function|General Exam|3080,3085|false|false|false|C0013604|Edema|edema
Anatomy|Body Location or Region|General Exam|3089,3094|false|false|false|C0230444|Shin|shins
Anatomy|Body Part, Organ, or Organ Component|General Exam|3099,3106|false|false|false|C0015811|Femur|femoral
Finding|Finding|General Exam|3107,3113|true|false|false|C0006318|Bruit|bruits
Drug|Food|General Exam|3117,3123|false|false|false|C5890763||PULSES
Finding|Physiologic Function|General Exam|3117,3123|false|false|false|C0391850|Physiologic pulse|PULSES
Procedure|Health Care Activity|General Exam|3117,3123|false|false|false|C0034107|Pulse taking|PULSES
Attribute|Clinical Attribute|General Exam|3126,3132|false|false|false|C4522154|Distal Resection Margin|Distal
Drug|Food|General Exam|3133,3139|false|false|false|C5890763||pulses
Finding|Physiologic Function|General Exam|3133,3139|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|3133,3139|false|false|false|C0034107|Pulse taking|pulses
Finding|Conceptual Entity|General Exam|3153,3162|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|General Exam|3153,3162|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Body Substance|General Exam|3164,3173|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|3164,3173|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|3164,3173|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|3164,3173|false|false|false|C0030685|Patient Discharge|DISCHARGE
Finding|Finding|General Exam|3174,3182|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|General Exam|3174,3182|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|General Exam|3174,3182|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|General Exam|3174,3194|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAMINATION
Procedure|Health Care Activity|General Exam|3174,3194|false|false|false|C0031809|Physical Examination|PHYSICAL EXAMINATION
Event|Activity|General Exam|3183,3194|false|false|false|C4321457|Examination|EXAMINATION
Procedure|Health Care Activity|General Exam|3183,3194|false|false|false|C0031809;C0582103|Medical Examination;Physical Examination|EXAMINATION
Attribute|Clinical Attribute|General Exam|3250,3256|false|false|false|C0944911||weight
Finding|Finding|General Exam|3250,3256|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|General Exam|3250,3256|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|General Exam|3250,3256|false|false|false|C1305866|Weighing patient|weight
Finding|Classification|General Exam|3263,3270|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|General Exam|3263,3270|false|false|false|C3812897|General medical service|GENERAL
Disorder|Disease or Syndrome|General Exam|3278,3283|false|false|false|C0028754|Obesity|obese
Finding|Finding|General Exam|3285,3300|false|false|false|C1280451|Sitting upright|sitting upright
Finding|Intellectual Product|General Exam|3293,3300|false|false|false|C1550127|Special Handling Code - Upright|upright
Phenomenon|Human-caused Phenomenon or Process|General Exam|3293,3300|false|false|false|C1550585|Entity Handling - upright|upright
Disorder|Disease or Syndrome|General Exam|3304,3307|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Finding|Intellectual Product|General Exam|3304,3307|false|false|false|C2346952|Bachelor of Education|bed
Disorder|Disease or Syndrome|General Exam|3312,3315|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|3312,3315|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|3312,3315|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|3312,3315|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|3312,3315|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Finding|Finding|General Exam|3312,3315|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Attribute|Clinical Attribute|General Exam|3324,3328|false|false|false|C2713234||Mood
Finding|Conceptual Entity|General Exam|3324,3328|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Finding|Finding|General Exam|3324,3328|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Finding|Mental Process|General Exam|3324,3328|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Anatomy|Body Location or Region|General Exam|3352,3357|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|General Exam|3365,3371|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|General Exam|3365,3371|false|false|false|C0036412|Scleral Diseases|Sclera
Procedure|Health Care Activity|General Exam|3365,3371|false|false|false|C2228481|examination of sclera|Sclera
Finding|Finding|General Exam|3372,3381|false|false|false|C0205180|Anicteric|anicteric
Finding|Finding|General Exam|3383,3388|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Anatomy|Body Part, Organ, or Organ Component|General Exam|3396,3407|false|false|false|C0009758;C0229274|Structure of palpebral conjunctiva;conjunctiva|Conjunctiva
Disorder|Disease or Syndrome|General Exam|3396,3407|false|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|Conjunctiva
Disorder|Neoplastic Process|General Exam|3396,3407|false|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|Conjunctiva
Finding|Body Substance|General Exam|3396,3407|false|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|Conjunctiva
Finding|Intellectual Product|General Exam|3396,3407|false|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|Conjunctiva
Procedure|Health Care Activity|General Exam|3396,3407|false|false|false|C0872390;C2228431|Procedure on conjunctiva;examination of conjunctiva|Conjunctiva
Finding|Finding|General Exam|3423,3429|true|false|false|C0241137|Pallor of skin|pallor
Finding|Sign or Symptom|General Exam|3433,3441|true|false|false|C0010520|Cyanosis|cyanosis
Anatomy|Body Space or Junction|General Exam|3449,3453|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|General Exam|3449,3453|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|General Exam|3449,3453|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|General Exam|3449,3453|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Anatomy|Body Part, Organ, or Organ Component|General Exam|3449,3460|false|false|false|C0026639|Oral mucous membrane structure|oral mucosa
Anatomy|Tissue|General Exam|3454,3460|false|false|false|C0026724|Mucous Membrane|mucosa
Finding|Intellectual Product|General Exam|3454,3460|false|false|false|C1561514||mucosa
Anatomy|Body Location or Region|General Exam|3462,3466|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|General Exam|3462,3466|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|General Exam|3462,3466|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Finding|Functional Concept|General Exam|3468,3474|false|false|false|C0332254|Supple|Supple
Finding|Finding|General Exam|3480,3483|false|false|false|C0428897|Jugular venous pressure|JVP
Anatomy|Body Part, Organ, or Organ Component|General Exam|3494,3501|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|General Exam|3494,3501|false|false|false|C1314974|Cardiac attachment|CARDIAC
Finding|Finding|General Exam|3503,3506|false|false|false|C1417244;C1418674;C1823304;C5238618;C5780972|MPI gene;PMM2 gene;PMM2 wt Allele;Point of Maximum Impulse;TMEM11 gene|PMI
Finding|Gene or Genome|General Exam|3503,3506|false|false|false|C1417244;C1418674;C1823304;C5238618;C5780972|MPI gene;PMM2 gene;PMM2 wt Allele;Point of Maximum Impulse;TMEM11 gene|PMI
Anatomy|Body Space or Junction|General Exam|3522,3539|false|false|false|C0230136;C4085247|Space of intercostal compartment;Structure of intercostal space|intercostal space
Phenomenon|Natural Phenomenon or Process|General Exam|3534,3539|false|false|false|C0282173|Space (Astronomy)|space
Drug|Biologically Active Substance|General Exam|3556,3560|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|3556,3560|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Substance|General Exam|3556,3560|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Finding|Intellectual Product|General Exam|3556,3560|false|false|false|C1546701|line source specimen code|line
Finding|Finding|General Exam|3589,3596|true|false|false|C0018808|Heart murmur|murmurs
Finding|Finding|General Exam|3597,3601|true|false|false|C0232267|Pericardial friction rub|rubs
Finding|Finding|General Exam|3615,3622|false|false|false|C0232269|Cardiac thrill (finding)|thrills
Anatomy|Body Part, Organ, or Organ Component|General Exam|3632,3637|false|false|false|C0024109|Lung|LUNGS
Attribute|Clinical Attribute|General Exam|3639,3643|false|false|false|C0231832|Respiratory rate|Resp
Disorder|Disease or Syndrome|General Exam|3639,3643|false|false|false|C0851355|Respiratory, thoracic and mediastinal disorders|Resp
Finding|Functional Concept|General Exam|3649,3658|false|false|false|C2983702|Unlabored|unlabored
Disorder|Congenital Abnormality|General Exam|3663,3679|true|false|false|C0158784|Accessory skeletal muscle|accessory muscle
Finding|Finding|General Exam|3663,3683|true|false|false|C1821466|Use of accessory muscles|accessory muscle use
Anatomy|Body Part, Organ, or Organ Component|General Exam|3673,3679|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|General Exam|3673,3679|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Finding|Functional Concept|General Exam|3680,3683|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|General Exam|3680,3683|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Finding|General Exam|3696,3704|false|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Finding|Functional Concept|General Exam|3705,3710|false|false|false|C1883002|Sequence Chromatogram|trace
Finding|Finding|General Exam|3712,3728|false|false|false|C2089439|diffuse wheezing|diffuse wheezing
Finding|Sign or Symptom|General Exam|3720,3728|false|false|false|C0043144|Wheezing|wheezing
Anatomy|Body Location or Region|General Exam|3732,3739|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|General Exam|3732,3739|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Finding|Finding|General Exam|3732,3739|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|General Exam|3741,3745|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Finding|Gene or Genome|General Exam|3756,3759|true|false|false|C1537594|LRRC4B gene|HSM
Finding|Mental Process|General Exam|3763,3773|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|General Exam|3763,3773|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Anatomy|Body Part, Organ, or Organ Component|General Exam|3777,3788|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Anatomy|Body Part, Organ, or Organ Component|General Exam|3798,3805|false|false|false|C0015811|Femur|femoral
Finding|Finding|General Exam|3806,3812|true|false|false|C0006318|Bruit|bruits
Drug|Food|General Exam|3816,3822|false|false|false|C5890763||PULSES
Finding|Physiologic Function|General Exam|3816,3822|false|false|false|C0391850|Physiologic pulse|PULSES
Procedure|Health Care Activity|General Exam|3816,3822|false|false|false|C0034107|Pulse taking|PULSES
Attribute|Clinical Attribute|General Exam|3825,3831|false|false|false|C4522154|Distal Resection Margin|Distal
Drug|Food|General Exam|3832,3838|false|false|false|C5890763||pulses
Finding|Physiologic Function|General Exam|3832,3838|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|3832,3838|false|false|false|C0034107|Pulse taking|pulses
Finding|Conceptual Entity|General Exam|3852,3861|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|General Exam|3852,3861|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Procedure|Health Care Activity|General Exam|3883,3892|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Lab|Laboratory or Test Result|General Exam|3893,3897|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|General Exam|3910,3915|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3910,3915|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|3916,3919|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|3924,3927|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|3924,3927|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|3924,3927|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|3934,3937|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|3934,3937|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|3934,3937|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|3934,3937|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|3943,3946|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|3943,3946|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|3954,3957|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|General Exam|3954,3957|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|3954,3957|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|3954,3957|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|3964,3967|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|3964,3967|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|General Exam|3964,3967|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|3964,3967|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|3964,3967|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|3973,3977|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|4006,4009|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|4026,4031|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4026,4031|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Body Substance|General Exam|4044,4050|false|false|false|C0024202|Lymph|Lymphs
Drug|Antibiotic|General Exam|4057,4062|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|General Exam|4057,4062|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|General Exam|4057,4062|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|General Exam|4068,4071|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Finding|Gene or Genome|General Exam|4068,4071|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|General Exam|4170,4175|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4170,4175|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|4180,4183|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Procedure|Laboratory Procedure|General Exam|4180,4183|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|General Exam|4205,4210|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4205,4210|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|4211,4214|false|false|false|C0389252|RET protein, human|Ret
Finding|Gene or Genome|General Exam|4211,4214|false|false|false|C0389252;C0694890;C0813143;C1704885|Oncogene RET;RET gene;RET protein, human;RET wt Allele|Ret
Finding|Receptor|General Exam|4211,4214|false|false|false|C0389252;C0694890;C0813143;C1704885|Oncogene RET;RET gene;RET protein, human;RET wt Allele|Ret
Disorder|Congenital Abnormality|General Exam|4224,4227|false|false|false|C0002636;C0220724|Amniotic Band Syndrome;CONSTRICTING BANDS, CONGENITAL|Abs
Disorder|Disease or Syndrome|General Exam|4224,4227|false|false|false|C0002636;C0220724|Amniotic Band Syndrome;CONSTRICTING BANDS, CONGENITAL|Abs
Finding|Gene or Genome|General Exam|4224,4227|false|false|false|C1425698;C4723885|DDX41 gene;DDX41 wt Allele|Abs
Drug|Amino Acid, Peptide, or Protein|General Exam|4228,4231|false|false|false|C0389252|RET protein, human|Ret
Finding|Gene or Genome|General Exam|4228,4231|false|false|false|C0389252;C0694890;C0813143;C1704885|Oncogene RET;RET gene;RET protein, human;RET wt Allele|Ret
Finding|Receptor|General Exam|4228,4231|false|false|false|C0389252;C0694890;C0813143;C1704885|Oncogene RET;RET gene;RET protein, human;RET wt Allele|Ret
Disorder|Disease or Syndrome|General Exam|4249,4254|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4249,4254|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|4249,4262|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|4249,4262|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|4249,4262|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|4255,4262|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|4255,4262|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|4255,4262|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|General Exam|4255,4262|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|4255,4262|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|4313,4317|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|4313,4317|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|4313,4317|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|4343,4348|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4343,4348|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|4349,4354|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|General Exam|4349,4354|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|General Exam|4349,4354|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|General Exam|4349,4354|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Drug|Pharmacologic Substance|General Exam|4352,4356|false|false|false|C4722362|MB-6|MB-6
Disorder|Disease or Syndrome|General Exam|4387,4392|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4387,4392|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|4393,4398|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|General Exam|4393,4398|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|General Exam|4393,4398|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|General Exam|4393,4398|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Drug|Pharmacologic Substance|General Exam|4396,4400|false|false|false|C4722362|MB-6|MB-6
Disorder|Disease or Syndrome|General Exam|4427,4432|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4427,4432|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|4427,4440|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|General Exam|4433,4440|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|4433,4440|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|4433,4440|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|4433,4440|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|4433,4440|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Finding|Physiologic Function|General Exam|4433,4440|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|4433,4440|false|false|false|C0201925|Calcium measurement|Calcium
Finding|Body Substance|General Exam|4462,4471|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|4462,4471|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|4462,4471|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|4462,4471|false|false|false|C0030685|Patient Discharge|DISCHARGE
Lab|Laboratory or Test Result|General Exam|4472,4476|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|General Exam|4495,4500|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4495,4500|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|4501,4504|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|4510,4513|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|4510,4513|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|4510,4513|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|4520,4523|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|4520,4523|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|4520,4523|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|4520,4523|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|4529,4532|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|4529,4532|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|4540,4543|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|General Exam|4540,4543|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|4540,4543|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|4540,4543|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|4547,4550|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|4547,4550|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|General Exam|4547,4550|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|4547,4550|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|4547,4550|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|4556,4560|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|4588,4591|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|4608,4613|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4608,4613|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|General Exam|4630,4635|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4630,4635|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|4630,4643|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|4630,4643|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|4630,4643|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|4636,4643|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|4636,4643|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|4636,4643|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|General Exam|4636,4643|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|4636,4643|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|4690,4694|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|4690,4694|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|4690,4694|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|4719,4724|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4719,4724|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|4719,4732|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|General Exam|4725,4732|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|4725,4732|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|4725,4732|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|4725,4732|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|4725,4732|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Finding|Physiologic Function|General Exam|4725,4732|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|4725,4732|false|false|false|C0201925|Calcium measurement|Calcium
Finding|Finding|General Exam|4754,4761|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|General Exam|4754,4761|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Procedure|Diagnostic Procedure|General Exam|4772,4775|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Intellectual Product|Findings|4796,4800|false|false|false|C1547225|Mild Severity of Illness Code|mild
Anatomy|Body Part, Organ, or Organ Component|Findings|4801,4810|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Findings|4801,4810|false|false|false|C2707265||pulmonary
Finding|Finding|Findings|4801,4810|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|Findings|4801,4816|false|false|false|C0034063|Pulmonary Edema|pulmonary edema
Attribute|Clinical Attribute|Findings|4811,4816|false|false|false|C1717255||edema
Finding|Pathologic Function|Findings|4811,4816|false|false|false|C0013604|Edema|edema
Drug|Amino Acid Sequence|Findings|4835,4841|false|false|false|C1514562|Protein Domain|region
Disorder|Disease or Syndrome|Findings|4861,4874|false|false|false|C0521530|Lung consolidation|consolidation
Finding|Functional Concept|Findings|4882,4886|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|Findings|4893,4897|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Findings|4893,4897|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Findings|4893,4897|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Findings|4893,4897|false|false|false|C0740941|Lung Problem|lung
Finding|Finding|Findings|4911,4919|false|false|false|C0332149|Possible|possible
Anatomy|Tissue|Findings|4936,4943|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|Findings|4936,4943|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Pathologic Function|Findings|4936,4953|false|false|false|C0032227|Pleural effusion (disorder)|pleural effusions
Finding|Pathologic Function|Findings|4944,4953|false|false|false|C0013687|effusion|effusions
Finding|Finding|Findings|4956,4964|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|Findings|4956,4964|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Finding|Findings|4966,4978|false|false|false|C0018800|Cardiomegaly|cardiomegaly
Finding|Finding|Findings|4996,5000|false|false|false|C5575035|Well (answer to question)|well
Finding|Functional Concept|Findings|5023,5033|false|false|false|C1547177|Sequencing - Descending|descending
Anatomy|Body Part, Organ, or Organ Component|Findings|5023,5048|false|false|false|C1522460;C3163626|Descending thoracic aorta;Thoracic aorta|descending thoracic aorta
Anatomy|Body Location or Region|Findings|5034,5042|false|false|false|C0817096|Chest|thoracic
Disorder|Disease or Syndrome|Findings|5034,5042|false|false|false|C5779551|Dissecting Thoracic Aortic Aneurysm|thoracic
Anatomy|Body Part, Organ, or Organ Component|Findings|5034,5048|false|false|false|C1522460;C4037977|Chest>Aorta.thoracic;Thoracic aorta|thoracic aorta
Anatomy|Body Part, Organ, or Organ Component|Findings|5043,5048|false|false|false|C0003483;C4037978|Aorta;Chest+Abdomen>Aorta|aorta
Procedure|Health Care Activity|Findings|5043,5048|false|false|false|C0869784|Procedure on aorta|aorta
Finding|Intellectual Product|Findings|5054,5059|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Part, Organ, or Organ Component|Findings|5060,5067|false|false|false|C0262950;C4520924|Bone Tissue, Human;Skeletal bone|osseous
Anatomy|Tissue|Findings|5060,5067|false|false|false|C0262950;C4520924|Bone Tissue, Human;Skeletal bone|osseous
Disorder|Congenital Abnormality|Findings|5068,5081|true|false|false|C0000768|Congenital Abnormality|abnormalities
Finding|Functional Concept|Findings|5068,5081|true|false|false|C0000769|teratologic|abnormalities
Finding|Intellectual Product|Impression|5098,5102|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Anatomy|Body Part, Organ, or Organ Component|Impression|5103,5112|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Impression|5103,5112|false|false|false|C2707265||pulmonary
Finding|Finding|Impression|5103,5112|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|Impression|5103,5118|false|false|false|C0034063|Pulmonary Edema|pulmonary edema
Attribute|Clinical Attribute|Impression|5113,5118|false|false|false|C1717255||edema
Finding|Pathologic Function|Impression|5113,5118|false|false|false|C0013604|Edema|edema
Finding|Functional Concept|Impression|5137,5141|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|Impression|5148,5152|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Impression|5148,5152|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Impression|5148,5152|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Impression|5148,5152|false|false|false|C0740941|Lung Problem|lung
Disorder|Disease or Syndrome|Impression|5154,5167|false|false|false|C0521530|Lung consolidation|consolidation
Attribute|Clinical Attribute|Impression|5196,5201|false|false|false|C1717255||edema
Finding|Pathologic Function|Impression|5196,5201|false|false|false|C0013604|Edema|edema
Disorder|Disease or Syndrome|Impression|5223,5232|false|false|false|C0009450|Communicable Diseases|infection
Finding|Pathologic Function|Impression|5223,5232|false|false|false|C3714514|Infection|infection
Finding|Idea or Concept|Hospital Course|5264,5268|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|Hospital Course|5264,5268|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Conceptual Entity|Hospital Course|5285,5292|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|5285,5292|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|5285,5292|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|5285,5295|false|false|false|C0262926|Medical History|history of
Finding|Finding|Hospital Course|5285,5308|false|false|false|C0455527||history of hypertension
Disorder|Disease or Syndrome|Hospital Course|5296,5308|false|false|false|C0020538|Hypertensive disease|hypertension
Disorder|Disease or Syndrome|Hospital Course|5310,5313|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5310,5313|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|5310,5313|false|false|false|C1504769|DFFB protein, human|CAD
Finding|Gene or Genome|Hospital Course|5310,5313|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|5310,5313|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|5310,5313|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5310,5313|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|Hospital Course|5318,5321|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5318,5321|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|Hospital Course|5318,5321|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|Hospital Course|5318,5321|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|Hospital Course|5318,5321|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|Hospital Course|5318,5321|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Finding|Gene or Genome|Hospital Course|5318,5321|false|false|false|C1413980|DES gene|DES
Finding|Functional Concept|Hospital Course|5328,5336|false|false|false|C0475224|Ischemic|ischemic
Finding|Organ or Tissue Function|Hospital Course|5344,5352|false|false|false|C0039155|Systole|systolic
Finding|Pathologic Function|Hospital Course|5344,5364|false|false|false|C0749225|Systolic dysfunction|systolic dysfunction
Disorder|Disease or Syndrome|Hospital Course|5353,5364|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Finding|Conceptual Entity|Hospital Course|5353,5364|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|Hospital Course|5353,5364|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|Hospital Course|5353,5364|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Anatomy|Body Location or Region|Hospital Course|5377,5380|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Hospital Course|5377,5380|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Hospital Course|5377,5380|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Anatomy|Body Space or Junction|Hospital Course|5400,5403|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|Hospital Course|5400,5403|false|false|false|C0018802|Congestive heart failure|CHF
Finding|Finding|Hospital Course|5404,5416|false|false|false|C4086268|Exacerbation|exacerbation
Finding|Intellectual Product|Hospital Course|5421,5426|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Finding|Intellectual Product|Hospital Course|5430,5437|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Hospital Course|5430,5437|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|Hospital Course|5438,5465|false|false|false|C0581377|Decompensated cardiac failure|decompensated heart failure
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5452,5457|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Hospital Course|5452,5457|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Hospital Course|5452,5457|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|Hospital Course|5452,5465|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Finding|Functional Concept|Hospital Course|5458,5465|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|Hospital Course|5458,5465|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|Hospital Course|5458,5465|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Mental Process|Hospital Course|5485,5492|false|false|false|C0542559|contextual factors|setting
Finding|Finding|Hospital Course|5496,5500|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|Hospital Course|5496,5500|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|Hospital Course|5496,5500|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Drug|Chemical Viewed Structurally|Hospital Course|5501,5505|false|false|false|C0036140;C0037494;C0206136|Salts;Sodium Chloride, Dietary;sodium chloride|salt
Drug|Food|Hospital Course|5501,5505|false|false|false|C0036140;C0037494;C0206136|Salts;Sodium Chloride, Dietary;sodium chloride|salt
Drug|Inorganic Chemical|Hospital Course|5501,5505|false|false|false|C0036140;C0037494;C0206136|Salts;Sodium Chloride, Dietary;sodium chloride|salt
Drug|Food|Hospital Course|5506,5510|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Finding|Functional Concept|Hospital Course|5506,5510|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|Hospital Course|5506,5510|false|false|false|C0012159|Diet therapy|diet
Finding|Finding|Hospital Course|5516,5523|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|Hospital Course|5516,5523|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|Hospital Course|5516,5535|false|false|false|C0231807|Dyspnea on exertion|dyspnea on exertion
Finding|Organism Function|Hospital Course|5527,5535|false|false|false|C0015264|Exertion|exertion
Finding|Daily or Recreational Activity|Hospital Course|5548,5556|false|false|false|C0015259|Exercise|exercise
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5548,5556|false|false|false|C1522704|Exercise Pain Management|exercise
Attribute|Clinical Attribute|Hospital Course|5548,5566|false|false|false|C0162521;C2709256|Exercise Tolerance|exercise tolerance
Finding|Finding|Hospital Course|5548,5566|false|false|false|C2024889||exercise tolerance
Finding|Finding|Hospital Course|5557,5566|false|false|false|C0013220;C0020963;C0220929;C0231197|Drug Tolerance;Immune Tolerance;Mental tolerance;Physiologic tolerance|tolerance
Finding|Mental Process|Hospital Course|5557,5566|false|false|false|C0013220;C0020963;C0220929;C0231197|Drug Tolerance;Immune Tolerance;Mental tolerance;Physiologic tolerance|tolerance
Finding|Pathologic Function|Hospital Course|5557,5566|false|false|false|C0013220;C0020963;C0220929;C0231197|Drug Tolerance;Immune Tolerance;Mental tolerance;Physiologic tolerance|tolerance
Finding|Physiologic Function|Hospital Course|5557,5566|false|false|false|C0013220;C0020963;C0220929;C0231197|Drug Tolerance;Immune Tolerance;Mental tolerance;Physiologic tolerance|tolerance
Attribute|Clinical Attribute|Hospital Course|5572,5577|false|false|false|C1717255||edema
Finding|Pathologic Function|Hospital Course|5572,5577|false|false|false|C0013604|Edema|edema
Finding|Finding|Hospital Course|5579,5587|false|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Finding|Functional Concept|Hospital Course|5591,5595|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|Hospital Course|5591,5595|false|false|false|C0582103|Medical Examination|exam
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5606,5609|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Hormone|Hospital Course|5606,5609|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Pharmacologic Substance|Hospital Course|5606,5609|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Finding|Gene or Genome|Hospital Course|5606,5609|false|false|false|C1417808;C2982014|NPPB gene;NPPB wt Allele|BNP
Procedure|Laboratory Procedure|Hospital Course|5606,5609|false|false|false|C1095989|Brain natriuretic peptide measurement|BNP
Attribute|Clinical Attribute|Hospital Course|5634,5640|false|false|false|C0944911||weight
Finding|Finding|Hospital Course|5634,5640|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|Hospital Course|5634,5640|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|Hospital Course|5634,5640|false|false|false|C1305866|Weighing patient|weight
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5645,5654|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Hospital Course|5645,5654|false|false|false|C2707265||pulmonary
Finding|Finding|Hospital Course|5645,5654|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Disorder|Disease or Syndrome|Hospital Course|5645,5665|false|false|false|C0242073|Pulmonary congestion|pulmonary congestion
Finding|Pathologic Function|Hospital Course|5655,5665|false|false|false|C0700148|Congestion|congestion
Procedure|Diagnostic Procedure|Hospital Course|5669,5672|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Intellectual Product|Hospital Course|5695,5703|false|false|false|C1547997;C3244303|Diagnostic Service Section ID - Pharmacy;Pharmacy domain|pharmacy
Procedure|Health Care Activity|Hospital Course|5695,5703|false|false|false|C0031321|Pharmaceutical Services|pharmacy
Finding|Idea or Concept|Hospital Course|5704,5710|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Intellectual Product|Hospital Course|5704,5710|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Body Substance|Hospital Course|5716,5723|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|5716,5723|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|5716,5723|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Organic Chemical|Hospital Course|5740,5749|false|false|false|C0076840|torsemide|torsemide
Drug|Pharmacologic Substance|Hospital Course|5740,5749|false|false|false|C0076840|torsemide|torsemide
Finding|Classification|Hospital Course|5761,5771|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|5761,5771|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Anatomy|Body System|Hospital Course|5772,5782|false|false|false|C0007226|Cardiovascular system|Cardiology
Event|Activity|Hospital Course|5783,5794|false|false|false|C0003629|Appointments|appointment
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5841,5850|false|false|false|C0041199|Troponin|Troponins
Drug|Biologically Active Substance|Hospital Course|5841,5850|false|false|false|C0041199|Troponin|Troponins
Finding|Classification|Hospital Course|5863,5871|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|5863,5871|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|5863,5871|false|false|false|C5237010|Expression Negative|negative
Procedure|Health Care Activity|Hospital Course|5876,5885|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Drug|Chemical Viewed Structurally|Hospital Course|5907,5911|false|false|false|C0036140;C0037494;C0206136|Salts;Sodium Chloride, Dietary;sodium chloride|salt
Drug|Food|Hospital Course|5907,5911|false|false|false|C0036140;C0037494;C0206136|Salts;Sodium Chloride, Dietary;sodium chloride|salt
Drug|Inorganic Chemical|Hospital Course|5907,5911|false|false|false|C0036140;C0037494;C0206136|Salts;Sodium Chloride, Dietary;sodium chloride|salt
Drug|Substance|Hospital Course|5916,5921|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|5916,5921|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Functional Concept|Hospital Course|5923,5933|false|false|false|C0443288;C1548390;C1549594;C1610594|Confidentiality - restricted;Confidentiality code - Restricted;Document Confidentiality Status - Restricted;Restricted|restricted
Finding|Idea or Concept|Hospital Course|5923,5933|false|false|false|C0443288;C1548390;C1549594;C1610594|Confidentiality - restricted;Confidentiality code - Restricted;Document Confidentiality Status - Restricted;Restricted|restricted
Finding|Intellectual Product|Hospital Course|5923,5933|false|false|false|C0443288;C1548390;C1549594;C1610594|Confidentiality - restricted;Confidentiality code - Restricted;Document Confidentiality Status - Restricted;Restricted|restricted
Procedure|Health Care Activity|Hospital Course|5923,5938|false|false|false|C0425422|Dietary Restriction|restricted diet
Drug|Food|Hospital Course|5934,5938|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Finding|Functional Concept|Hospital Course|5934,5938|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|Hospital Course|5934,5938|false|false|false|C0012159|Diet therapy|diet
Drug|Organic Chemical|Hospital Course|5965,5970|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|Hospital Course|5965,5970|false|false|false|C0699992|Lasix|Lasix
Finding|Intellectual Product|Hospital Course|5992,5996|false|false|false|C1720594|Then - dosing instruction fragment|then
Drug|Organic Chemical|Hospital Course|6016,6025|false|false|false|C0076840|torsemide|torsemide
Drug|Pharmacologic Substance|Hospital Course|6016,6025|false|false|false|C0076840|torsemide|torsemide
Attribute|Clinical Attribute|Hospital Course|6043,6049|false|false|false|C0944911||weight
Finding|Finding|Hospital Course|6043,6049|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|Hospital Course|6043,6049|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|Hospital Course|6043,6049|false|false|false|C1305866|Weighing patient|weight
Anatomy|Cell Component|Hospital Course|6063,6066|false|false|false|C3850088|Neutrophil Extracellular Traps|net
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6063,6066|false|false|false|C1456447;C3853572|Ephrin Type-B Receptor 1, human;SLC6A2 protein, human|net
Drug|Biologically Active Substance|Hospital Course|6063,6066|false|false|false|C1456447;C3853572|Ephrin Type-B Receptor 1, human;SLC6A2 protein, human|net
Drug|Enzyme|Hospital Course|6063,6066|false|false|false|C1456447;C3853572|Ephrin Type-B Receptor 1, human;SLC6A2 protein, human|net
Finding|Gene or Genome|Hospital Course|6063,6066|false|false|false|C0812375;C0815327;C1366441;C1420212;C1704819;C1705456;C3853572;C3890893|ELK3 gene;ELK3 wt Allele;EPHB1 gene;EPHB1 wt Allele;Ephrin Type-B Receptor 1, human;NET questionnaire;SLC6A2 gene;SLC6A2 wt Allele|net
Finding|Intellectual Product|Hospital Course|6063,6066|false|false|false|C0812375;C0815327;C1366441;C1420212;C1704819;C1705456;C3853572;C3890893|ELK3 gene;ELK3 wt Allele;EPHB1 gene;EPHB1 wt Allele;Ephrin Type-B Receptor 1, human;NET questionnaire;SLC6A2 gene;SLC6A2 wt Allele|net
Finding|Receptor|Hospital Course|6063,6066|false|false|false|C0812375;C0815327;C1366441;C1420212;C1704819;C1705456;C3853572;C3890893|ELK3 gene;ELK3 wt Allele;EPHB1 gene;EPHB1 wt Allele;Ephrin Type-B Receptor 1, human;NET questionnaire;SLC6A2 gene;SLC6A2 wt Allele|net
Finding|Classification|Hospital Course|6067,6075|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|6067,6075|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|6067,6075|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|Hospital Course|6067,6089|false|false|false|C0429652|Negative fluid balance|negative fluid balance
Drug|Substance|Hospital Course|6076,6081|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|6076,6081|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Organism Function|Hospital Course|6076,6089|false|false|false|C0016284|Fluid Balance|fluid balance
Drug|Organic Chemical|Hospital Course|6082,6089|false|false|false|C4319618|Balance (substance)|balance
Drug|Pharmacologic Substance|Hospital Course|6082,6089|false|false|false|C4319618|Balance (substance)|balance
Finding|Finding|Hospital Course|6082,6089|false|false|false|C0014653;C0560184|Ability to balance;Equilibrium|balance
Finding|Organism Function|Hospital Course|6082,6089|false|false|false|C0014653;C0560184|Ability to balance;Equilibrium|balance
Procedure|Diagnostic Procedure|Hospital Course|6082,6089|false|false|false|C2174421|examination of balance|balance
Finding|Idea or Concept|Hospital Course|6093,6097|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Finding|Intellectual Product|Hospital Course|6093,6097|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Finding|Intellectual Product|Hospital Course|6108,6114|false|false|false|C1547311|Patient Condition Code - Stable|stable
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6115,6120|false|false|false|C0022646|Kidney|renal
Disorder|Disease or Syndrome|Hospital Course|6115,6120|false|false|false|C0042075|Urologic Diseases|renal
Finding|Organ or Tissue Function|Hospital Course|6115,6129|false|false|false|C0232804|Renal function|renal function
Procedure|Laboratory Procedure|Hospital Course|6115,6129|false|false|false|C0022662|Kidney Function Tests|renal function
Finding|Finding|Hospital Course|6121,6129|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|Hospital Course|6121,6129|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|Hospital Course|6121,6129|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|Hospital Course|6121,6129|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Drug|Inorganic Chemical|Hospital Course|6131,6143|false|false|false|C0013832;C3536863|Electrolyte [EPC];Electrolytes|Electrolytes
Drug|Pharmacologic Substance|Hospital Course|6131,6143|false|false|false|C0013832;C3536863|Electrolyte [EPC];Electrolytes|Electrolytes
Finding|Idea or Concept|Hospital Course|6157,6161|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Finding|Intellectual Product|Hospital Course|6157,6161|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Finding|Idea or Concept|Hospital Course|6198,6202|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|6198,6202|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|6198,6202|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|6203,6213|false|false|false|C0054836|carvedilol|carvedilol
Drug|Pharmacologic Substance|Hospital Course|6203,6213|false|false|false|C0054836|carvedilol|carvedilol
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6221,6224|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6221,6224|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|6221,6224|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|6221,6224|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|6227,6239|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|Hospital Course|6227,6239|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6255,6265|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|Hospital Course|6255,6265|false|false|false|C0065374|lisinopril|lisinopril
Disorder|Disease or Syndrome|Hospital Course|6281,6286|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|Hospital Course|6281,6286|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|Hospital Course|6288,6296|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|Hospital Course|6288,6296|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|Hospital Course|6288,6296|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|Hospital Course|6288,6296|false|false|false|C0033095||pressure
Drug|Organic Chemical|Hospital Course|6297,6304|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|Hospital Course|6297,6304|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|Hospital Course|6297,6304|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Finding|Conceptual Entity|Hospital Course|6297,6304|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|Hospital Course|6297,6304|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|Hospital Course|6297,6304|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|Hospital Course|6319,6323|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|6319,6323|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|6319,6323|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|6324,6334|false|false|false|C0028066|nifedipine|nifedipine
Drug|Pharmacologic Substance|Hospital Course|6324,6334|false|false|false|C0028066|nifedipine|nifedipine
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6355,6358|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6355,6358|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|6355,6358|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|6355,6358|false|false|false|C1332410|BID gene|BID
Finding|Idea or Concept|Hospital Course|6370,6374|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Finding|Intellectual Product|Hospital Course|6370,6374|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Attribute|Clinical Attribute|Hospital Course|6375,6378|false|false|false|C0871470|Systolic Pressure|SBP
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6375,6378|false|false|false|C0085805|Androgen Binding Protein|SBP
Drug|Biologically Active Substance|Hospital Course|6375,6378|false|false|false|C0085805|Androgen Binding Protein|SBP
Finding|Gene or Genome|Hospital Course|6375,6378|false|false|false|C1705296;C3274833|CCHCR1 wt Allele;SHBG wt Allele|SBP
Procedure|Diagnostic Procedure|Hospital Course|6375,6378|false|false|false|C1306620|Systolic blood pressure measurement|SBP
Finding|Finding|Hospital Course|6401,6406|false|false|false|C0587267;C3810854|Close;Closed|close
Finding|Functional Concept|Hospital Course|6401,6406|false|false|false|C0587267;C3810854|Close;Closed|close
Disorder|Disease or Syndrome|Hospital Course|6407,6410|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6407,6410|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|Hospital Course|6407,6410|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6407,6410|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|Hospital Course|6407,6410|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|Hospital Course|6407,6410|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|Hospital Course|6407,6410|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|Hospital Course|6407,6410|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Finding|Gene or Genome|Hospital Course|6407,6410|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|Hospital Course|6407,6410|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Daily or Recreational Activity|Hospital Course|6431,6438|false|false|false|C3812400|Weights - exercise activity|weights
Disorder|Disease or Syndrome|Hospital Course|6443,6448|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|Hospital Course|6443,6448|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|Hospital Course|6443,6457|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Finding|Organism Function|Hospital Course|6443,6457|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Procedure|Health Care Activity|Hospital Course|6443,6457|false|false|false|C0005824|Blood pressure determination|blood pressure
Finding|Finding|Hospital Course|6449,6457|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|Hospital Course|6449,6457|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|Hospital Course|6449,6457|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|Hospital Course|6449,6457|false|false|false|C0033095||pressure
Drug|Organic Chemical|Hospital Course|6459,6466|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|Hospital Course|6459,6466|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|Hospital Course|6459,6466|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Finding|Conceptual Entity|Hospital Course|6459,6466|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|Hospital Course|6459,6466|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|Hospital Course|6459,6466|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Disorder|Disease or Syndrome|Hospital Course|6471,6483|false|false|false|C0020538|Hypertensive disease|Hypertension
Finding|Idea or Concept|Hospital Course|6506,6510|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|6506,6510|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|6506,6510|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|6511,6521|false|false|false|C0054836|carvedilol|carvedilol
Drug|Pharmacologic Substance|Hospital Course|6511,6521|false|false|false|C0054836|carvedilol|carvedilol
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6529,6532|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6529,6532|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|6529,6532|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|6529,6532|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|6535,6547|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|Hospital Course|6535,6547|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6563,6573|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|Hospital Course|6563,6573|false|false|false|C0065374|lisinopril|lisinopril
Disorder|Disease or Syndrome|Hospital Course|6589,6594|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|Hospital Course|6589,6594|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|Hospital Course|6596,6604|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|Hospital Course|6596,6604|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|Hospital Course|6596,6604|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|Hospital Course|6596,6604|false|false|false|C0033095||pressure
Drug|Organic Chemical|Hospital Course|6605,6612|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|Hospital Course|6605,6612|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|Hospital Course|6605,6612|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Finding|Conceptual Entity|Hospital Course|6605,6612|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|Hospital Course|6605,6612|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|Hospital Course|6605,6612|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|Hospital Course|6627,6631|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|6627,6631|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|6627,6631|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|6632,6642|false|false|false|C0028066|nifedipine|nifedipine
Drug|Pharmacologic Substance|Hospital Course|6632,6642|false|false|false|C0028066|nifedipine|nifedipine
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6663,6666|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6663,6666|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|6663,6666|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|6663,6666|false|false|false|C1332410|BID gene|BID
Finding|Idea or Concept|Hospital Course|6678,6682|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Finding|Intellectual Product|Hospital Course|6678,6682|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Attribute|Clinical Attribute|Hospital Course|6683,6686|false|false|false|C0871470|Systolic Pressure|SBP
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6683,6686|false|false|false|C0085805|Androgen Binding Protein|SBP
Drug|Biologically Active Substance|Hospital Course|6683,6686|false|false|false|C0085805|Androgen Binding Protein|SBP
Finding|Gene or Genome|Hospital Course|6683,6686|false|false|false|C1705296;C3274833|CCHCR1 wt Allele;SHBG wt Allele|SBP
Procedure|Diagnostic Procedure|Hospital Course|6683,6686|false|false|false|C1306620|Systolic blood pressure measurement|SBP
Disorder|Cell or Molecular Dysfunction|Hospital Course|6697,6705|false|false|false|C4727483|BRAF Gene Rearrangement|Positive
Finding|Classification|Hospital Course|6697,6705|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|Positive
Finding|Finding|Hospital Course|6697,6705|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|Positive
Finding|Body Substance|Hospital Course|6711,6718|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|6711,6718|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|6711,6718|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|Hospital Course|6719,6731|false|false|false|C0231221;C0332151|Asymptomatic (finding);Asymptomatic diagnosis of|asymptomatic
Finding|Functional Concept|Hospital Course|6756,6764|false|false|false|C1510439|bacteria aspects|bacteria
Finding|Finding|Hospital Course|6784,6796|false|false|false|C0231221;C0332151|Asymptomatic (finding);Asymptomatic diagnosis of|Asymptomatic
Finding|Sign or Symptom|Hospital Course|6806,6812|false|false|false|C0015967|Fever|fevers
Finding|Sign or Symptom|Hospital Course|6813,6820|false|false|false|C0013428|Dysuria|dysuria
Finding|Sign or Symptom|Hospital Course|6821,6828|false|false|false|C0231218|Malaise|malaise
Finding|Body Substance|Hospital Course|6830,6835|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Functional Concept|Hospital Course|6830,6835|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Intellectual Product|Hospital Course|6830,6835|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Procedure|Laboratory Procedure|Hospital Course|6830,6843|false|false|false|C0430404|Urine culture|Urine culture
Lab|Laboratory or Test Result|Hospital Course|6830,6852|false|false|false|C0853721|Culture urine negative|Urine culture negative
Drug|Biomedical or Dental Material|Hospital Course|6836,6843|false|false|false|C1706355|Culture Dose Form|culture
Finding|Functional Concept|Hospital Course|6836,6843|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Finding|Idea or Concept|Hospital Course|6836,6843|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Procedure|Laboratory Procedure|Hospital Course|6836,6843|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|culture
Lab|Laboratory or Test Result|Hospital Course|6836,6852|false|false|false|C0855652|Culture negative|culture negative
Finding|Classification|Hospital Course|6844,6852|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|6844,6852|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|6844,6852|false|false|false|C5237010|Expression Negative|negative
Finding|Functional Concept|Hospital Course|6857,6861|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Location or Region|Hospital Course|6868,6872|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6868,6872|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Hospital Course|6868,6872|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Hospital Course|6868,6872|false|false|false|C0740941|Lung Problem|lung
Disorder|Disease or Syndrome|Hospital Course|6868,6886|false|false|false|C0521530|Lung consolidation|lung consolidation
Disorder|Disease or Syndrome|Hospital Course|6873,6886|false|false|false|C0521530|Lung consolidation|consolidation
Finding|Functional Concept|Hospital Course|6888,6898|false|false|false|C0332448;C1546677;C1549537|Administration Method - Infiltrate;Infiltration|infiltrate
Finding|Intellectual Product|Hospital Course|6888,6898|false|false|false|C0332448;C1546677;C1549537|Administration Method - Infiltrate;Infiltration|infiltrate
Finding|Pathologic Function|Hospital Course|6888,6898|false|false|false|C0332448;C1546677;C1549537|Administration Method - Infiltrate;Infiltration|infiltrate
Finding|Finding|Hospital Course|6903,6912|false|false|false|C1405978;C1548000;C1548429|Encounter due to radiological examination;Radiology Section ID;radiology referral type|Radiology
Finding|Idea or Concept|Hospital Course|6903,6912|false|false|false|C1405978;C1548000;C1548429|Encounter due to radiological examination;Radiology Section ID;radiology referral type|Radiology
Finding|Intellectual Product|Hospital Course|6903,6912|false|false|false|C1405978;C1548000;C1548429|Encounter due to radiological examination;Radiology Section ID;radiology referral type|Radiology
Procedure|Diagnostic Procedure|Hospital Course|6903,6912|false|false|false|C0043299;C0807679;C1962945|Diagnostic radiologic examination;Radiographic imaging procedure;Radiology studies|Radiology
Finding|Conceptual Entity|Hospital Course|6913,6917|false|false|false|C0034754;C1705179;C4722184|Do Reading Question;Reading (activity);Reading (datum presentation)|read
Finding|Daily or Recreational Activity|Hospital Course|6913,6917|false|false|false|C0034754;C1705179;C4722184|Do Reading Question;Reading (activity);Reading (datum presentation)|read
Finding|Intellectual Product|Hospital Course|6913,6917|false|false|false|C0034754;C1705179;C4722184|Do Reading Question;Reading (activity);Reading (datum presentation)|read
Procedure|Laboratory Procedure|Hospital Course|6913,6917|false|false|false|C4723641|Nucleotide Sequence Read|read
Procedure|Health Care Activity|Hospital Course|6922,6931|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Procedure|Diagnostic Procedure|Hospital Course|6932,6935|false|false|false|C0039985|Plain chest X-ray|CXR
Drug|Organic Chemical|Hospital Course|6940,6945|true|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|Hospital Course|6940,6945|true|false|false|C3815497|Cough (guaifenesin)|cough
Finding|Sign or Symptom|Hospital Course|6940,6945|true|false|false|C0010200|Coughing|cough
Finding|Sign or Symptom|Hospital Course|6947,6953|true|false|false|C0015967|Fever|fevers
Disorder|Disease or Syndrome|Hospital Course|6955,6967|true|false|false|C0023518|Leukocytosis|leukocytosis
Finding|Finding|Hospital Course|6955,6967|true|false|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Finding|Functional Concept|Hospital Course|6989,6993|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Gene or Genome|Hospital Course|6989,6993|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Intellectual Product|Hospital Course|6989,6993|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Mental Process|Hospital Course|6989,6993|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Intellectual Product|Hospital Course|6994,7005|false|false|false|C1549438|Procedure Practitioner Identifier Code Type - Radiologist|radiologist
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7018,7027|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Hospital Course|7018,7027|false|false|false|C2707265||pulmonary
Finding|Finding|Hospital Course|7018,7027|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|Hospital Course|7018,7033|false|false|false|C0034063|Pulmonary Edema|pulmonary edema
Attribute|Clinical Attribute|Hospital Course|7028,7033|false|false|false|C1717255||edema
Finding|Pathologic Function|Hospital Course|7028,7033|false|false|false|C0013604|Edema|edema
Finding|Functional Concept|Hospital Course|7052,7058|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Finding|Finding|Hospital Course|7059,7066|false|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|Hospital Course|7059,7066|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Hospital Course|7070,7073|false|false|false|C0600500|Peptide Nucleic Acids|PNA
Finding|Conceptual Entity|Hospital Course|7074,7083|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Hospital Course|7074,7083|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Hospital Course|7074,7083|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7074,7083|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Finding|Idea or Concept|Hospital Course|7136,7147|false|false|false|C0750502|Significant|significant
Finding|Intellectual Product|Hospital Course|7148,7156|false|false|false|C1315013|Clinical NEC (not elsewhere classified in LNC)|clinical
Finding|Sign or Symptom|Hospital Course|7148,7165|true|false|false|C0037088|Signs and Symptoms|clinical findings
Attribute|Clinical Attribute|Hospital Course|7157,7165|true|false|false|C2926606||findings
Finding|Functional Concept|Hospital Course|7157,7165|true|false|false|C2607943|findings aspects|findings
Anatomy|Body Location or Region|Hospital Course|7170,7173|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Hospital Course|7170,7173|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Hospital Course|7170,7173|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Drug|Organic Chemical|Hospital Course|7193,7201|false|false|false|C0699129|Coumadin|Coumadin
Drug|Pharmacologic Substance|Hospital Course|7193,7201|false|false|false|C0699129|Coumadin|Coumadin
Finding|Idea or Concept|Hospital Course|7202,7206|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Finding|Intellectual Product|Hospital Course|7202,7206|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Finding|Finding|Hospital Course|7219,7224|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Hospital Course|7219,7224|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Pathologic Function|Hospital Course|7229,7237|false|false|false|C0087086;C0302148|Blood Clot;Thrombus|thrombus
Finding|Functional Concept|Hospital Course|7241,7245|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|Hospital Course|7241,7245|false|false|false|C0582103|Medical Examination|exam
Attribute|Clinical Attribute|Hospital Course|7253,7256|false|false|false|C0368980|Coagulation tissue factor induced.INR|INR
Procedure|Laboratory Procedure|Hospital Course|7253,7256|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7253,7256|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Finding|Idea or Concept|Hospital Course|7282,7286|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|7282,7286|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|7282,7286|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|7288,7296|false|false|false|C0699129|Coumadin|Coumadin
Drug|Pharmacologic Substance|Hospital Course|7288,7296|false|false|false|C0699129|Coumadin|Coumadin
Disorder|Disease or Syndrome|Hospital Course|7312,7318|false|false|false|C0002871|Anemia|Anemia
Finding|Finding|Hospital Course|7323,7328|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Hospital Course|7323,7328|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Anatomy|Body Location or Region|Hospital Course|7332,7340|false|false|false|C1548801|Body Site Modifier - External|external
Finding|Functional Concept|Hospital Course|7332,7340|false|false|false|C0521134|External route|external
Finding|Finding|Hospital Course|7341,7345|true|false|false|C5890125|Loss (adaptation)|loss
Finding|Pathologic Function|Hospital Course|7373,7379|false|false|false|C0025222|Melena|melena
Finding|Finding|Hospital Course|7393,7399|false|false|false|C0857322|Anemic|anemic
Drug|Biomedical or Dental Material|Hospital Course|7405,7413|false|false|false|C0168634|BaseLine dental cement|baseline
Finding|Idea or Concept|Hospital Course|7405,7413|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7434,7437|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Hospital Course|7434,7437|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|Hospital Course|7434,7437|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Hospital Course|7434,7437|false|false|false|C0019029|Hemoglobin concentration|Hgb
Finding|Finding|Hospital Course|7442,7448|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Idea or Concept|Hospital Course|7442,7448|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7453,7458|false|false|false|C0022646|Kidney|renal
Disorder|Disease or Syndrome|Hospital Course|7453,7458|false|false|false|C0042075|Urologic Diseases|renal
Disorder|Disease or Syndrome|Hospital Course|7453,7466|false|false|false|C0022658|Kidney Diseases|renal disease
Disorder|Disease or Syndrome|Hospital Course|7459,7466|false|false|false|C0012634|Disease|disease
Disorder|Disease or Syndrome|Hospital Course|7471,7474|false|false|false|C0002873;C1275685;C4554601;C5960004|Amyloidosis cutis dyschromia;Anemia of chronic disease;Angiokeratoma Corporis Diffusum;Avellino corneal dystrophy|ACD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7471,7474|false|false|false|C0050552;C1565285|ACD protein, human;acid citrate dextrose|ACD
Drug|Biologically Active Substance|Hospital Course|7471,7474|false|false|false|C0050552;C1565285|ACD protein, human;acid citrate dextrose|ACD
Drug|Indicator, Reagent, or Diagnostic Aid|Hospital Course|7471,7474|false|false|false|C0050552;C1565285|ACD protein, human;acid citrate dextrose|ACD
Drug|Organic Chemical|Hospital Course|7471,7474|false|false|false|C0050552;C1565285|ACD protein, human;acid citrate dextrose|ACD
Finding|Gene or Genome|Hospital Course|7471,7474|false|false|false|C1538901|ACD gene|ACD
Finding|Finding|Hospital Course|7483,7495|false|true|false|C0302845|Mean corpuscular volume above reference range|elevated MCV
Disorder|Virus|Hospital Course|7492,7495|false|true|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|Hospital Course|7492,7495|false|true|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|Hospital Course|7492,7495|false|true|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7492,7495|false|true|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Finding|Finding|Hospital Course|7507,7515|false|false|false|C0332149|Possible|possible
Finding|Finding|Hospital Course|7516,7531|false|true|false|C0206160|Reticulocytosis|reticulocytosis
Finding|Finding|Hospital Course|7544,7547|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Hospital Course|7544,7547|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Mental Process|Hospital Course|7548,7557|false|false|false|C0242114|Suspicion|suspicion
Drug|Organic Chemical|Hospital Course|7570,7578|false|false|false|C0699129|Coumadin|Coumadin
Drug|Pharmacologic Substance|Hospital Course|7570,7578|false|false|false|C0699129|Coumadin|Coumadin
Anatomy|Cell|Hospital Course|7594,7607|false|false|false|C0035286|Reticulocytes|Reticulocytes
Finding|Intellectual Product|Hospital Course|7652,7657|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Finding|Hospital Course|7658,7662|false|false|false|C5890125|Loss (adaptation)|loss
Anatomy|Cell Component|Hospital Course|7678,7681|false|false|false|C2263086|Nuclear cap binding complex location|CBC
Procedure|Laboratory Procedure|Hospital Course|7678,7681|false|false|false|C0009555|Complete Blood Count|CBC
Finding|Body Substance|Hospital Course|7706,7715|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|7706,7715|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|7706,7715|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|7706,7715|false|false|false|C0030685|Patient Discharge|discharge
Finding|Intellectual Product|Hospital Course|7720,7727|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|Hospital Course|7720,7727|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Disorder|Disease or Syndrome|Hospital Course|7720,7742|false|false|false|C1561643|Chronic Kidney Diseases|Chronic kidney disease
Finding|Classification|Hospital Course|7720,7749|false|false|false|C2074731|chronic kidney disease stage|Chronic kidney disease, stage
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7728,7734|false|false|false|C0022646;C0227665|Both kidneys;Kidney|kidney
Disorder|Neoplastic Process|Hospital Course|7728,7734|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|kidney
Finding|Sign or Symptom|Hospital Course|7728,7734|false|false|false|C0812426|Kidney problem|kidney
Procedure|Diagnostic Procedure|Hospital Course|7728,7734|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7728,7734|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Disorder|Disease or Syndrome|Hospital Course|7728,7742|false|false|false|C0022658|Kidney Diseases|kidney disease
Disorder|Disease or Syndrome|Hospital Course|7735,7742|false|false|false|C0012634|Disease|disease
Attribute|Clinical Attribute|Hospital Course|7744,7749|false|false|false|C1300072|Tumor stage|stage
Finding|Intellectual Product|Hospital Course|7744,7752|false|false|false|C0441772|Stage level 4|stage IV
Drug|Biomedical or Dental Material|Hospital Course|7754,7762|false|false|false|C0168634|BaseLine dental cement|baseline
Finding|Idea or Concept|Hospital Course|7754,7762|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Finding|Hospital Course|7768,7774|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|7768,7774|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Disorder|Disease or Syndrome|Hospital Course|7780,7783|false|false|false|C0020538|Hypertensive disease|HTN
Attribute|Clinical Attribute|Hospital Course|7806,7817|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Hospital Course|7806,7817|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|Hospital Course|7806,7817|false|false|false|C4284232|Medications|medications
Finding|Idea or Concept|Hospital Course|7842,7853|false|false|false|C0750502|Significant|significant
Finding|Functional Concept|Hospital Course|7854,7860|false|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7854,7860|false|false|false|C4319952|Change - procedure|change
Finding|Idea or Concept|Hospital Course|7880,7884|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|7880,7884|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|7880,7884|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|7885,7897|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|Hospital Course|7885,7897|false|false|false|C0286651|atorvastatin|atorvastatin
Finding|Idea or Concept|Hospital Course|7909,7913|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|7909,7913|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|7909,7913|false|false|false|C1553498|home health encounter|home
Finding|Body Substance|Hospital Course|7926,7933|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|7926,7933|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|7926,7933|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7948,7954|false|false|false|C0123677|insulin aspart, human|aspart
Drug|Hormone|Hospital Course|7948,7954|false|false|false|C0123677|insulin aspart, human|aspart
Drug|Pharmacologic Substance|Hospital Course|7948,7954|false|false|false|C0123677|insulin aspart, human|aspart
Disorder|Congenital Abnormality|Hospital Course|7955,7958|false|false|false|C1845118|SHORT STATURE, IDIOPATHIC, X-LINKED|ISS
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7964,7972|false|false|false|C0907402|insulin glargine|glargine
Drug|Hormone|Hospital Course|7964,7972|false|false|false|C0907402|insulin glargine|glargine
Drug|Pharmacologic Substance|Hospital Course|7964,7972|false|false|false|C0907402|insulin glargine|glargine
Finding|Idea or Concept|Hospital Course|7982,7986|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7987,8003|false|false|false|C5392125|Glycemic Control|glycemic control
Drug|Organic Chemical|Hospital Course|7996,8003|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|Hospital Course|7996,8003|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|Hospital Course|7996,8003|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Finding|Conceptual Entity|Hospital Course|7996,8003|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|Hospital Course|7996,8003|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|Hospital Course|7996,8003|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|Hospital Course|8006,8018|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Anatomy|Body Space or Junction|Hospital Course|8045,8048|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|Hospital Course|8045,8048|false|false|false|C0018802|Congestive heart failure|CHF
Drug|Organic Chemical|Hospital Course|8067,8072|false|false|false|C0699992|Lasix|lasix
Drug|Pharmacologic Substance|Hospital Course|8067,8072|false|false|false|C0699992|Lasix|lasix
Drug|Pharmacologic Substance|Hospital Course|8093,8102|false|false|false|C0012798|Diuretics|diuretics
Finding|Idea or Concept|Hospital Course|8116,8120|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|8116,8120|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|8116,8120|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|8132,8141|false|false|false|C0076840|torsemide|torsemide
Drug|Pharmacologic Substance|Hospital Course|8132,8141|false|false|false|C0076840|torsemide|torsemide
Procedure|Health Care Activity|Hospital Course|8165,8169|false|false|false|C1515187|Take|take
Drug|Food|Hospital Course|8173,8179|false|false|false|C0004722;C0939797;C2722028|Banana;banana allergenic extract;banana extract|banana
Drug|Immunologic Factor|Hospital Course|8173,8179|false|false|false|C0004722;C0939797;C2722028|Banana;banana allergenic extract;banana extract|banana
Drug|Organic Chemical|Hospital Course|8173,8179|false|false|false|C0004722;C0939797;C2722028|Banana;banana allergenic extract;banana extract|banana
Drug|Pharmacologic Substance|Hospital Course|8173,8179|false|false|false|C0004722;C0939797;C2722028|Banana;banana allergenic extract;banana extract|banana
Finding|Idea or Concept|Hospital Course|8217,8227|false|false|false|C1548386|Document Completion - incomplete|incomplete
Finding|Finding|Hospital Course|8228,8235|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|hearing
Finding|Physiologic Function|Hospital Course|8228,8235|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|hearing
Finding|Finding|Hospital Course|8237,8241|false|false|false|C5890125|Loss (adaptation)|loss
Finding|Idea or Concept|Hospital Course|8245,8248|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|8245,8248|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Body Substance|Hospital Course|8252,8261|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|8252,8261|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|8252,8261|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|8252,8261|false|false|false|C0030685|Patient Discharge|discharge
Drug|Organic Chemical|Hospital Course|8282,8289|false|false|false|C0163712|Relate - vinyl resin|related
Finding|Finding|Hospital Course|8282,8289|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|Hospital Course|8282,8289|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Drug|Pharmacologic Substance|Hospital Course|8294,8303|false|false|false|C0012798|Diuretics|diuretics
Disorder|Disease or Syndrome|Hospital Course|8319,8322|false|false|false|C0020538|Hypertensive disease|HTN
Drug|Organic Chemical|Hospital Course|8334,8344|false|false|false|C0028066|nifedipine|nifedipine
Drug|Pharmacologic Substance|Hospital Course|8334,8344|false|false|false|C0028066|nifedipine|nifedipine
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8356,8359|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8356,8359|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8356,8359|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|8356,8359|false|false|false|C1332410|BID gene|BID
Anatomy|Body Space or Junction|Hospital Course|8375,8379|false|false|false|C0228216|Structure of subparietal sulcus|SBPs
Finding|Idea or Concept|Hospital Course|8396,8400|false|false|false|C1552851|next - HtmlLinkType|next
Event|Activity|Hospital Course|8401,8413|false|false|false|C0003629|Appointments|appointments
Disorder|Disease or Syndrome|Hospital Course|8415,8421|false|false|false|C0002871|Anemia|Anemia
Disorder|Disease or Syndrome|Hospital Course|8454,8457|false|false|false|C0002873;C1275685;C4554601;C5960004|Amyloidosis cutis dyschromia;Anemia of chronic disease;Angiokeratoma Corporis Diffusum;Avellino corneal dystrophy|ACD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8454,8457|false|false|false|C0050552;C1565285|ACD protein, human;acid citrate dextrose|ACD
Drug|Biologically Active Substance|Hospital Course|8454,8457|false|false|false|C0050552;C1565285|ACD protein, human;acid citrate dextrose|ACD
Drug|Indicator, Reagent, or Diagnostic Aid|Hospital Course|8454,8457|false|false|false|C0050552;C1565285|ACD protein, human;acid citrate dextrose|ACD
Drug|Organic Chemical|Hospital Course|8454,8457|false|false|false|C0050552;C1565285|ACD protein, human;acid citrate dextrose|ACD
Finding|Gene or Genome|Hospital Course|8454,8457|false|false|false|C1538901|ACD gene|ACD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8459,8462|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Hospital Course|8459,8462|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|Hospital Course|8459,8462|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Hospital Course|8459,8462|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Health Care Activity|Hospital Course|8474,8483|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Anatomy|Body Location or Region|Hospital Course|8490,8493|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Hospital Course|8490,8493|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Hospital Course|8490,8493|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8508,8519|false|false|false|C0851145|on warfarin|on warfarin
Drug|Hazardous or Poisonous Substance|Hospital Course|8511,8519|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|Hospital Course|8511,8519|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|Hospital Course|8511,8519|false|false|false|C0043031|warfarin|warfarin
Finding|Idea or Concept|Hospital Course|8531,8540|false|false|false|C0549178|Continuous|continued
Event|Activity|Hospital Course|8542,8552|false|false|false|C1283169||monitoring
Procedure|Health Care Activity|Hospital Course|8542,8552|false|false|false|C0150369|Preventive monitoring|monitoring
Finding|Idea or Concept|Hospital Course|8565,8569|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|8565,8569|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|8565,8569|false|false|false|C1553498|home health encounter|home
Finding|Idea or Concept|Hospital Course|8582,8590|false|false|false|C4288901|In-House|in-house
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8603,8609|false|false|false|C0123677|insulin aspart, human|aspart
Drug|Hormone|Hospital Course|8603,8609|false|false|false|C0123677|insulin aspart, human|aspart
Drug|Pharmacologic Substance|Hospital Course|8603,8609|false|false|false|C0123677|insulin aspart, human|aspart
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8610,8618|false|false|false|C0907402|insulin glargine|glargine
Drug|Hormone|Hospital Course|8610,8618|false|false|false|C0907402|insulin glargine|glargine
Drug|Pharmacologic Substance|Hospital Course|8610,8618|false|false|false|C0907402|insulin glargine|glargine
Finding|Idea or Concept|Hospital Course|8634,8638|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|8634,8638|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|8634,8638|false|false|false|C1553498|home health encounter|home
Finding|Intellectual Product|Hospital Course|8639,8646|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8639,8646|false|false|false|C0040808|Treatment Protocols|regimen
Finding|Body Substance|Hospital Course|8648,8657|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|8648,8657|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|8648,8657|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|8648,8657|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|8658,8664|false|false|false|C0944911||weight
Finding|Finding|Hospital Course|8658,8664|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|Hospital Course|8658,8664|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|Hospital Course|8658,8664|false|false|false|C1305866|Weighing patient|weight
Finding|Body Substance|Hospital Course|8671,8680|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|8671,8680|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|8671,8680|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|8671,8680|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|8691,8702|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|8691,8702|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Hospital Course|8691,8702|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|8691,8715|false|false|false|C1627937|Medications on admission|Medications on Admission
Procedure|Health Care Activity|Hospital Course|8706,8715|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|Hospital Course|8734,8744|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Hospital Course|8734,8744|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|Hospital Course|8734,8749|false|false|false|C0746470|MEDICATION LIST|Medication list
Finding|Intellectual Product|Hospital Course|8745,8749|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Drug|Organic Chemical|Hospital Course|8766,8774|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Hospital Course|8766,8774|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Hospital Course|8766,8774|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Finding|Functional Concept|Hospital Course|8766,8774|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|8766,8774|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|Hospital Course|8779,8792|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|8779,8792|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|8779,8792|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|Hospital Course|8811,8814|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|8815,8819|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|8815,8819|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|8815,8819|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Hospital Course|8823,8828|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|Hospital Course|8823,8828|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Drug|Organic Chemical|Hospital Course|8833,8840|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Hospital Course|8833,8840|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|Hospital Course|8860,8872|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|8860,8872|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|Hospital Course|8890,8900|false|false|false|C0054836|carvedilol|Carvedilol
Drug|Pharmacologic Substance|Hospital Course|8890,8900|false|false|false|C0054836|carvedilol|Carvedilol
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8912,8915|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8912,8915|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8912,8915|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|8912,8915|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|8920,8928|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|8920,8928|false|false|false|C1692318|docusate|Docusate
Drug|Organic Chemical|Hospital Course|8920,8935|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|Hospital Course|8920,8935|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|Hospital Course|8929,8935|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|8929,8935|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|8929,8935|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Finding|Physiologic Function|Hospital Course|8929,8935|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|8929,8935|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8946,8949|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8946,8949|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8946,8949|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|8946,8949|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|8954,8964|false|false|false|C0060926|gabapentin|Gabapentin
Drug|Pharmacologic Substance|Hospital Course|8954,8964|false|false|false|C0060926|gabapentin|Gabapentin
Finding|Finding|Hospital Course|8979,8995|false|false|false|C0027796;C3714625|Neuralgia;Neuropathic pain|neuropathic pain
Finding|Sign or Symptom|Hospital Course|8979,8995|false|false|false|C0027796;C3714625|Neuralgia;Neuropathic pain|neuropathic pain
Attribute|Clinical Attribute|Hospital Course|8991,8995|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|8991,8995|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|8991,8995|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9000,9010|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|Hospital Course|9000,9010|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Organic Chemical|Hospital Course|9030,9043|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|Hospital Course|9030,9043|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|Hospital Course|9030,9043|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Biomedical or Dental Material|Hospital Course|9046,9049|false|false|false|C0039225|Tablet Dosage Form|TAB
Drug|Organic Chemical|Hospital Course|9063,9073|false|false|false|C0028066|nifedipine|NIFEdipine
Drug|Pharmacologic Substance|Hospital Course|9063,9073|false|false|false|C0028066|nifedipine|NIFEdipine
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9086,9089|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9086,9089|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9086,9089|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|9086,9089|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|9095,9108|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Pharmacologic Substance|Hospital Course|9095,9108|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Finding|Gene or Genome|Hospital Course|9128,9131|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Location or Region|Hospital Course|9132,9137|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|9132,9137|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|9132,9142|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Hospital Course|9132,9142|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Hospital Course|9138,9142|false|true|false|C2598155||pain
Finding|Functional Concept|Hospital Course|9138,9142|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|9138,9142|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|9148,9160|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Pharmacologic Substance|Hospital Course|9148,9160|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Biomedical or Dental Material|Hospital Course|9180,9192|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Drug|Organic Chemical|Hospital Course|9180,9192|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Drug|Organic Chemical|Hospital Course|9180,9199|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Pharmacologic Substance|Hospital Course|9180,9199|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Hazardous or Poisonous Substance|Hospital Course|9193,9199|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Drug|Organic Chemical|Hospital Course|9193,9199|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Drug|Organic Chemical|Hospital Course|9219,9224|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|Hospital Course|9219,9224|false|false|false|C3489575|sennosides, USP|Senna
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9235,9238|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9235,9238|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9235,9238|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|9235,9238|false|false|false|C1332410|BID gene|BID
Finding|Sign or Symptom|Hospital Course|9239,9251|false|false|false|C0009806|Constipation|constipation
Drug|Organic Chemical|Hospital Course|9257,9264|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|9257,9264|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|9257,9264|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|Hospital Course|9257,9266|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|Hospital Course|9257,9266|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|Hospital Course|9257,9266|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|Hospital Course|9257,9266|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|Hospital Course|9257,9266|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Drug|Hazardous or Poisonous Substance|Hospital Course|9290,9298|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|Hospital Course|9290,9298|false|false|false|C0043031|warfarin|Warfarin
Drug|Pharmacologic Substance|Hospital Course|9290,9298|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|Hospital Course|9320,9331|false|false|false|C0002144|allopurinol|Allopurinol
Drug|Pharmacologic Substance|Hospital Course|9320,9331|false|false|false|C0002144|allopurinol|Allopurinol
Finding|Idea or Concept|Hospital Course|9354,9357|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|DAY
Finding|Intellectual Product|Hospital Course|9354,9357|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|DAY
Drug|Organic Chemical|Hospital Course|9363,9372|false|false|false|C0076840|torsemide|Torsemide
Drug|Pharmacologic Substance|Hospital Course|9363,9372|false|false|false|C0076840|torsemide|Torsemide
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9393,9400|false|false|false|C0020171;C0020172;C3538423|Humulin;Humulin S;Humulin insulin|HumuLIN
Drug|Hormone|Hospital Course|9393,9400|false|false|false|C0020171;C0020172;C3538423|Humulin;Humulin S;Humulin insulin|HumuLIN
Drug|Pharmacologic Substance|Hospital Course|9393,9400|false|false|false|C0020171;C0020172;C3538423|Humulin;Humulin S;Humulin insulin|HumuLIN
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9393,9406|false|false|false|C0306367|HumuLIN 70/30|HumuLIN 70/30
Drug|Hormone|Hospital Course|9393,9406|false|false|false|C0306367|HumuLIN 70/30|HumuLIN 70/30
Drug|Pharmacologic Substance|Hospital Course|9393,9406|false|false|false|C0306367|HumuLIN 70/30|HumuLIN 70/30
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9408,9415|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|Hospital Course|9408,9415|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|Hospital Course|9408,9415|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Finding|Gene or Genome|Hospital Course|9408,9415|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|Hospital Course|9408,9415|false|false|false|C0202098|Insulin measurement|insulin
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9408,9419|false|false|false|C0021658|insulin isophane|insulin NPH
Drug|Hormone|Hospital Course|9408,9419|false|false|false|C0021658|insulin isophane|insulin NPH
Drug|Pharmacologic Substance|Hospital Course|9408,9419|false|false|false|C0021658|insulin isophane|insulin NPH
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9416,9419|false|false|false|C0027442|Nasopharynx|NPH
Disorder|Disease or Syndrome|Hospital Course|9416,9419|false|false|false|C0020258|Hydrocephalus, Normal Pressure|NPH
Finding|Functional Concept|Hospital Course|9460,9472|false|false|false|C1522438|Subcutaneous Route of Administration|subcutaneous
Finding|Daily or Recreational Activity|Hospital Course|9487,9493|false|false|false|C4048877|Dinner|dinner
Finding|Body Substance|Hospital Course|9498,9507|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|9498,9507|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|9498,9507|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|9498,9507|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|9498,9519|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|9508,9519|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|9508,9519|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Hospital Course|9508,9519|false|false|false|C4284232|Medications|Medications
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9524,9531|false|false|false|C0020171;C0020172;C3538423|Humulin;Humulin S;Humulin insulin|HumuLIN
Drug|Hormone|Hospital Course|9524,9531|false|false|false|C0020171;C0020172;C3538423|Humulin;Humulin S;Humulin insulin|HumuLIN
Drug|Pharmacologic Substance|Hospital Course|9524,9531|false|false|false|C0020171;C0020172;C3538423|Humulin;Humulin S;Humulin insulin|HumuLIN
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9524,9537|false|false|false|C0306367|HumuLIN 70/30|HumuLIN 70/30
Drug|Hormone|Hospital Course|9524,9537|false|false|false|C0306367|HumuLIN 70/30|HumuLIN 70/30
Drug|Pharmacologic Substance|Hospital Course|9524,9537|false|false|false|C0306367|HumuLIN 70/30|HumuLIN 70/30
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9539,9546|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|Hospital Course|9539,9546|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|Hospital Course|9539,9546|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Finding|Gene or Genome|Hospital Course|9539,9546|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|Hospital Course|9539,9546|false|false|false|C0202098|Insulin measurement|insulin
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9539,9550|false|false|false|C0021658|insulin isophane|insulin NPH
Drug|Hormone|Hospital Course|9539,9550|false|false|false|C0021658|insulin isophane|insulin NPH
Drug|Pharmacologic Substance|Hospital Course|9539,9550|false|false|false|C0021658|insulin isophane|insulin NPH
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9547,9550|false|false|false|C0027442|Nasopharynx|NPH
Disorder|Disease or Syndrome|Hospital Course|9547,9550|false|false|false|C0020258|Hydrocephalus, Normal Pressure|NPH
Finding|Functional Concept|Hospital Course|9591,9603|false|false|false|C1522438|Subcutaneous Route of Administration|subcutaneous
Finding|Daily or Recreational Activity|Hospital Course|9618,9624|false|false|false|C4048877|Dinner|dinner
Drug|Hazardous or Poisonous Substance|Hospital Course|9629,9637|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|Hospital Course|9629,9637|false|false|false|C0043031|warfarin|Warfarin
Drug|Pharmacologic Substance|Hospital Course|9629,9637|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|Hospital Course|9658,9665|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|9658,9665|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|9658,9665|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|Hospital Course|9658,9667|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|Hospital Course|9658,9667|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|Hospital Course|9658,9667|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|Hospital Course|9658,9667|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|Hospital Course|9658,9667|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Drug|Organic Chemical|Hospital Course|9690,9703|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|9690,9703|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|9690,9703|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|Hospital Course|9722,9725|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|9726,9730|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|9726,9730|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|9726,9730|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Hospital Course|9734,9739|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|Hospital Course|9734,9739|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Drug|Organic Chemical|Hospital Course|9744,9755|false|false|false|C0002144|allopurinol|Allopurinol
Drug|Pharmacologic Substance|Hospital Course|9744,9755|false|false|false|C0002144|allopurinol|Allopurinol
Finding|Idea or Concept|Hospital Course|9778,9781|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|DAY
Finding|Intellectual Product|Hospital Course|9778,9781|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|DAY
Drug|Organic Chemical|Hospital Course|9786,9793|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Hospital Course|9786,9793|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|Hospital Course|9813,9825|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|9813,9825|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|Hospital Course|9843,9851|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|9843,9851|false|false|false|C1692318|docusate|Docusate
Drug|Organic Chemical|Hospital Course|9843,9858|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|Hospital Course|9843,9858|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|Hospital Course|9852,9858|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|9852,9858|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|9852,9858|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Finding|Physiologic Function|Hospital Course|9852,9858|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|9852,9858|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9869,9872|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9869,9872|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9869,9872|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|9869,9872|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|9877,9887|false|false|false|C0060926|gabapentin|Gabapentin
Drug|Pharmacologic Substance|Hospital Course|9877,9887|false|false|false|C0060926|gabapentin|Gabapentin
Finding|Finding|Hospital Course|9902,9918|false|false|false|C0027796;C3714625|Neuralgia;Neuropathic pain|neuropathic pain
Finding|Sign or Symptom|Hospital Course|9902,9918|false|false|false|C0027796;C3714625|Neuralgia;Neuropathic pain|neuropathic pain
Attribute|Clinical Attribute|Hospital Course|9914,9918|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|9914,9918|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|9914,9918|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9924,9934|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|Hospital Course|9924,9934|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Organic Chemical|Hospital Course|9955,9968|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|Hospital Course|9955,9968|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|Hospital Course|9955,9968|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Biomedical or Dental Material|Hospital Course|9971,9974|false|false|false|C0039225|Tablet Dosage Form|TAB
Drug|Organic Chemical|Hospital Course|9989,10002|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Pharmacologic Substance|Hospital Course|9989,10002|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Finding|Gene or Genome|Hospital Course|10022,10025|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Location or Region|Hospital Course|10026,10031|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|10026,10031|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|10026,10036|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Hospital Course|10026,10036|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Hospital Course|10032,10036|false|true|false|C2598155||pain
Finding|Functional Concept|Hospital Course|10032,10036|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|10032,10036|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Biomedical or Dental Material|Hospital Course|10042,10054|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Drug|Organic Chemical|Hospital Course|10042,10054|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Drug|Organic Chemical|Hospital Course|10042,10061|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Pharmacologic Substance|Hospital Course|10042,10061|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Hazardous or Poisonous Substance|Hospital Course|10055,10061|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Drug|Organic Chemical|Hospital Course|10055,10061|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Drug|Organic Chemical|Hospital Course|10081,10086|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|Hospital Course|10081,10086|false|false|false|C3489575|sennosides, USP|Senna
Disorder|Mental or Behavioral Dysfunction|Hospital Course|10097,10100|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10097,10100|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|10097,10100|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|10097,10100|false|false|false|C1332410|BID gene|BID
Finding|Sign or Symptom|Hospital Course|10101,10113|false|false|false|C0009806|Constipation|constipation
Drug|Organic Chemical|Hospital Course|10119,10128|false|false|false|C0076840|torsemide|Torsemide
Drug|Pharmacologic Substance|Hospital Course|10119,10128|false|false|false|C0076840|torsemide|Torsemide
Drug|Organic Chemical|Hospital Course|10149,10158|false|false|false|C0076840|torsemide|torsemide
Drug|Pharmacologic Substance|Hospital Course|10149,10158|false|false|false|C0076840|torsemide|torsemide
Drug|Biomedical or Dental Material|Hospital Course|10167,10173|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|10177,10185|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|10180,10185|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|10180,10185|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Intellectual Product|Hospital Course|10186,10190|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Biomedical or Dental Material|Hospital Course|10208,10214|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|10215,10222|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|10230,10242|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Pharmacologic Substance|Hospital Course|10230,10242|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Organic Chemical|Hospital Course|10262,10272|false|false|false|C0054836|carvedilol|Carvedilol
Drug|Pharmacologic Substance|Hospital Course|10262,10272|false|false|false|C0054836|carvedilol|Carvedilol
Disorder|Mental or Behavioral Dysfunction|Hospital Course|10282,10285|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10282,10285|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|10282,10285|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|10282,10285|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|10291,10301|false|false|false|C0028066|nifedipine|NIFEdipine
Drug|Pharmacologic Substance|Hospital Course|10291,10301|false|false|false|C0028066|nifedipine|NIFEdipine
Disorder|Mental or Behavioral Dysfunction|Hospital Course|10314,10317|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10314,10317|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|10314,10317|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|10314,10317|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|10323,10333|false|false|false|C0028066|nifedipine|nifedipine
Drug|Pharmacologic Substance|Hospital Course|10323,10333|false|false|false|C0028066|nifedipine|nifedipine
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10342,10349|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|Hospital Course|10342,10349|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|Hospital Course|10342,10349|false|false|false|C0006935|capsule (pharmacologic)|capsule
Finding|Functional Concept|Hospital Course|10353,10361|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|10356,10361|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|10356,10361|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10386,10393|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|10386,10393|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|10386,10393|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Finding|Idea or Concept|Hospital Course|10394,10401|false|false|false|C0807726|refill|Refills
Finding|Body Substance|Hospital Course|10408,10417|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|10408,10417|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|10408,10417|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|10408,10417|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|10408,10429|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|10408,10429|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|10418,10429|false|false|false|C2926604||Disposition
Procedure|Health Care Activity|Hospital Course|10418,10429|false|false|false|C0184758|Patient disposition|Disposition
Finding|Idea or Concept|Hospital Course|10431,10435|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|10431,10435|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|10431,10435|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|Hospital Course|10441,10448|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|Hospital Course|10441,10448|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Finding|Intellectual Product|Hospital Course|10451,10459|false|false|false|C4695111|ADMIN.FACILITY|Facility
Finding|Body Substance|Hospital Course|10467,10476|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|10467,10476|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|10467,10476|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|10467,10476|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|10467,10486|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|10477,10486|false|false|false|C0945731||Diagnosis
Finding|Classification|Hospital Course|10477,10486|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|10477,10486|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|10477,10486|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Intellectual Product|Principle Diagnosis|10507,10512|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Finding|Intellectual Product|Principle Diagnosis|10516,10523|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Principle Diagnosis|10516,10523|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|Principle Diagnosis|10538,10562|false|false|false|C0018802|Congestive heart failure|congestive Heart Failure
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|10549,10554|false|false|false|C0018787;C4037974|Chest>Heart;Heart|Heart
Disorder|Neoplastic Process|Principle Diagnosis|10549,10554|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|Heart
Finding|Sign or Symptom|Principle Diagnosis|10549,10554|false|false|false|C0795691|HEART PROBLEM|Heart
Disorder|Disease or Syndrome|Principle Diagnosis|10549,10562|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|Heart Failure
Finding|Functional Concept|Principle Diagnosis|10555,10562|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|Failure
Finding|Idea or Concept|Principle Diagnosis|10555,10562|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|Failure
Finding|Individual Behavior|Principle Diagnosis|10555,10562|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|Failure
Disorder|Disease or Syndrome|Principle Diagnosis|10563,10575|false|false|false|C0020538|Hypertensive disease|Hypertension
Disorder|Neoplastic Process|Principle Diagnosis|10577,10586|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Finding|Functional Concept|Principle Diagnosis|10577,10586|false|false|false|C1522484|metastatic qualifier|Secondary
Procedure|Diagnostic Procedure|Principle Diagnosis|10587,10596|false|false|false|C0011900|Diagnosis|Diagnoses
Disorder|Disease or Syndrome|Principle Diagnosis|10598,10604|false|false|false|C0002871|Anemia|Anemia
Disorder|Disease or Syndrome|Principle Diagnosis|10605,10613|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|Diabetes
Disorder|Disease or Syndrome|Principle Diagnosis|10605,10622|false|false|false|C0011849|Diabetes Mellitus|Diabetes mellitus
Attribute|Clinical Attribute|Principle Diagnosis|10629,10633|false|false|false|C4318566|Deep Resection Margin|deep
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|10629,10638|false|false|false|C0226514|Structure of deep vein|deep vein
Disorder|Disease or Syndrome|Principle Diagnosis|10629,10649|false|false|false|C0149871;C0340708|Deep Vein Thrombosis;Deep vein thrombosis of lower limb|deep vein thrombosis
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|10634,10638|false|false|false|C0042449|Veins|vein
Finding|Pathologic Function|Principle Diagnosis|10634,10649|false|false|false|C0042487|Venous Thrombosis|vein thrombosis
Finding|Pathologic Function|Principle Diagnosis|10639,10649|false|false|false|C0040053|Thrombosis|thrombosis
Finding|Intellectual Product|Principle Diagnosis|10650,10657|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|Principle Diagnosis|10650,10657|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Disorder|Disease or Syndrome|Principle Diagnosis|10650,10672|false|false|false|C1561643|Chronic Kidney Diseases|Chronic Kidney Disease
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|10658,10664|false|false|false|C0022646;C0227665|Both kidneys;Kidney|Kidney
Disorder|Neoplastic Process|Principle Diagnosis|10658,10664|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|Kidney
Finding|Sign or Symptom|Principle Diagnosis|10658,10664|false|false|false|C0812426|Kidney problem|Kidney
Procedure|Diagnostic Procedure|Principle Diagnosis|10658,10664|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|Kidney
Procedure|Therapeutic or Preventive Procedure|Principle Diagnosis|10658,10664|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|Kidney
Disorder|Disease or Syndrome|Principle Diagnosis|10658,10672|false|false|false|C0022658|Kidney Diseases|Kidney Disease
Disorder|Disease or Syndrome|Principle Diagnosis|10665,10672|false|false|false|C0012634|Disease|Disease
Finding|Mental Process|Discharge Condition|10697,10703|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|10697,10710|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|10697,10710|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|10704,10710|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|10704,10710|false|false|false|C1546481|What subject filter - Status|Status
Finding|Idea or Concept|Discharge Condition|10712,10717|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Finding|Discharge Condition|10722,10730|false|false|false|C4068804|Coherent|coherent
Attribute|Clinical Attribute|Discharge Condition|10732,10754|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|10732,10754|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Finding|Finding|Discharge Condition|10741,10754|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|10741,10754|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|10756,10761|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|10756,10761|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|10756,10761|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|Discharge Condition|10756,10761|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|10756,10761|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|10756,10761|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|10766,10777|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|10779,10787|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|10779,10787|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|10779,10787|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|10788,10794|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|10788,10794|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|Discharge Condition|10796,10806|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|10796,10806|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|10796,10806|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|10796,10806|false|false|false|C1561560|ambulatory encounter|Ambulatory
Finding|Finding|Discharge Condition|10809,10820|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Condition|10809,10820|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Conceptual Entity|Discharge Instructions|10890,10899|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Discharge Instructions|10890,10899|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Discharge Instructions|10890,10899|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10890,10899|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|10920,10925|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|10920,10925|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Discharge Instructions|10920,10925|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|Discharge Instructions|10920,10933|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Finding|Functional Concept|Discharge Instructions|10926,10933|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|Discharge Instructions|10926,10933|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|Discharge Instructions|10926,10933|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Disorder|Disease or Syndrome|Discharge Instructions|10938,10950|false|false|false|C0020538|Hypertensive disease|hypertension
Drug|Pharmacologic Substance|Discharge Instructions|10970,10979|false|false|false|C0012798|Diuretics|diuretics
Finding|Conceptual Entity|Discharge Instructions|10986,10997|false|false|false|C2986411|Improvement|improvement
Finding|Functional Concept|Discharge Instructions|11006,11014|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Discharge Instructions|11006,11014|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Lab|Laboratory or Test Result|Discharge Instructions|11016,11020|false|false|false|C0587081|Laboratory test finding|labs
Finding|Functional Concept|Discharge Instructions|11025,11029|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|Discharge Instructions|11025,11029|false|false|false|C0582103|Medical Examination|exam
Disorder|Disease or Syndrome|Discharge Instructions|11057,11062|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|Discharge Instructions|11057,11062|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|Discharge Instructions|11057,11071|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Finding|Organism Function|Discharge Instructions|11057,11071|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Procedure|Health Care Activity|Discharge Instructions|11057,11071|false|false|false|C0005824|Blood pressure determination|blood pressure
Finding|Finding|Discharge Instructions|11063,11071|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|Discharge Instructions|11063,11071|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|Discharge Instructions|11063,11071|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|Discharge Instructions|11063,11071|false|false|false|C0033095||pressure
Attribute|Clinical Attribute|Discharge Instructions|11072,11083|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|11072,11083|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|Discharge Instructions|11072,11083|false|false|false|C4284232|Medications|medications
Finding|Idea or Concept|Discharge Instructions|11109,11113|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Discharge Instructions|11109,11113|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Discharge Instructions|11109,11113|false|false|false|C1553498|home health encounter|home
Drug|Pharmacologic Substance|Discharge Instructions|11115,11124|false|false|false|C0013227|Pharmaceutical Preparations|medicines
Finding|Intellectual Product|Discharge Instructions|11137,11145|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|Discharge Instructions|11137,11145|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|Discharge Instructions|11153,11157|false|false|false|C1947933|care activity|care
Finding|Finding|Discharge Instructions|11153,11157|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|11153,11157|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|11153,11160|false|false|false|C1555558|care of - AddressPartType|care of
Drug|Amino Acid, Peptide, or Protein|Discharge Instructions|11186,11190|false|false|false|C3273412|NCK-Interacting Protein with SH3 Domain|wish
Finding|Gene or Genome|Discharge Instructions|11186,11190|false|false|false|C1423524;C3273411|NCKIPSD gene;NCKIPSD wt Allele|wish
Disorder|Disease or Syndrome|Discharge Instructions|11204,11208|false|false|false|C0339510|Vitelliform Macular Dystrophy|best
Finding|Gene or Genome|Discharge Instructions|11204,11208|false|false|false|C1826421;C5781213|BEST1 gene;BEST1 wt Allele|best
Procedure|Health Care Activity|Discharge Instructions|11229,11237|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|11238,11250|false|false|false|C3263700||Instructions
Finding|Intellectual Product|Discharge Instructions|11238,11250|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

