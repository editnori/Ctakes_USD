CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Known|Modifier|false|false||Knownnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Adverse reaction to drug|Finding|true|false||Adverse Drug Reactionsnull|Adverse reaction to drug|Finding|true|false||Drug Reactionsnull|Pharmaceutical Preparations|Drug|false|false||Drug
null|Pharmacologic Substance|Drug|false|false||Drugnull|Drug problem|Finding|false|false||Drugnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Chief complaint (finding)|Finding|false|false||Chief Complaintnull|Complaint (finding)|Finding|false|false||Complaintnull|null|Attribute|false|false||Complaintnull|Chest Pain|Finding|false|false||Chest painnull|null|Attribute|false|false||Chest painnull|Chest problem|Finding|false|false||Chestnull|Chest|Anatomy|false|false||Chest
null|Anterior thoracic region|Anatomy|false|false||Chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Cardiac catheterisation as the cause of abnormal reaction of the patient, or of later complication, without mention of misadventure at the time of the procedure|Disorder|false|false||Cardiac catheterizationnull|Diagnostic Service Section ID - Cardiac Catheterization|Finding|false|false||Cardiac catheterizationnull|Consent Type - Cardiac Catheterization|Procedure|false|false||Cardiac catheterization
null|Cardiac Catheterization Procedures|Procedure|false|false||Cardiac catheterizationnull|Cardiac attachment|Finding|false|false||Cardiacnull|Heart|Anatomy|false|false||Cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||Cardiacnull|Catheterization|Procedure|false|false||catheterizationnull|Stenting|Procedure|false|false||stentingnull|null|Device|false|false||stentingnull|Drug-Eluting Stents|Device|false|false||drug eluting stentnull|Pharmaceutical Preparations|Drug|false|false||drug
null|Pharmacologic Substance|Drug|false|false||drugnull|Drug problem|Finding|false|false||drugnull|null|Device|false|false||stentnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Circumflex|Modifier|false|false||circumflexnull|History of present illness (finding)|Finding|false|false||History of Present Illnessnull|null|Attribute|false|false||History of Present Illnessnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Present illness|Finding|false|false||Present Illnessnull|Present|Finding|false|false||Present
null|Presentation|Finding|false|false||Presentnull|Illness (finding)|Finding|false|false||Illnessnull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Old|Time|false|false||oldnull|Woman|Subject|false|false||woman
null|Human, Female adult|Subject|false|false||womannull|diastolic congestive heart failure|Disorder|false|false||diastolic CHFnull|Diastole|Attribute|false|false||diastolicnull|Congestive heart failure|Disorder|false|false||CHFnull|Choroidal fissure|Anatomy|false|false||CHFnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Hypertensive disease|Disorder|false|false||HTNnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Leukocyte adhesion deficiency type 1|Disorder|false|false||LAD
null|Leukocyte adhesion deficiency|Disorder|false|false||LADnull|ITGB2 wt Allele|Finding|false|false||LAD
null|DLD gene|Finding|false|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false||LADnull|Ladino Language|Entity|false|false||LADnull|Stenting|Procedure|false|false||stentingnull|null|Device|false|false||stentingnull|Repeat Object|Finding|false|false||repeat
null|Repeat|Finding|false|false||repeatnull|Repeat Pattern|Time|false|false||repeatnull|Stenting|Procedure|false|false||stentingnull|null|Device|false|false||stentingnull|DES protein, human|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|DES protein, human|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DESnull|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|Disorder|false|false||DESnull|DES gene|Finding|false|false||DESnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Episode of|Time|false|false||episodesnull|Past 2 Weeks|Time|false|false||past 2 weeksnull|2 Weeks|Time|false|false||2 weeksnull|week|Time|false|false||weeksnull|Tightness sensation quality|Modifier|false|false||tightnessnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Usually|Finding|false|false||usuallynull|Usual|Modifier|false|false||usuallynull|Exertion|Finding|false|false||exertionnull|Residential flat|Device|false|false||flatnull|Flat shape|Modifier|false|false||flatnull|Night time|Time|false|false||at nightnull|Night time|Time|false|false||nightnull|At rest (qualifier value)|Finding|false|false||at restnull|REST protein, human|Drug|false|false||rest
null|REST protein, human|Drug|false|false||restnull|REST gene|Finding|false|false||rest
null|site-specific telomere resolvase activity|Finding|false|false||rest
null|Rest|Finding|false|false||restnull|To the left (qualifier value)|Modifier|false|false||to the leftnull|Left upper arm structure|Anatomy|false|false||left arm
null|Left arm|Anatomy|false|false||left armnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Anorectal Malformations|Disorder|false|false||armnull|AKR1A1 wt Allele|Finding|false|false||arm
null|ARMC9 gene|Finding|false|false||armnull|Protocol Treatment Arm|Procedure|false|false||arm
null|Axillary Reverse Mapping|Procedure|false|false||arm
null|Study Arm|Procedure|false|false||armnull|Upper arm|Anatomy|false|false||arm
null|null|Anatomy|false|false||arm
null|Upper Extremity|Anatomy|false|false||armnull|GLAUCOMA, NORMAL TENSION, SUSCEPTIBILITY TO|Finding|false|false||NTG
null|OPA1 wt Allele|Finding|false|false||NTG
null|OPA1 gene|Finding|false|false||NTGnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Somewhat|Finding|false|false||Somewhatnull|Different|Modifier|false|false||differentnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|null|Time|false|false||prior tonull|null|Time|false|false||priornull|Act Relationship Subset - previous|Time|false|false||previous
null|Previous|Time|false|false||previousnull|Structure of cisterna pontis|Anatomy|false|false||PCIsnull|Lightheadedness|Finding|false|false||lightheadednessnull|More|LabModifier|false|false||morenull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Episode of|Time|false|false||episodenull|Initial (abbreviation)|Finding|false|false||initialnull|Initially|Time|false|false||initialnull|Firstly|Modifier|false|false||initialnull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Plain chest X-ray|Procedure|false|false||CXRnull|Negative|Finding|false|false||negative fornull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Process Pharmacologic Substance|Drug|false|false||processnull|Process (qualifier value)|Finding|false|false||processnull|bony process|Anatomy|false|false||processnull|Process|Phenomenon|false|false||processnull|Laboratory test finding|Lab|false|false||Labsnull|Negative|Finding|false|false||for negativenull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Troponin|Drug|false|false||troponin
null|Troponin|Drug|false|false||troponinnull|Troponin measurement|Procedure|false|false||troponinnull|null|Time|false|false||prior tonull|null|Time|false|false||priornull|Arylsulfatase A, human|Drug|false|false||ASA
null|Arylsulfatase A, human|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASAnull|ARSA gene|Finding|false|false||ASAnull|null|Time|false|false||prior tonull|null|Time|false|false||priornull|Transfer - product ownership|Finding|false|false||transfer
null|Transfer Technique|Finding|false|false||transfer
null|ActClass - transfer|Finding|false|false||transfer
null|null|Finding|false|false||transfernull|Transfer (immobility management)|Procedure|false|false||transfernull|arrival - ActRelationshipType|Finding|false|false||arrivalnull|null|Event|false|false||arrivalnull|Floor (anatomic)|Anatomy|false|false||floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Feeling comfortable|Finding|false|false||comfortablenull|Chest problem|Finding|true|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Review of systems (procedure)|Procedure|false|false||REVIEW OF SYSTEMSnull|null|Attribute|false|false||REVIEW OF SYSTEMS
null|null|Attribute|false|false||REVIEW OF SYSTEMSnull|Review of|Finding|false|false||REVIEW OFnull|Review (Publication Type)|Finding|false|false||REVIEW
null|Act Class - review|Finding|false|false||REVIEWnull|System|Finding|false|false||SYSTEMSnull|Proline dehydrogenase deficiency|Disorder|false|false||HPInull|History of present illness (finding)|Finding|false|false||HPI
null|allene oxide synthase activity|Finding|false|false||HPInull|In addition to|Finding|false|false||addition
null|Add - instruction imperative|Finding|false|false||additionnull|Fever|Finding|true|false||feversnull|Chills|Finding|false|false||chillsnull|Sweating|Finding|false|false||sweats
null|Sweat|Finding|false|false||sweatsnull|Presyncope|Finding|false|false||presyncopenull|Syncope|Finding|false|false||syncopenull|Syncope <Gastrophryninae>|Entity|false|false||syncopenull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Paroxysmal nocturnal dyspnea|Disorder|false|false||PNDnull|NPPA wt Allele|Finding|false|false||PND
null|NPPA gene|Finding|false|false||PNDnull|sleeping upright or using specific number of extra pillows (orthopnea)|Finding|false|false||orthopnea
null|Orthopnea|Finding|false|false||orthopneanull|Leg|Anatomy|false|false||leg
null|Lower Extremity|Anatomy|false|false||legnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Abdominal Pain|Finding|false|false||abdominal painnull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Vomiting|Finding|false|false||vomitingnull|Hematemesis|Finding|false|false||hematemesisnull|rectal discharge diarrhea (physical finding)|Finding|false|false||diarrhea
null|Diarrhea|Finding|false|false||diarrheanull|Constipation|Finding|false|false||constipationnull|DYRK3 gene|Finding|false|false||red
null|Redness|Finding|false|false||red
null|IK gene|Finding|false|false||rednull|Radiological Exposure Device|Device|false|false||rednull|Red color|Modifier|false|false||rednull|null|Finding|false|false||black stools
null|Melena|Finding|false|false||black stoolsnull|Black - ethnic group (ethnic group)|Subject|false|false||black
null|Black race|Subject|false|false||black
null|African|Subject|false|false||blacknull|Black - Structured Product Labeling Color|Modifier|false|false||black
null|Black color|Modifier|false|false||blacknull|Feces|Finding|false|false||stoolsnull|null|Attribute|false|false||stoolsnull|Stool seat|Device|false|false||stoolsnull|Dysuria|Finding|false|false||dysurianull|Hematuria|Disorder|false|false||hematurianull|Myalgia|Finding|false|false||myalgiasnull|Arthralgia|Finding|false|false||arthralgiasnull|Eruption of skin (disorder)|Disorder|false|false||rashnull|Skin rash|Finding|false|false||rash
null|Eruptions|Finding|false|false||rash
null|Exanthema|Finding|false|false||rashnull|Medical History|Finding|true|false||history ofnull|History of present illness (finding)|Finding|true|false||history
null|History of previous events|Finding|true|false||history
null|Historical aspects qualifier|Finding|true|false||history
null|Medical History|Finding|true|false||history
null|Concept History|Finding|true|false||historynull|History|Subject|false|false||historynull|Deep thrombophlebitis|Disorder|true|false||DVT
null|Deep Vein Thrombosis|Disorder|true|false||DVTnull|area DVT|Anatomy|true|false||DVTnull|null|Attribute|true|false||DVTnull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Leukocyte adhesion deficiency type 1|Disorder|false|false||LAD
null|Leukocyte adhesion deficiency|Disorder|false|false||LADnull|ITGB2 wt Allele|Finding|false|false||LAD
null|DLD gene|Finding|false|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false||LADnull|Ladino Language|Entity|false|false||LADnull|Stenting|Procedure|false|false||stentingnull|null|Device|false|false||stentingnull|Repeat Object|Finding|false|false||repeat
null|Repeat|Finding|false|false||repeatnull|Repeat Pattern|Time|false|false||repeatnull|Stenting|Procedure|false|false||stentingnull|null|Device|false|false||stentingnull|DES protein, human|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|DES protein, human|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DESnull|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|Disorder|false|false||DESnull|DES gene|Finding|false|false||DESnull|diastolic congestive heart failure|Disorder|false|false||Diastolic CHFnull|Diastole|Attribute|false|false||Diastolicnull|Congestive heart failure|Disorder|false|false||CHFnull|Choroidal fissure|Anatomy|false|false||CHFnull|Hypertensive disease|Disorder|false|false||HTNnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Cancer patients and suicide and depression|Disorder|false|false||Depression
null|Mental Depression|Disorder|false|false||Depression
null|Depressive disorder|Disorder|false|false||Depression
null|Depressed mood|Disorder|false|false||Depressionnull|Depression - motion|Finding|false|false||Depression
null|null|Finding|false|false||Depressionnull|Depression - recess|Modifier|false|false||Depressionnull|Pain of right shoulder region|Finding|false|false||Right shoulder pain
null|right shoulder joint pain|Finding|false|false||Right shoulder painnull|Structure of right shoulder region|Anatomy|false|false||Right shouldernull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Shoulder Pain|Finding|false|false||shoulder painnull|Examination of shoulder(s)|Procedure|false|false||shoulder
null|Procedures on Shoulder|Procedure|false|false||shouldernull|Upper extremity>Shoulder|Anatomy|false|false||shoulder
null|Shoulder|Anatomy|false|false||shouldernull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Bursitis|Disorder|false|false||bursitisnull|Rotator Cuff Injuries|Disorder|false|false||rotator cuff injurynull|Rotator Cuff|Anatomy|false|false||rotator cuffnull|null|Device|false|false||rotatornull|Cuffing (morphologic abnormality)|Finding|false|false||cuffnull|Cuff - body part|Anatomy|false|false||cuffnull|Cuff Device|Device|false|false||cuffnull|Traumatic AND/OR non-traumatic injury|Disorder|false|false||injury
null|Traumatic injury|Disorder|false|false||injurynull|Social and personal history|Finding|false|false||Social History
null|Social History|Finding|false|false||Social Historynull|Social|Finding|false|false||Socialnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Family Medical History|Finding|false|false||Family Historynull|Entity Name Part Type - family|Finding|false|false||Family
null|Last Name|Finding|false|false||Family
null|Living Arrangement - Family|Finding|false|false||Family
null|Family (taxonomic)|Finding|false|false||Family
null|Family Collection|Finding|false|false||Familynull|Family|Subject|false|false||Familynull|History of present illness (finding)|Finding|false|true||History
null|History of previous events|Finding|false|true||History
null|Historical aspects qualifier|Finding|false|true||History
null|Medical History|Finding|false|true||History
null|Concept History|Finding|false|true||Historynull|History|Subject|false|false||Historynull|Ward (environment)|Device|false|false||wardnull|Ward (person)|Subject|false|false||wardnull|Ward (environment)|Entity|false|false||wardnull|ErbB Receptors|Drug|false|false||her family
null|ErbB Receptors|Drug|false|false||her familynull|ErbB Receptors|Finding|false|false||her familynull|Entity Name Part Type - family|Finding|true|false||family
null|Last Name|Finding|true|false||family
null|Living Arrangement - Family|Finding|true|false||family
null|Family (taxonomic)|Finding|true|false||family
null|Family Collection|Finding|true|false||familynull|Family|Subject|false|false||familynull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|physical examination (physical finding)|Finding|false|false||physical examnull|Physical Examination|Procedure|false|false||physical examnull|physical examination (physical finding)|Finding|false|false||physical
null|Physical|Finding|false|false||physicalnull|Physical Examination|Procedure|false|false||physicalnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GENERALnull|General medical service|Procedure|false|false||GENERALnull|Generalized|Modifier|false|false||GENERALnull|Woman|Subject|false|false||woman
null|Human, Female adult|Subject|false|false||womannull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|Oriented to place|Finding|false|false||Orientednull|Orientation, Spatial|Modifier|false|false||Orientednull|Mood (psychological function)|Finding|false|false||Mood
null|mood (physical finding)|Finding|false|false||Mood
null|Mood (attribute)|Finding|false|false||Moodnull|null|Attribute|false|false||Moodnull|Affect (mental function)|Finding|false|false||affectnull|assessment of affect|Procedure|false|false||affectnull|Appropriate|Modifier|false|false||appropriatenull|HEENT|Anatomy|false|false||HEENTnull|Scleral Diseases|Disorder|false|false||Scleranull|examination of sclera|Procedure|false|false||Scleranull|Sclera|Anatomy|false|false||Scleranull|Anicteric|Finding|false|false||anictericnull|Pupil equal round and reacting to light|Finding|false|false||PERRLnull|Malignant neoplasm of conjunctiva|Disorder|false|false||Conjunctiva
null|Benign neoplasm of conjunctiva|Disorder|false|false||Conjunctiva
null|Conjunctival Diseases|Disorder|false|false||Conjunctivanull|Specimen Type - Conjunctiva|Finding|false|false||Conjunctiva
null|null|Finding|false|false||Conjunctivanull|examination of conjunctiva|Procedure|false|false||Conjunctiva
null|Procedure on conjunctiva|Procedure|false|false||Conjunctivanull|Structure of palpebral conjunctiva|Anatomy|false|false||Conjunctiva
null|conjunctiva|Anatomy|false|false||Conjunctivanull|Pink color|Modifier|false|false||pinknull|Pallor of skin|Finding|true|false||pallornull|Cyanosis|Finding|true|false||cyanosisnull|Oral mucous membrane structure|Anatomy|false|false||oral mucosanull|Oral Dosage Form|Drug|false|false||oralnull|Oral Route of Administration|Finding|false|false||oral
null|Oral (intended site)|Finding|false|false||oralnull|Oral cavity|Anatomy|false|false||oralnull|Oral|Modifier|false|false||oralnull|null|Finding|false|false||mucosanull|Mucous Membrane|Anatomy|false|false||mucosanull|Passive joint movement of neck (finding)|Finding|false|false||NECK
null|Neck problem|Finding|false|false||NECKnull|dendritic spine neck|Anatomy|false|false||NECK
null|Neck|Anatomy|false|false||NECKnull|Supple|Finding|false|false||Supplenull|Jugular venous pressure|Finding|false|false||JVPnull|Cardiac attachment|Finding|false|false||CARDIACnull|Heart|Anatomy|false|false||CARDIACnull|Cardiac - anatomy qualifier|Modifier|false|false||CARDIACnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Palpation|Procedure|false|false||palpationnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||breastnull|Breast problem|Finding|false|false||breastnull|Procedures on breast|Procedure|false|false||breastnull|Breast|Anatomy|false|false||breastnull|Lung|Anatomy|false|false||LUNGSnull|Respiratory, thoracic and mediastinal disorders|Disorder|false|false||Respnull|Respiratory rate|Attribute|false|false||Respnull|Unlabored|Finding|false|false||unlaborednull|Use of accessory muscles|Finding|true|false||accessory muscle usenull|Accessory skeletal muscle|Disorder|true|false||accessory musclenull|Accessory|Device|true|false||accessorynull|Muscle (organ)|Anatomy|false|false||muscle
null|Muscle Tissue|Anatomy|false|false||musclenull|Use - dosing instruction imperative|Finding|true|false||use
null|utilization qualifier|Finding|true|false||use
null|Usage|Finding|true|false||usenull|cetrimonium bromide|Drug|false|false||CTABnull|Malignant neoplasm of abdomen|Disorder|false|false||ABDOMENnull|Abdomen problem|Finding|false|false||ABDOMENnull|Abdomen|Anatomy|false|false||ABDOMEN
null|Abdominal Cavity|Anatomy|false|false||ABDOMENnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|LRRC4B gene|Finding|true|false||HSMnull|Emotional tenderness|Finding|true|false||tenderness
null|Sore to touch|Finding|true|false||tendernessnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false||Abdnull|ABD (body structure)|Anatomy|false|false||Abd
null|Abdomen|Anatomy|false|false||Abdnull|Procedure on aorta|Procedure|false|false||aortanull|Chest+Abdomen>Aorta|Anatomy|false|false||aorta
null|Aorta|Anatomy|false|false||aortanull|Palpation|Procedure|false|false||palpationnull|Bruit|Finding|true|false||bruitsnull|All extremities|Anatomy|false|false||EXTREMITIES
null|Limb structure|Anatomy|false|false||EXTREMITIESnull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||SKIN
null|Skin and subcutaneous tissue disorders|Disorder|false|false||SKINnull|Skin Specimen Source Code|Finding|false|false||SKIN
null|Skin Specimen|Finding|false|false||SKINnull|Skin, Human|Anatomy|false|false||SKIN
null|Skin|Anatomy|false|false||SKINnull|Stasis dermatitis|Disorder|true|false||stasis dermatitisnull|Stasis|Finding|false|false||stasisnull|Dermatitis|Disorder|true|false||dermatitisnull|Ulcer|Finding|true|false||ulcersnull|Scar Tissue|Finding|true|false||scars
null|Cicatrix|Finding|true|false||scarsnull|Xanthoma|Disorder|true|false||xanthomasnull|null|Drug|false|false||PULSESnull|Physiologic pulse|Finding|false|false||PULSESnull|Pulse taking|Procedure|false|false||PULSESnull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Carotid Arteries|Anatomy|false|false||Carotidnull|Femur|Anatomy|false|false||Femoralnull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Carotid Arteries|Anatomy|false|false||Carotidnull|Femur|Anatomy|false|false||Femoralnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|physical examination (physical finding)|Finding|false|false||physical examnull|Physical Examination|Procedure|false|false||physical examnull|physical examination (physical finding)|Finding|false|false||physical
null|Physical|Finding|false|false||physicalnull|Physical Examination|Procedure|false|false||physicalnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|SAT1 protein, human|Drug|false|false||Sat
null|SAT1 protein, human|Drug|false|false||Satnull|College Entrance Examination Board Scholastic Aptitude Test|Finding|false|false||Sat
null|SAT1 wt Allele|Finding|false|false||Sat
null|SAT1 gene|Finding|false|false||Satnull|Santali language|Entity|false|false||Satnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Generalnull|General medical service|Procedure|false|false||Generalnull|Generalized|Modifier|false|false||Generalnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|BORNHOLM EYE DISEASE|Disorder|false|false||bednull|Bachelor of Education|Finding|false|false||bednull|Beds|Device|false|false||bednull|Patient Location - Bed|Modifier|false|false||bednull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|HEENT|Anatomy|false|false||HEENTnull|Myelofibrosis|Disorder|false|false||MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false||MMMnull|Passive joint movement of neck (finding)|Finding|false|false||Neck
null|Neck problem|Finding|false|false||Necknull|dendritic spine neck|Anatomy|false|false||Neck
null|Neck|Anatomy|false|false||Necknull|Supple|Finding|false|false||Supplenull|Jugular venous engorgement|Finding|true|false||JVDnull|Lung|Anatomy|false|false||Lungsnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Auscultation|Procedure|false|false||auscultationnull|Basilar Rales|Finding|true|false||crackles
null|Rales|Finding|true|false||cracklesnull|Wheezing|Finding|false|false||wheezesnull|Lymphoma, Mixed-Cell, Follicular|Disorder|false|false||Nmlnull|RRP8 gene|Finding|false|false||Nmlnull|Work of Breathing|Finding|false|false||work of breathingnull|Work|Event|false|false||worknull|outcomes otolaryngology breathing|Finding|false|false||breathing
null|Inspiration (function)|Finding|false|false||breathing
null|Respiration|Finding|false|false||breathingnull|null|Attribute|false|false||breathingnull|respiratory system process|Phenomenon|false|false||breathingnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false||Abdnull|ABD (body structure)|Anatomy|false|false||Abd
null|Abdomen|Anatomy|false|false||Abdnull|Obesity|Disorder|false|false||Obesenull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|Hereditary Multiple Exostoses|Disorder|false|false||Extnull|EXT1 wt Allele|Finding|false|false||Ext
null|EXT1 gene|Finding|false|false||Extnull|PDSS1 gene|Finding|false|false||DPsnull|Disintegration per Second|LabModifier|false|false||DPsnull|Clubbing|Disorder|true|false||clubbingnull|Cyanosis|Finding|true|false||cyanosisnull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|Laboratory test finding|Lab|false|false||labsnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Monos|Drug|false|false||Monos
null|Mono-S|Drug|false|false||Monos
null|Monos|Drug|false|false||Monosnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||Eos
null|Familial eosinophilia|Disorder|false|false||Eosnull|PRSS33 gene|Finding|false|false||Eos
null|IKZF4 gene|Finding|false|false||Eosnull|Eos <Loriini>|Entity|false|false||Eosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Maxillary left lateral incisor mesial prosthesis|Device|false|false||10PMnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Laboratory test finding|Lab|false|false||labsnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Cardiac enzymes|Drug|false|false||Cardiac enzymes
null|Cardiac enzymes|Drug|false|false||Cardiac enzymesnull|Cardiac enzymes/isoenzymes measurement|Procedure|false|false||Cardiac enzymesnull|null|Attribute|false|false||Cardiac enzymesnull|Cardiac attachment|Finding|false|false||Cardiacnull|Heart|Anatomy|false|false||Cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||Cardiacnull|Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM|Drug|false|false||enzymes
null|Enzymes, peripheral vasodilators|Drug|false|false||enzymes
null|Enzymes, peripheral vasodilators|Drug|false|false||enzymes
null|Enzymes, peripheral vasodilators|Drug|false|false||enzymes
null|Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM|Drug|false|false||enzymes
null|Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM|Drug|false|false||enzymes
null|Enzymes, antithrombotic|Drug|false|false||enzymes
null|Enzymes, antithrombotic|Drug|false|false||enzymes
null|Enzymes, antithrombotic|Drug|false|false||enzymes
null|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS|Drug|false|false||enzymes
null|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS|Drug|false|false||enzymes
null|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS|Drug|false|false||enzymes
null|Enzymes, hematological|Drug|false|false||enzymes
null|Enzymes, hematological|Drug|false|false||enzymes
null|Enzymes, hematological|Drug|false|false||enzymes
null|Enzymes|Drug|false|false||enzymes
null|Enzymes|Drug|false|false||enzymes
null|Enzymes for ALIMENTARY TRACT AND METABOLISM|Drug|false|false||enzymes
null|Enzymes for ALIMENTARY TRACT AND METABOLISM|Drug|false|false||enzymes
null|Enzymes for ALIMENTARY TRACT AND METABOLISM|Drug|false|false||enzymesnull|enzymology|Finding|false|false||enzymesnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Creatine Kinase|Drug|false|false||CPK
null|Creatine Kinase|Drug|false|false||CPKnull|PIK3C2A gene|Finding|false|false||CPKnull|Creatine kinase measurement|Procedure|false|false||CPKnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MB
null|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MBnull|creatine kinase activity|Finding|false|false||CK-MBnull|Serum creatine phosphokinase MB isoenzyme measurement|Procedure|false|false||CK-MB
null|Creatine kinase MB measurement|Procedure|false|false||CK-MBnull|MB 2|Drug|false|false||MB-2null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|Sinus rhythm|Finding|false|false||Sinus rhythm
null|null|Finding|false|false||Sinus rhythmnull|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false||Sinus
null|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false||Sinusnull|pathologic fistula|Disorder|false|false||Sinusnull|Sinus - general anatomical term|Anatomy|false|false||Sinus
null|Nasal sinus|Anatomy|false|false||Sinusnull|Rhythm|Finding|false|false||rhythm
null|rhythmic process (biological)|Finding|false|false||rhythmnull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Fracture of second cervical vertebra|Disorder|false|false||axisnull|Axis vertebra|Anatomy|false|false||axisnull|Genus Axis|Entity|false|false||axisnull|Axis|Modifier|false|false||axisnull|Finding of electrocardiogram PR interval|Finding|false|false||PR intervalnull|PR interval feature|Attribute|false|false||PR intervalnull|Parameterized Data Type - Interval|Finding|false|false||intervalnull|Interval|Time|false|false||intervalnull|Slightly (qualifier value)|Modifier|false|false||slightly
null|Slight (qualifier value)|Modifier|false|false||slightlynull|Greater Than|LabModifier|false|false||more thannull|More|LabModifier|false|false||morenull|null|Time|false|false||priornull|Electrocardiogram image|Finding|false|false||ekg
null|Electrocardiogram|Finding|false|false||ekgnull|Electrocardiography|Procedure|false|false||ekgnull|null|Procedure|false|false||Q wavenull|Q wave|Attribute|false|false||Q wavenull|WASF1 gene|Finding|false|false||wavenull|null|Phenomenon|false|false||wavenull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Nuclear stress test|Procedure|false|false||Nuclear Stress Testnull|Nuclear (incident type)|Modifier|false|false||Nuclear
null|Nuclear (nucleus)|Modifier|false|false||Nuclearnull|Exercise stress test|Procedure|false|false||Stress Test
null|Stress Test|Procedure|false|false||Stress Testnull|Stress bismuth subsalicylate|Drug|false|false||Stress
null|Stress bismuth subsalicylate|Drug|false|false||Stressnull|Stress|Finding|false|false||Stressnull|W stress|Attribute|false|false||Stressnull|Tests (qualifier value)|Finding|false|false||Test
null|Testing|Finding|false|false||Testnull|Laboratory Procedures|Procedure|false|false||Testnull|Test - temporal region|Anatomy|false|false||Testnull|Test Result|Lab|false|false||Testnull|Test Dosing Unit|LabModifier|false|false||Testnull|Interpretation Process|Finding|false|false||INTERPRETATIONnull|null|Attribute|false|false||INTERPRETATIONnull|Image Quality|Modifier|false|false||image qualitynull|Intrauterine growth restriction, metaphyseal dysplasia, adrenal hypoplasia congenita, and genital anomaly syndrome|Disorder|false|false||imagenull|Image (foundation metadata concept)|Finding|false|false||image
null|Image|Finding|false|false||image
null|Medical Image|Finding|false|false||image
null|image - dosage form|Finding|false|false||imagenull|Integrated Molecular Analysis of Genomes and their Expression Consortium|Entity|false|false||imagenull|Quality|Modifier|false|false||qualitynull|Adequate|Modifier|false|false||adequate
null|Sufficient|Modifier|false|false||adequatenull|Limited component (foundation metadata concept)|Finding|false|false||limited
null|Limited (extensiveness)|Finding|false|false||limitednull|Neck+Chest>Soft tissue|Anatomy|false|false||soft tissue
null|soft tissue|Anatomy|false|false||soft tissuenull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|Tissue Specimen Code|Finding|false|false||tissuenull|Body tissue|Anatomy|false|false||tissuenull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||breastnull|Breast problem|Finding|false|false||breastnull|Procedures on breast|Procedure|false|false||breastnull|Breast|Anatomy|false|false||breastnull|Attenuation|Event|false|false||attenuationnull|Activity (animal life circumstance)|Finding|false|false||activity
null|Physical activity|Finding|false|false||activitynull|Activities|Event|false|false||activitynull|null|Modifier|false|false||activitynull|Adjacent|Modifier|false|false||adjacent tonull|Adjacent|Modifier|false|false||adjacentnull|Malignant neoplasm of heart|Disorder|false|false||heart
null|benign neoplasm of heart|Disorder|false|false||heartnull|HEART PROBLEM|Finding|false|false||heartnull|Chest>Heart|Anatomy|false|false||heart
null|Heart|Anatomy|false|false||heartnull|REST protein, human|Drug|false|false||rest
null|REST protein, human|Drug|false|false||restnull|REST gene|Finding|false|false||rest
null|site-specific telomere resolvase activity|Finding|false|false||rest
null|Rest|Finding|false|false||restnull|Stress bismuth subsalicylate|Drug|false|false||stress
null|Stress bismuth subsalicylate|Drug|false|false||stressnull|Stress|Finding|false|false||stressnull|W stress|Attribute|false|false||stressnull|Left ventricular cavity size|Attribute|false|false||Left ventricular cavity sizenull|Cavity of left ventricle|Anatomy|false|false||Left ventricular cavitynull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Cavity of ventricle|Anatomy|false|false||ventricular cavitynull|Heart Ventricle|Anatomy|false|false||ventricularnull|Ventricular|Modifier|false|false||ventricularnull|Dental caries|Disorder|false|false||cavity
null|Cavitation|Disorder|false|false||cavitynull|Body cavities|Anatomy|false|false||cavitynull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|REST protein, human|Drug|false|false||Rest
null|REST protein, human|Drug|false|false||Restnull|REST gene|Finding|false|false||Rest
null|site-specific telomere resolvase activity|Finding|false|false||Rest
null|Rest|Finding|false|false||Restnull|Stress bismuth subsalicylate|Drug|false|false||stress
null|Stress bismuth subsalicylate|Drug|false|false||stressnull|Stress|Finding|false|false||stressnull|W stress|Attribute|false|false||stressnull|Perfusion (biological)|Finding|false|false||perfusion
null|Perfusion route|Finding|false|false||perfusionnull|Chemotherapeutic Perfusion|Procedure|false|false||perfusion
null|Perfusion (procedure)|Procedure|false|false||perfusionnull|Reversible|Finding|false|false||reversiblenull|Moderate - Severity of Illness Code|Finding|false|false||moderate
null|Moderate|Finding|false|false||moderatenull|Moderate (severity modifier)|Modifier|false|false||moderate
null|Moderate - Allergy Severity|Modifier|false|false||moderate
null|Moderation|Modifier|false|false||moderatenull|Reduced|Finding|false|false||reductionnull|Reduction procedure|Procedure|false|false||reduction
null|Surgical reduction|Procedure|false|false||reductionnull|Reduction (chemical)|Phenomenon|false|false||reductionnull|Photons|Drug|false|false||photonnull|counts|LabModifier|false|false||countsnull|Middle|Modifier|false|false||midnull|Basal|Modifier|false|false||basalnull|Inferolateral|Modifier|false|false||inferolateralnull|Walls of a building|Device|false|false||wallsnull|Distal Resection Margin|Attribute|false|false||distalnull|Distal (qualifier value)|Modifier|false|false||distalnull|Lateral|Modifier|false|false||lateralnull|Walls of a building|Device|false|false||wallnull|Wall motion|Attribute|false|false||wall motionnull|Walls of a building|Device|false|false||wallnull|Motion|Phenomenon|false|false||motionnull|Calculated Left Ventricular Ejection Fraction|Procedure|false|false||calculated left ventricular ejection fractionnull|Left ventricular ejection fraction|Attribute|false|false||left ventricular ejection fraction
null|null|Attribute|false|false||left ventricular ejection fractionnull|Left ventricular ejection|Finding|false|false||left ventricular ejectionnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Ventricular Ejection Fraction|Lab|false|false||ventricular ejection fractionnull|Ventricular ejection|Finding|false|false||ventricular ejectionnull|Heart Ventricle|Anatomy|false|false||ventricularnull|Ventricular|Modifier|false|false||ventricularnull|stress echo measurements ejection fraction|Finding|false|false||ejection fraction
null|Ejection fraction|Finding|false|false||ejection fractionnull|Ejection fraction (procedure)|Procedure|false|false||ejection fractionnull|Ejection as a Sports activity|Finding|false|false||ejectionnull|Ejection time|Attribute|false|false||ejectionnull|Ejection as a Circumstance of Injury|Phenomenon|false|false||ejectionnull|MDFAttributeType - Fraction|Finding|false|false||fractionnull|Fraction of|LabModifier|false|false||fractionnull|End Diastolic Volume Imaging|Procedure|false|false||EDVnull|Workstation|Device|false|false||workstationnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Reversible|Finding|false|false||Reversiblenull|Medium (Substance)|Drug|false|false||medium
null|Culture Media|Drug|false|false||mediumnull|A Medium Amount of Time|Finding|false|false||medium
null|Communications Media|Finding|false|false||medium
null|A Medium Amount|Finding|false|false||mediumnull|Message Waiting Priority - Medium|Modifier|false|false||medium
null|medium exposure|Modifier|false|false||mediumnull|Medium|LabModifier|false|false||mediumnull|Moderate (severity modifier)|Modifier|false|false||moderate severitynull|Moderate - Severity of Illness Code|Finding|false|false||moderate
null|Moderate|Finding|false|false||moderatenull|Moderate (severity modifier)|Modifier|false|false||moderate
null|Moderate - Allergy Severity|Modifier|false|false||moderate
null|Moderation|Modifier|false|false||moderatenull|With intensity|Modifier|false|false||severity
null|Severities|Modifier|false|false||severitynull|Perfusion (biological)|Finding|false|false||perfusion
null|Perfusion route|Finding|false|false||perfusionnull|Chemotherapeutic Perfusion|Procedure|false|false||perfusion
null|Perfusion (procedure)|Procedure|false|false||perfusionnull|THYROID HORMONE PLASMA MEMBRANE TRANSPORT DEFECT|Disorder|false|false||defectnull|Defect|Finding|false|false||defectnull|Methylcytosine Dioxygenase TET1|Drug|false|false||LCx
null|Methylcytosine Dioxygenase TET1|Drug|false|false||LCxnull|TET1 wt Allele|Finding|false|false||LCx
null|TET1 gene|Finding|false|false||LCxnull|Territory|Entity|false|false||territory
null|Geographic state|Entity|false|false||territorynull|Left ventricular cavity size|Attribute|false|false||left ventricular cavity sizenull|Cavity of left ventricle|Anatomy|false|false||left ventricular cavitynull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Cavity of ventricle|Anatomy|false|false||ventricular cavitynull|Heart Ventricle|Anatomy|false|false||ventricularnull|Ventricular|Modifier|false|false||ventricularnull|Dental caries|Disorder|false|false||cavity
null|Cavitation|Disorder|false|false||cavitynull|Body cavities|Anatomy|false|false||cavitynull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Systole|Finding|false|false||systolicnull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|null|Time|false|false||priornull|Study Object|Finding|false|false||studynull|Scientific Study|Procedure|false|false||study
null|Study|Procedure|false|false||study
null|Clinical Research|Procedure|false|false||studynull|Room of building - Study|Device|false|false||studynull|THYROID HORMONE PLASMA MEMBRANE TRANSPORT DEFECT|Disorder|false|false||defectnull|Defect|Finding|false|false||defectnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Cardiac catheterisation as the cause of abnormal reaction of the patient, or of later complication, without mention of misadventure at the time of the procedure|Disorder|false|false||Cardiac catheterizationnull|Diagnostic Service Section ID - Cardiac Catheterization|Finding|false|false||Cardiac catheterizationnull|Consent Type - Cardiac Catheterization|Procedure|false|false||Cardiac catheterization
null|Cardiac Catheterization Procedures|Procedure|false|false||Cardiac catheterizationnull|Cardiac attachment|Finding|false|false||Cardiacnull|Heart|Anatomy|false|false||Cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||Cardiacnull|Catheterization|Procedure|false|false||catheterizationnull|Published Comment|Finding|false|false||COMMENTS
null|Comment|Finding|false|false||COMMENTSnull|Consent Type - Coronary Angiography|Procedure|false|false||coronary angiography
null|Coronary angiography|Procedure|false|false||coronary angiographynull|Heart|Anatomy|false|false||coronarynull|Coronary|Modifier|false|false||coronarynull|angiogram|Procedure|false|false||angiographynull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Dominant|Finding|false|false||dominantnull|System (basic dose form)|Drug|false|false||systemnull|System, LOINC Axis 4|Finding|false|false||system
null|System|Finding|false|false||systemnull|Device system|Device|false|false||system
null|System - kit|Device|false|false||systemnull|System (unit of presentation)|LabModifier|false|false||systemnull|Coronary Vessels|Anatomy|false|false||vessel coronarynull|Vessel Positions|Anatomy|false|false||vessel
null|Blood Vessel|Anatomy|false|false||vesselnull|Vessel (unit of presentation)|LabModifier|false|false||vesselnull|Coronary Artery Disease|Disorder|false|false||coronary artery disease
null|Coronary Arteriosclerosis|Disorder|false|false||coronary artery diseasenull|Coronary artery|Anatomy|false|false||coronary arterynull|Heart|Anatomy|false|false||coronarynull|Coronary|Modifier|false|false||coronarynull|Arteriopathic disease|Disorder|false|false||artery diseasenull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Disease|Disorder|false|false||diseasenull|apparent|Finding|false|false||apparentnull|Flow|Phenomenon|false|false||flownull|Stenosis|Finding|false|false||stenosesnull|Leukocyte adhesion deficiency type 1|Disorder|false|false||LAD
null|Leukocyte adhesion deficiency|Disorder|false|false||LADnull|ITGB2 wt Allele|Finding|false|false||LAD
null|DLD gene|Finding|false|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false||LADnull|Ladino Language|Entity|false|false||LADnull|Stent restenosis|Finding|false|false||stent restenosisnull|null|Device|false|false||stentnull|Restenosis|Finding|false|false||restenosisnull|Junction Device|Device|false|false||junctionnull|Junctional|Modifier|false|false||junctionnull|Old|Time|false|false||oldnull|LDB3 wt Allele|Finding|false|false||Cypher
null|LDB3 gene|Finding|false|false||Cyphernull|null|Device|false|false||stentnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|null|Device|false|false||stentnull|Macromolecular Branch|Drug|false|false||branchnull|Branch of|Modifier|false|false||branchnull|Participation Type - origin|Finding|false|false||origin
null|National origin|Finding|false|false||originnull|Beginning|Time|false|false||originnull|Stenosis|Finding|false|false||stenosisnull|Stenosis <Pimeliinae>|Entity|false|false||stenosisnull|Stenosis Morphology|Modifier|false|false||stenosisnull|Methylcytosine Dioxygenase TET1|Drug|false|false||LCx
null|Methylcytosine Dioxygenase TET1|Drug|false|false||LCxnull|TET1 wt Allele|Finding|false|false||LCx
null|TET1 gene|Finding|false|false||LCxnull|Stenosis|Finding|false|false||stenosisnull|Stenosis <Pimeliinae>|Entity|false|false||stenosisnull|Stenosis Morphology|Modifier|false|false||stenosisnull|Participation Type - origin|Finding|false|false||origin
null|National origin|Finding|false|false||originnull|Beginning|Time|false|false||originnull|Stenosis|Finding|false|false||stenosisnull|Stenosis <Pimeliinae>|Entity|false|false||stenosisnull|Stenosis Morphology|Modifier|false|false||stenosisnull|Macromolecular Branch|Drug|false|false||branchnull|Branch of|Modifier|false|false||branchnull|Stenosis|Finding|false|false||stenosisnull|Stenosis <Pimeliinae>|Entity|false|false||stenosisnull|Stenosis Morphology|Modifier|false|false||stenosisnull|Limited component (foundation metadata concept)|Finding|false|false||Limited
null|Limited (extensiveness)|Finding|false|false||Limitednull|Hemodynamics|Finding|false|false||hemodynamicsnull|hemodynamics (procedure)|Procedure|false|false||hemodynamicsnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Systemic Route of Administration|Finding|false|false||systemic
null|Systemic|Finding|false|false||systemicnull|Arteries|Anatomy|false|false||arterialnull|Arterial|Modifier|false|false||arterialnull|Hypertensive disease|Disorder|false|false||hypertensionnull|Central brand of multivitamin with minerals|Drug|false|false||central
null|Central brand of multivitamin with minerals|Drug|false|false||centralnull|Central Minus|Procedure|false|false||centralnull|Central|Modifier|false|false||centralnull|Aortic Pressure|Lab|false|false||aortic pressurenull|Aorta|Anatomy|false|false||aorticnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|mmHg|LabModifier|false|false||mmHgnull|Success|Finding|false|false||Successfulnull|Successful|Modifier|false|false||Successfulnull|Percutaneous Transluminal Coronary Angioplasty|Procedure|false|false||PTCAnull|Stenting|Procedure|false|false||stentingnull|null|Device|false|false||stentingnull|null|Device|false|false||stentnull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|angiogram|Procedure|false|false||angiographynull|Residual|Modifier|false|false||residualnull|Stenosis|Finding|false|false||stenosisnull|Stenosis <Pimeliinae>|Entity|false|false||stenosisnull|Stenosis Morphology|Modifier|false|false||stenosisnull|apparent|Finding|false|false||apparentnull|Dissecting hemorrhage|Finding|false|false||dissectionnull|Tissue Dissection|Procedure|false|false||dissectionnull|Flow|Phenomenon|false|false||flownull|Vision|Finding|false|false||seenull|See|Event|false|false||seenull|Percutaneous Transluminal Coronary Angioplasty|Procedure|false|false||PTCAnull|Published Comment|Finding|false|false||comments
null|Comment|Finding|false|false||commentsnull|Final diagnosis (discharge)|Modifier|false|false||FINAL DIAGNOSISnull|Diagnosis Type - Final|Finding|false|false||FINALnull|Final|Time|false|false||FINALnull|End-stage|Modifier|false|false||FINALnull|Diagnosis Classification - Diagnosis|Finding|false|false||DIAGNOSIS
null|diagnosis aspects|Finding|false|false||DIAGNOSISnull|Diagnosis|Procedure|false|false||DIAGNOSISnull|null|Attribute|false|false||DIAGNOSISnull|Coronary Vessels|Anatomy|false|false||vessel coronarynull|Vessel Positions|Anatomy|false|false||vessel
null|Blood Vessel|Anatomy|false|false||vesselnull|Vessel (unit of presentation)|LabModifier|false|false||vesselnull|Coronary Artery Disease|Disorder|false|false||coronary artery disease
null|Coronary Arteriosclerosis|Disorder|false|false||coronary artery diseasenull|Coronary artery|Anatomy|false|false||coronary arterynull|Heart|Anatomy|false|false||coronarynull|Coronary|Modifier|false|false||coronarynull|Arteriopathic disease|Disorder|false|false||artery diseasenull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Disease|Disorder|false|false||diseasenull|Success|Finding|false|false||Successfulnull|Successful|Modifier|false|false||Successfulnull|Percutaneous Transluminal Coronary Angioplasty|Procedure|false|false||PTCAnull|Stenting|Procedure|false|false||stentingnull|null|Device|false|false||stentingnull|DES protein, human|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|DES protein, human|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DESnull|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|Disorder|false|false||DESnull|DES gene|Finding|false|false||DESnull|BRIEF Health Literacy Screening Tool|Finding|false|false||Brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||Briefnull|Brief|Time|false|false||Briefnull|Shortened|Modifier|false|false||Briefnull|Hospital course|Finding|false|false||Hospital Coursenull|null|Attribute|false|false||Hospital Coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||Coursenull|Angina, Unstable|Disorder|false|false||Unstable anginanull|Unstable status|Finding|false|false||Unstablenull|Angina Pectoris|Finding|false|false||angina
null|null|Finding|false|false||anginanull|null|Attribute|false|false||anginanull|Description|Finding|false|false||Descriptionnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Somewhat|Finding|false|false||somewhatnull|atypia morphology|Finding|false|false||atypicalnull|Atypical|Modifier|false|false||atypicalnull|Angina Pectoris|Finding|false|false||angina
null|null|Finding|false|false||anginanull|null|Attribute|false|false||anginanull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|Numerous|LabModifier|false|false||multiplenull|Structure of cisterna pontis|Anatomy|false|false||PCIsnull|risk factors - observation list|Finding|false|false||risk factors
null|risk factors|Finding|false|false||risk factors
null|History of - risk factor|Finding|false|false||risk factorsnull|null|Attribute|false|false||risk factorsnull|Risk|Finding|false|false||risknull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Exercise stress test|Procedure|false|false||stress test
null|Stress Test|Procedure|false|false||stress testnull|Stress bismuth subsalicylate|Drug|false|false||stress
null|Stress bismuth subsalicylate|Drug|false|false||stressnull|Stress|Finding|false|false||stressnull|W stress|Attribute|false|false||stressnull|Tests (qualifier value)|Finding|false|false||test
null|Testing|Finding|false|false||testnull|Laboratory Procedures|Procedure|false|false||testnull|Test - temporal region|Anatomy|false|false||testnull|Test Result|Lab|false|false||testnull|Test Dosing Unit|LabModifier|false|false||testnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Nuclear stress test|Procedure|false|false||Nuclear stress testnull|Nuclear (incident type)|Modifier|false|false||Nuclear
null|Nuclear (nucleus)|Modifier|false|false||Nuclearnull|Exercise stress test|Procedure|false|false||stress test
null|Stress Test|Procedure|false|false||stress testnull|Stress bismuth subsalicylate|Drug|false|false||stress
null|Stress bismuth subsalicylate|Drug|false|false||stressnull|Stress|Finding|false|false||stressnull|W stress|Attribute|false|false||stressnull|Tests (qualifier value)|Finding|false|false||test
null|Testing|Finding|false|false||testnull|Laboratory Procedures|Procedure|false|false||testnull|Test - temporal region|Anatomy|false|false||testnull|Test Result|Lab|false|false||testnull|Test Dosing Unit|LabModifier|false|false||testnull|Reversible|Finding|false|false||reversiblenull|Medium (Substance)|Drug|false|false||medium
null|Culture Media|Drug|false|false||mediumnull|A Medium Amount of Time|Finding|false|false||medium
null|Communications Media|Finding|false|false||medium
null|A Medium Amount|Finding|false|false||mediumnull|Message Waiting Priority - Medium|Modifier|false|false||medium
null|medium exposure|Modifier|false|false||mediumnull|Medium|LabModifier|false|false||mediumnull|Moderate (severity modifier)|Modifier|false|false||moderate severitynull|Moderate - Severity of Illness Code|Finding|false|false||moderate
null|Moderate|Finding|false|false||moderatenull|Moderate (severity modifier)|Modifier|false|false||moderate
null|Moderate - Allergy Severity|Modifier|false|false||moderate
null|Moderation|Modifier|false|false||moderatenull|With intensity|Modifier|false|false||severity
null|Severities|Modifier|false|false||severitynull|Perfusion (biological)|Finding|false|false||perfusion
null|Perfusion route|Finding|false|false||perfusionnull|Chemotherapeutic Perfusion|Procedure|false|false||perfusion
null|Perfusion (procedure)|Procedure|false|false||perfusionnull|THYROID HORMONE PLASMA MEMBRANE TRANSPORT DEFECT|Disorder|false|false||defectnull|Defect|Finding|false|false||defectnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Circumflex|Modifier|false|false||circumflexnull|Territory|Entity|false|false||territory
null|Geographic state|Entity|false|false||territorynull|TNFSF14 protein, human|Drug|false|false||light
null|TNFSF14 protein, human|Drug|false|false||lightnull|Light - subjective measurement|Finding|false|false||light
null|TNFSF14 wt Allele|Finding|false|false||light
null|TNFSF14 gene|Finding|false|false||light
null|Light color|Finding|false|false||lightnull|Phototherapy|Procedure|false|false||lightnull|Light|Phenomenon|false|false||lightnull|Light (qualifier)|Modifier|false|false||lightnull|Exercise stress test|Procedure|false|false||stress test
null|Stress Test|Procedure|false|false||stress testnull|Stress bismuth subsalicylate|Drug|false|false||stress
null|Stress bismuth subsalicylate|Drug|false|false||stressnull|Stress|Finding|false|false||stressnull|W stress|Attribute|false|false||stressnull|Tests (qualifier value)|Finding|false|false||test
null|Testing|Finding|false|false||testnull|Laboratory Procedures|Procedure|false|false||testnull|Test - temporal region|Anatomy|false|false||testnull|Test Result|Lab|false|false||testnull|Test Dosing Unit|LabModifier|false|false||testnull|findings aspects|Finding|false|false||findingsnull|null|Attribute|false|false||findingsnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Cardiac attachment|Finding|false|false||cardiacnull|Heart|Anatomy|false|false||cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||cardiacnull|Catheterization|Procedure|false|false||catheterizationnull|null|Time|false|false||Prior tonull|null|Time|false|false||Priornull|Cardiac catheterisation as the cause of abnormal reaction of the patient, or of later complication, without mention of misadventure at the time of the procedure|Disorder|false|false||cardiac catheterizationnull|Diagnostic Service Section ID - Cardiac Catheterization|Finding|false|false||cardiac catheterizationnull|Consent Type - Cardiac Catheterization|Procedure|false|false||cardiac catheterization
null|Cardiac Catheterization Procedures|Procedure|false|false||cardiac catheterizationnull|Cardiac attachment|Finding|false|false||cardiacnull|Heart|Anatomy|false|false||cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||cardiacnull|Catheterization|Procedure|false|false||catheterizationnull|Acute kidney injury|Disorder|false|false||acute kidney injury
null|Kidney Failure, Acute|Disorder|false|false||acute kidney injurynull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Injury of kidney|Disorder|false|false||kidney injurynull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false||kidney
null|Benign neoplasm of kidney|Disorder|false|false||kidneynull|Kidney problem|Finding|false|false||kidneynull|examination of kidney|Procedure|false|false||kidney
null|Procedures on Kidney|Procedure|false|false||kidneynull|Kidney|Anatomy|false|false||kidney
null|Both kidneys|Anatomy|false|false||kidneynull|Traumatic AND/OR non-traumatic injury|Disorder|false|false||injury
null|Traumatic injury|Disorder|false|false||injurynull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Pharmaceutical Preparations|Drug|false|false||drug
null|Pharmacologic Substance|Drug|false|false||drugnull|Drug problem|Finding|false|false||drugnull|null|Device|false|false||stentnull|Obtuse|Modifier|false|false||obtusenull|Target Awareness - marginal|Finding|false|false||marginalnull|Marginal (quality)|Modifier|false|false||marginal
null|Marginal|Modifier|false|false||marginalnull|Macromolecular Branch|Drug|false|false||branchnull|Branch of|Modifier|false|false||branchnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Hypertensive (finding)|Finding|false|false||hypertensivenull|Cardiac attachment|Finding|false|false||cardiacnull|Heart|Anatomy|false|false||cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||cardiacnull|Catheterization|Procedure|false|false||catheterizationnull|nitroglycerin|Drug|false|false||nitroglycerin
null|nitroglycerin|Drug|false|false||nitroglycerinnull|Discussion (communication)|Finding|false|false||discussionnull|Discussion (procedure)|Procedure|false|false||discussionnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|aspirin|Drug|false|false||aspirin
null|aspirin|Drug|false|false||aspirinnull|Full|Modifier|false|false||fullnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Plavix|Drug|false|false||plavix
null|Plavix|Drug|false|false||plavixnull|metoprolol|Drug|false|false||metoprolol
null|metoprolol|Drug|false|false||metoprololnull|Imdur|Drug|false|false||imdur
null|Imdur|Drug|false|false||imdurnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|atorvastatin|Drug|false|false||atorvastatin
null|atorvastatin|Drug|false|false||atorvastatinnull|Evidence of (contextual qualifier)|Finding|false|false||evidence ofnull|Evidence|Finding|false|false||evidencenull|Coronary Artery Disease|Disorder|false|false||coronary artery disease
null|Coronary Arteriosclerosis|Disorder|false|false||coronary artery diseasenull|Coronary artery|Anatomy|false|false||coronary arterynull|Heart|Anatomy|false|false||coronarynull|Coronary|Modifier|false|false||coronarynull|Arteriopathic disease|Disorder|false|false||artery diseasenull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Disease|Disorder|false|false||diseasenull|Periodicals|Finding|false|false||Serialnull|Serial|Time|false|false||Serialnull|Cardiac enzymes|Drug|false|false||cardiac enzymes
null|Cardiac enzymes|Drug|false|false||cardiac enzymesnull|Cardiac enzymes/isoenzymes measurement|Procedure|false|false||cardiac enzymesnull|null|Attribute|false|false||cardiac enzymesnull|Cardiac attachment|Finding|false|false||cardiacnull|Heart|Anatomy|false|false||cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||cardiacnull|Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM|Drug|false|false||enzymes
null|Enzymes, peripheral vasodilators|Drug|false|false||enzymes
null|Enzymes, peripheral vasodilators|Drug|false|false||enzymes
null|Enzymes, peripheral vasodilators|Drug|false|false||enzymes
null|Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM|Drug|false|false||enzymes
null|Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM|Drug|false|false||enzymes
null|Enzymes, antithrombotic|Drug|false|false||enzymes
null|Enzymes, antithrombotic|Drug|false|false||enzymes
null|Enzymes, antithrombotic|Drug|false|false||enzymes
null|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS|Drug|false|false||enzymes
null|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS|Drug|false|false||enzymes
null|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS|Drug|false|false||enzymes
null|Enzymes, hematological|Drug|false|false||enzymes
null|Enzymes, hematological|Drug|false|false||enzymes
null|Enzymes, hematological|Drug|false|false||enzymes
null|Enzymes|Drug|false|false||enzymes
null|Enzymes|Drug|false|false||enzymes
null|Enzymes for ALIMENTARY TRACT AND METABOLISM|Drug|false|false||enzymes
null|Enzymes for ALIMENTARY TRACT AND METABOLISM|Drug|false|false||enzymes
null|Enzymes for ALIMENTARY TRACT AND METABOLISM|Drug|false|false||enzymesnull|enzymology|Finding|false|false||enzymesnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Referral category - Outpatient|Finding|false|false||OUTPATIENT
null|Patient Class - Outpatient|Finding|false|false||OUTPATIENTnull|Outpatients|Subject|false|false||OUTPATIENTnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|aspirin|Drug|false|false||aspirin
null|aspirin|Drug|false|false||aspirinnull|Plavix|Drug|false|false||plavix
null|Plavix|Drug|false|false||plavixnull|Daily|Time|false|false||dailynull|next - HtmlLinkType|Finding|false|false||nextnull|Following|Time|false|false||next
null|Then|Time|false|false||nextnull|Adjacent|Modifier|false|false||nextnull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Cardiovascular system|Anatomy|false|false||cardiologynull|cardiology (field)|Title|false|false||cardiologynull|Cardiology service|Entity|false|false||cardiologynull|Follow-up status|Finding|false|false||follow-upnull|follow-up|Procedure|false|false||follow-upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Group Specimen|Finding|false|false||group
null|Stage Grouping|Finding|false|false||group
null|Group Object|Finding|false|false||group
null|Groups|Finding|false|false||groupnull|Population Group|Subject|false|false||group
null|Social group|Subject|false|false||group
null|User Group|Subject|false|false||groupnull|Acute kidney injury|Disorder|false|false||Acute kidney injury
null|Kidney Failure, Acute|Disorder|false|false||Acute kidney injurynull|Admission Level of Care Code - Acute|Finding|false|false||Acute
null|Acute - Triage Code|Finding|false|false||Acutenull|acute|Time|false|false||Acutenull|Injury of kidney|Disorder|false|false||kidney injurynull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false||kidney
null|Benign neoplasm of kidney|Disorder|false|false||kidneynull|Kidney problem|Finding|false|false||kidneynull|examination of kidney|Procedure|false|false||kidney
null|Procedures on Kidney|Procedure|false|false||kidneynull|Kidney|Anatomy|false|false||kidney
null|Both kidneys|Anatomy|false|false||kidneynull|Traumatic AND/OR non-traumatic injury|Disorder|false|false||injury
null|Traumatic injury|Disorder|false|false||injurynull|creatinine|Drug|false|false||Creatinine
null|creatinine|Drug|false|false||Creatininenull|Creatinine metabolic function|Finding|false|false||Creatininenull|Creatinine measurement|Procedure|false|false||Creatininenull|Current (present time)|Time|false|false||currentlynull|Renal function|Finding|false|false||Renal functionnull|Kidney Function Tests|Procedure|false|false||Renal functionnull|Urologic Diseases|Disorder|false|false||Renalnull|Kidney|Anatomy|false|false||Renalnull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|lisinopril|Drug|false|false||lisinopril
null|lisinopril|Drug|false|false||lisinoprilnull|furosemide|Drug|false|false||furosemide
null|furosemide|Drug|false|false||furosemidenull|ACOT8 gene|Finding|false|false||htenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|furosemide|Drug|false|false||furosemide
null|furosemide|Drug|false|false||furosemidenull|Approximate|Modifier|false|false||approximatelynull|month|Time|false|false||monthsnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|Growth and Development function|Finding|false|false||development
null|development aspects|Finding|false|false||development
null|biological development|Finding|false|false||development
null|Development|Finding|false|false||developmentnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Serum creatinine raised|Finding|false|false||elevated serum creatininenull|Elevated|Modifier|false|false||elevated
null|High|Modifier|false|false||elevatednull|Serum creatinine level|Finding|false|false||serum creatininenull|Creatinine measurement, serum (procedure)|Procedure|false|false||serum creatininenull|Cell Culture Serum|Drug|false|false||serumnull|Serum specimen|Finding|false|false||serum
null|null|Finding|false|false||serum
null|Serum|Finding|false|false||serumnull|creatinine|Drug|false|false||creatinine
null|creatinine|Drug|false|false||creatininenull|Creatinine metabolic function|Finding|false|false||creatininenull|Creatinine measurement|Procedure|false|false||creatininenull|Serum creatinine level|Finding|false|false||Serum creatininenull|Creatinine measurement, serum (procedure)|Procedure|false|false||Serum creatininenull|Cell Culture Serum|Drug|false|false||Serumnull|Serum specimen|Finding|false|false||Serum
null|null|Finding|false|false||Serum
null|Serum|Finding|false|false||Serumnull|creatinine|Drug|false|false||creatinine
null|creatinine|Drug|false|false||creatininenull|Creatinine metabolic function|Finding|false|false||creatininenull|Creatinine measurement|Procedure|false|false||creatininenull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|lisinopril|Drug|false|false||lisinopril
null|lisinopril|Drug|false|false||lisinoprilnull|Serum creatinine level|Finding|false|false||serum creatininenull|Creatinine measurement, serum (procedure)|Procedure|false|false||serum creatininenull|Cell Culture Serum|Drug|false|false||serumnull|Serum specimen|Finding|false|false||serum
null|null|Finding|false|false||serum
null|Serum|Finding|false|false||serumnull|creatinine|Drug|false|false||creatinine
null|creatinine|Drug|false|false||creatininenull|Creatinine metabolic function|Finding|false|false||creatininenull|Creatinine measurement|Procedure|false|false||creatininenull|Instructions|Finding|false|false||instructions
null|Instruction [Publication Type]|Finding|false|false||instructionsnull|null|Attribute|false|false||instructionsnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Follow-up status|Finding|false|false||follow-upnull|follow-up|Procedure|false|false||follow-upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|Primary Care Physicians|Subject|false|false||primary care physician
null|Primary care provider|Subject|false|false||primary care physiciannull|Location Service Code - Primary Care|Finding|false|false||primary carenull|Primary Health Care|Procedure|false|false||primary carenull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|null|Attribute|false|false||physiciannull|Physicians|Subject|false|false||physiciannull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Basic metabolic panel|Procedure|false|false||basic metabolic panelnull|Base|Drug|false|false||basicnull|Basis - conceptual entity|Finding|false|false||basicnull|Basic (cigarettes)|Device|false|false||basicnull|Metabolic Process, Cellular|Finding|false|false||metabolic
null|Metabolic|Finding|false|false||metabolicnull|Multisection metabolic|Procedure|false|false||metabolicnull|Groups|Finding|false|false||panelnull|Panel Device|Device|false|false||panelnull|Heart Failure, Diastolic|Disorder|false|false||Diastolic heart failurenull|Diastole|Attribute|false|false||Diastolicnull|Congestive heart failure|Disorder|false|false||heart failure
null|Heart failure|Disorder|false|false||heart failurenull|Malignant neoplasm of heart|Disorder|false|false||heart
null|benign neoplasm of heart|Disorder|false|false||heartnull|HEART PROBLEM|Finding|false|false||heartnull|Chest>Heart|Anatomy|false|false||heart
null|Heart|Anatomy|false|false||heartnull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Lasix|Drug|false|false||lasix
null|Lasix|Drug|false|false||lasixnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Acute kidney injury|Disorder|false|false||acute kidney injury
null|Kidney Failure, Acute|Disorder|false|false||acute kidney injurynull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Injury of kidney|Disorder|false|false||kidney injurynull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false||kidney
null|Benign neoplasm of kidney|Disorder|false|false||kidneynull|Kidney problem|Finding|false|false||kidneynull|examination of kidney|Procedure|false|false||kidney
null|Procedures on Kidney|Procedure|false|false||kidneynull|Kidney|Anatomy|false|false||kidney
null|Both kidneys|Anatomy|false|false||kidneynull|Traumatic AND/OR non-traumatic injury|Disorder|false|false||injury
null|Traumatic injury|Disorder|false|false||injurynull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Primary Care Physicians|Subject|false|false||primary care physician
null|Primary care provider|Subject|false|false||primary care physiciannull|Location Service Code - Primary Care|Finding|false|false||primary carenull|Primary Health Care|Procedure|false|false||primary carenull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|null|Attribute|false|false||physiciannull|Physicians|Subject|false|false||physiciannull|Lasix|Drug|false|false||lasix
null|Lasix|Drug|false|false||lasixnull|Referral category - Outpatient|Finding|false|false||OUTPATIENT
null|Patient Class - Outpatient|Finding|false|false||OUTPATIENTnull|Outpatients|Subject|false|false||OUTPATIENTnull|Referral category - Outpatient|Finding|false|false||Outpatient
null|Patient Class - Outpatient|Finding|false|false||Outpatientnull|Outpatients|Subject|false|false||Outpatientnull|Bone Morphogenetic Proteins|Drug|false|false||BMP
null|Bone Morphogenetic Proteins|Drug|false|false||BMPnull|carmustine/methotrexate/procarbazine protocol|Procedure|false|false||BMPnull|Preventive monitoring|Procedure|false|false||monitoringnull|null|Event|false|false||monitoringnull|Cell Culture Serum|Drug|false|false||serumnull|Serum specimen|Finding|false|false||serum
null|null|Finding|false|false||serum
null|Serum|Finding|false|false||serumnull|creatinine|Drug|false|false||creatinine
null|creatinine|Drug|false|false||creatininenull|Creatinine metabolic function|Finding|false|false||creatininenull|Creatinine measurement|Procedure|false|false||creatininenull|Lasix|Drug|false|false||lasix
null|Lasix|Drug|false|false||lasixnull|Location Service Code - Primary Care|Finding|false|false||primary carenull|Primary Health Care|Procedure|false|false||primary carenull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|Continuity Assessment Record and Evaluation|Finding|false|false||care
null|In care (finding)|Finding|false|false||carenull|care activity|Event|false|false||carenull|null|Attribute|false|false||physiciannull|Physicians|Subject|false|false||physiciannull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Type 2 Diabetesnull|Type 2|Finding|false|false||Type 2null|Type - ParameterizedDataType|Finding|false|false||Type
null|SGCG gene|Finding|false|false||Typenull|null|Modifier|false|false||Typenull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Diabetes
null|Diabetes|Disorder|false|false||Diabetes
null|Diabetes Mellitus|Disorder|false|false||Diabetesnull|insulin, regular, human|Drug|false|false||insulin
null|Insulin [EPC]|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulinnull|INS gene|Finding|false|false||insulinnull|Insulin measurement|Procedure|false|false||insulinnull|dependent|Finding|false|false||dependentnull|Dependent - ability|Modifier|false|false||dependent
null|Conditional|Modifier|false|false||dependentnull|Moderate Response|Finding|false|false||Moderately
null|Moderate|Finding|false|false||Moderately
null|Moderate Effect|Finding|false|false||Moderatelynull|Moderate (severity modifier)|Modifier|false|false||Moderately
null|Moderation|Modifier|false|false||Moderatelynull|Last|Modifier|false|false||lastnull|United States Military enlisted E3 (qualifier value)|Finding|false|false||A1cnull|Hemoglobin A1c measurement|Procedure|false|false||A1cnull|Lantus|Drug|false|false||Lantus
null|Lantus|Drug|false|false||Lantusnull|Sliding|Finding|false|false||slidingnull|Scale, LOINC Axis 5|Finding|false|false||scale
null|Base Number|Finding|false|false||scale
null|Scale - rank|Finding|false|false||scalenull|Integumentary scale|Anatomy|false|false||scalenull|Weight measurement scales|Device|false|false||scalenull|Scaling|Event|false|false||scalenull|Hospitalization|Procedure|false|false||hospitalizationnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Dosage|LabModifier|false|false||dosesnull|Lantus|Drug|false|false||lantus
null|Lantus|Drug|false|false||lantusnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|insulin, regular, human|Drug|false|false||insulin
null|Insulin [EPC]|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulinnull|INS gene|Finding|false|false||insulinnull|Insulin measurement|Procedure|false|false||insulinnull|Scale, LOINC Axis 5|Finding|false|false||scale
null|Base Number|Finding|false|false||scale
null|Scale - rank|Finding|false|false||scalenull|Integumentary scale|Anatomy|false|false||scalenull|Weight measurement scales|Device|false|false||scalenull|Scaling|Event|false|false||scalenull|Hypertensive disease|Disorder|false|false||Hypertensionnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Blood pressure finding|Finding|false|false||blood pressure
null|Systemic arterial pressure|Finding|false|false||blood pressure
null|Blood Pressure|Finding|false|false||blood pressurenull|Blood pressure determination|Procedure|false|false||blood pressurenull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|objective (goal)|Finding|false|false||goal
null|Act Mood - Goal|Finding|false|false||goalnull|Continuous|Finding|false|false||continuednull|metoprolol|Drug|false|false||metoprolol
null|metoprolol|Drug|false|false||metoprololnull|Imdur|Drug|false|false||imdur
null|Imdur|Drug|false|false||imdurnull|furosemide|Drug|false|false||furosemide
null|furosemide|Drug|false|false||furosemidenull|lisinopril|Drug|false|false||lisinopril
null|lisinopril|Drug|false|false||lisinoprilnull|TNFSF14 protein, human|Drug|false|false||light
null|TNFSF14 protein, human|Drug|false|false||lightnull|Light - subjective measurement|Finding|false|false||light
null|TNFSF14 wt Allele|Finding|false|false||light
null|TNFSF14 gene|Finding|false|false||light
null|Light color|Finding|false|false||lightnull|Phototherapy|Procedure|false|false||lightnull|Light|Phenomenon|false|false||lightnull|Light (qualifier)|Modifier|false|false||lightnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Elevated|Modifier|false|false||elevated
null|High|Modifier|false|false||elevatednull|Serum creatinine level|Finding|false|false||serum creatininenull|Creatinine measurement, serum (procedure)|Procedure|false|false||serum creatininenull|Cell Culture Serum|Drug|false|false||serumnull|Serum specimen|Finding|false|false||serum
null|null|Finding|false|false||serum
null|Serum|Finding|false|false||serumnull|creatinine|Drug|false|false||creatinine
null|creatinine|Drug|false|false||creatininenull|Creatinine metabolic function|Finding|false|false||creatininenull|Creatinine measurement|Procedure|false|false||creatininenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Cardiac attachment|Finding|false|false||cardiacnull|Heart|Anatomy|false|false||cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||cardiacnull|Catheterization|Procedure|false|false||catheterizationnull|Elevated|Modifier|false|false||elevated
null|High|Modifier|false|false||elevatednull|Systole|Finding|false|false||systolicnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Pressure (finding)|Finding|false|false||pressuresnull|null|Phenomenon|false|false||pressuresnull|nitroglycerin|Drug|false|false||nitroglycerin
null|nitroglycerin|Drug|false|false||nitroglycerinnull|Control brand of phenylpropanolamine|Drug|false|false||control
null|CONTROL veterinary product|Drug|false|false||control
null|control substance|Drug|false|false||control
null|Control brand of phenylpropanolamine|Drug|false|false||controlnull|Control - Relationship modifier|Finding|false|false||control
null|Control function|Finding|false|false||control
null|Scientific Control|Finding|false|false||controlnull|Control Groups|Subject|false|false||controlnull|True Control Status|Modifier|false|false||control
null|control aspects|Modifier|false|false||controlnull|Systemic arterial pressure|Finding|false|false||blood pressuresnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Pressure (finding)|Finding|false|false||pressuresnull|null|Phenomenon|false|false||pressuresnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|nitroglycerin|Drug|false|false||nitroglycerin
null|nitroglycerin|Drug|false|false||nitroglycerinnull|4 Hours|Time|false|false||4 hoursnull|Hour|Time|false|false||hoursnull|Cardiac catheterisation as the cause of abnormal reaction of the patient, or of later complication, without mention of misadventure at the time of the procedure|Disorder|false|false||cardiac catheterizationnull|Diagnostic Service Section ID - Cardiac Catheterization|Finding|false|false||cardiac catheterizationnull|Consent Type - Cardiac Catheterization|Procedure|false|false||cardiac catheterization
null|Cardiac Catheterization Procedures|Procedure|false|false||cardiac catheterizationnull|Cardiac attachment|Finding|false|false||cardiacnull|Heart|Anatomy|false|false||cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||cardiacnull|Catheterization|Procedure|false|false||catheterizationnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|lisinopril|Drug|false|false||lisinopril
null|lisinopril|Drug|false|false||lisinoprilnull|Cell Culture Serum|Drug|false|false||serumnull|Serum specimen|Finding|false|false||serum
null|null|Finding|false|false||serum
null|Serum|Finding|false|false||serumnull|creatinine|Drug|false|false||creatinine
null|creatinine|Drug|false|false||creatininenull|Creatinine metabolic function|Finding|false|false||creatininenull|Creatinine measurement|Procedure|false|false||creatininenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|next - HtmlLinkType|Finding|false|false||nextnull|Following|Time|false|false||next
null|Then|Time|false|false||nextnull|Adjacent|Modifier|false|false||nextnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Referral category - Outpatient|Finding|false|false||OUTPATIENT
null|Patient Class - Outpatient|Finding|false|false||OUTPATIENTnull|Outpatients|Subject|false|false||OUTPATIENTnull|Primary Care Physicians|Subject|false|false||primary care physician
null|Primary care provider|Subject|false|false||primary care physiciannull|Location Service Code - Primary Care|Finding|false|false||primary carenull|Primary Health Care|Procedure|false|false||primary carenull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|null|Attribute|false|false||physiciannull|Physicians|Subject|false|false||physiciannull|History of recent hospitalization|Finding|false|false||recent hospitalizationnull|Recent|Time|false|false||recentnull|Hospitalization|Procedure|false|false||hospitalizationnull|Antihypertensive Agents|Drug|false|false||anti-hypertensivenull|GDC Regimen Terminology|Finding|false|false||regimennull|Treatment Protocols|Procedure|false|false||regimennull|TNFSF14 protein, human|Drug|false|false||light
null|TNFSF14 protein, human|Drug|false|false||lightnull|Light - subjective measurement|Finding|false|false||light
null|TNFSF14 wt Allele|Finding|false|false||light
null|TNFSF14 gene|Finding|false|false||light
null|Light color|Finding|false|false||lightnull|Phototherapy|Procedure|false|false||lightnull|Light|Phenomenon|false|false||lightnull|Light (qualifier)|Modifier|false|false||lightnull|Serum creatinine raised|Finding|false|false||elevated serum creatininenull|Elevated|Modifier|false|false||elevated
null|High|Modifier|false|false||elevatednull|Serum creatinine level|Finding|false|false||serum creatininenull|Creatinine measurement, serum (procedure)|Procedure|false|false||serum creatininenull|Cell Culture Serum|Drug|false|false||serumnull|Serum specimen|Finding|false|false||serum
null|null|Finding|false|false||serum
null|Serum|Finding|false|false||serumnull|creatinine|Drug|false|false||creatinine
null|creatinine|Drug|false|false||creatininenull|Creatinine metabolic function|Finding|false|false||creatininenull|Creatinine measurement|Procedure|false|false||creatininenull|Hyperlipidemia|Disorder|false|false||Hyperlipidemia
null|Hyperlipoproteinemias|Disorder|false|false||Hyperlipidemianull|Serum lipids high (finding)|Finding|false|false||Hyperlipidemianull|Well (answer to question)|Finding|false|false||Wellnull|Well (container)|Device|false|false||Wellnull|Microplate Well|Modifier|false|false||Well
null|Good|Modifier|false|false||Well
null|Healthy|Modifier|false|false||Wellnull|Last|Modifier|false|false||lastnull|Low-Density Lipoproteins|Drug|false|false||LDL
null|Low-Density Lipoproteins|Drug|false|false||LDLnull|Low density lipoprotein cholesterol measurement|Procedure|false|false||LDLnull|objective (goal)|Finding|false|false||goal
null|Act Mood - Goal|Finding|false|false||goalnull|Low-Density Lipoproteins|Drug|false|false||LDL
null|Low-Density Lipoproteins|Drug|false|false||LDLnull|Low density lipoprotein cholesterol measurement|Procedure|false|false||LDLnull|Triglycerides|Drug|false|false||triglycerides
null|Triglycerides|Drug|false|false||triglyceridesnull|Triglycerides metabolic function|Finding|false|false||triglyceridesnull|Triglycerides measurement|Procedure|false|false||triglyceridesnull|MILDLY|Modifier|false|false||mildly
null|Mild (qualifier value)|Modifier|false|false||mildlynull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|Daily|Time|false|false||dailynull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Lesion|Finding|false|false||lesionsnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Fasting lipid profile|Procedure|false|false||fasting lipid panelnull|Fasting|Finding|false|false||fastingnull|Fasting (regime/therapy)|Procedure|false|false||fastingnull|Lipid panel|Procedure|false|false||lipid panel
null|null|Procedure|false|false||lipid panelnull|null|Attribute|false|false||lipid panelnull|Lipids|Drug|false|false||lipidnull|Groups|Finding|false|false||panelnull|Panel Device|Device|false|false||panelnull|Pending - Allergy Clinical Status|Finding|false|false||pending
null|Pending - referral status|Finding|false|false||pendingnull|Pending - status|Time|false|false||pendingnull|pending - ManagedParticipationStatus|Modifier|false|false||pending
null|pending - RoleStatus|Modifier|false|false||pending
null|Pending - Day type|Modifier|false|false||pendingnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Referral category - Outpatient|Finding|false|false||OUTPATIENT
null|Patient Class - Outpatient|Finding|false|false||OUTPATIENTnull|Outpatients|Subject|false|false||OUTPATIENTnull|Pending - Allergy Clinical Status|Finding|false|false||pending
null|Pending - referral status|Finding|false|false||pendingnull|Pending - status|Time|false|false||pendingnull|pending - ManagedParticipationStatus|Modifier|false|false||pending
null|pending - RoleStatus|Modifier|false|false||pending
null|Pending - Day type|Modifier|false|false||pendingnull|Fasting lipid profile|Procedure|false|false||fasting lipid panelnull|Fasting|Finding|false|false||fastingnull|Fasting (regime/therapy)|Procedure|false|false||fastingnull|Lipid panel|Procedure|false|false||lipid panel
null|null|Procedure|false|false||lipid panelnull|null|Attribute|false|false||lipid panelnull|Lipids|Drug|false|false||lipidnull|Groups|Finding|false|false||panelnull|Panel Device|Device|false|false||panelnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Current (present time)|Time|false|false||Currentlynull|Asymptomatic diagnosis of|Finding|false|false||asymptomatic
null|Asymptomatic (finding)|Finding|false|false||asymptomaticnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|fluticasone|Drug|false|false||fluticasone
null|fluticasone|Drug|false|false||fluticasonenull|albuterol|Drug|false|false||albuterol
null|albuterol|Drug|false|false||albuterolnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|clopidogrel|Drug|false|false||Clopidogrel
null|clopidogrel|Drug|false|false||Clopidogrelnull|Daily|Time|false|false||dailynull|Daily|Time|false|false||dailynull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|Daily|Time|false|false||dailynull|lisinopril|Drug|false|false||Lisinopril
null|lisinopril|Drug|false|false||Lisinoprilnull|Daily|Time|false|false||dailynull|metoprolol succinate|Drug|false|false||Metoprolol succinate
null|metoprolol succinate|Drug|false|false||Metoprolol succinatenull|metoprolol|Drug|false|false||Metoprolol
null|metoprolol|Drug|false|false||Metoprololnull|succinate|Drug|false|false||succinate
null|Succinates|Drug|false|false||succinatenull|Daily|Time|false|false||dailynull|isosorbide mononitrate|Drug|false|false||Isosorbide mononitrate
null|isosorbide mononitrate|Drug|false|false||Isosorbide mononitratenull|isosorbide|Drug|false|false||Isosorbide
null|isosorbide|Drug|false|false||Isosorbidenull|Daily|Time|false|false||dailynull|furosemide|Drug|false|false||Furosemide
null|furosemide|Drug|false|false||Furosemidenull|Daily|Time|false|false||dailynull|nitroglycerin|Drug|false|false||Nitroglycerin
null|nitroglycerin|Drug|false|false||Nitroglycerinnull|CIAO3 gene|Finding|false|false||prnnull|As required|Time|false|false||prn
null|Pro Re Nata|Time|false|false||prnnull|insulin glargine|Drug|false|false||Glargine insulin
null|insulin glargine|Drug|false|false||Glargine insulin
null|insulin glargine|Drug|false|false||Glargine insulinnull|insulin glargine|Drug|false|false||Glargine
null|insulin glargine|Drug|false|false||Glargine
null|insulin glargine|Drug|false|false||Glarginenull|insulin, regular, human|Drug|false|false||insulin
null|Insulin [EPC]|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulinnull|INS gene|Finding|false|false||insulinnull|Insulin measurement|Procedure|false|false||insulinnull|Unit - NCI Thesaurus Property|LabModifier|false|false||units
null|Unit of Measure|LabModifier|false|false||units
null|Unit|LabModifier|false|false||unitsnull|Once a day, at bedtime|Time|false|false||QHSnull|insulin lispro|Drug|false|false||Lispro insulin
null|insulin lispro|Drug|false|false||Lispro insulin
null|insulin lispro|Drug|false|false||Lispro insulinnull|insulin lispro|Drug|false|false||Lispro
null|insulin lispro|Drug|false|false||Lispro
null|insulin lispro|Drug|false|false||Lispronull|insulin, regular, human|Drug|false|false||insulin
null|Insulin [EPC]|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulinnull|INS gene|Finding|false|false||insulinnull|Insulin measurement|Procedure|false|false||insulinnull|Scale, LOINC Axis 5|Finding|false|false||scale
null|Base Number|Finding|false|false||scale
null|Scale - rank|Finding|false|false||scalenull|Integumentary scale|Anatomy|false|false||scalenull|Weight measurement scales|Device|false|false||scalenull|Scaling|Event|false|false||scalenull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|microgram|LabModifier|false|false||mcgnull|Puff Dosing Unit|LabModifier|false|false||puffsnull|HGS protein, human|Drug|false|false||hrs
null|HGS protein, human|Drug|false|false||hrsnull|Dentatorubral-Pallidoluysian Atrophy|Disorder|false|false||hrsnull|HARS1 wt Allele|Finding|false|false||hrs
null|HARS1 gene|Finding|false|false||hrs
null|HGS wt Allele|Finding|false|false||hrs
null|HGS gene|Finding|false|false||hrs
null|ATN1 wt Allele|Finding|false|false||hrs
null|SRSF5 gene|Finding|false|false||hrsnull|Hour|Time|false|false||hrsnull|CIAO3 gene|Finding|false|false||prnnull|As required|Time|false|false||prn
null|Pro Re Nata|Time|false|false||prnnull|fluticasone|Drug|false|false||Fluticasone
null|fluticasone|Drug|false|false||Fluticasonenull|microgram|LabModifier|false|false||mcgnull|Puff Dosing Unit|LabModifier|false|false||puffsnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|pantoprazole|Drug|false|false||Pantoprazole
null|pantoprazole|Drug|false|false||Pantoprazolenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|CIAO3 gene|Finding|false|false||prnnull|As required|Time|false|false||prn
null|Pro Re Nata|Time|false|false||prnnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|potassium chloride|Drug|false|false||Potassium chloride
null|potassium chloride|Drug|false|false||Potassium chloridenull|Potassium Drug Class|Drug|false|false||Potassium
null|Dietary Potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassiumnull|Potassium metabolic function|Finding|false|false||Potassiumnull|Potassium measurement|Procedure|false|false||Potassiumnull|chloride ion|Drug|false|false||chloride
null|Chlorides|Drug|false|false||chloridenull|Chloride metabolic function|Finding|false|false||chloridenull|Chloride measurement|Procedure|false|false||chloridenull|mEq|LabModifier|false|false||mEqnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|cholecalciferol|Drug|false|false||Cholecalciferol
null|cholecalciferol|Drug|false|false||Cholecalciferol
null|cholecalciferol|Drug|false|false||Cholecalciferolnull|Storage Unit|Device|false|false||unit
null|Unit device|Device|false|false||unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||unit
null|Unit of Measure|LabModifier|false|false||unit
null|Unit|LabModifier|false|false||unit
null|Enzyme Unit|LabModifier|false|false||unitnull|Daily|Time|false|false||dailynull|metronidazole|Drug|false|false||Metronidazole
null|metronidazole|Drug|false|false||Metronidazolenull|Lotion|Drug|false|false||lotionnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|clopidogrel|Drug|false|false||clopidogrel
null|clopidogrel|Drug|false|false||clopidogrelnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|aspirin|Drug|false|false||aspirin
null|aspirin|Drug|false|false||aspirinnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|atorvastatin|Drug|false|false||atorvastatin
null|atorvastatin|Drug|false|false||atorvastatinnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|metoprolol succinate|Drug|false|false||metoprolol succinate
null|metoprolol succinate|Drug|false|false||metoprolol succinatenull|metoprolol|Drug|false|false||metoprolol
null|metoprolol|Drug|false|false||metoprololnull|succinate|Drug|false|false||succinate
null|Succinates|Drug|false|false||succinatenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|isosorbide mononitrate|Drug|false|false||isosorbide mononitrate
null|isosorbide mononitrate|Drug|false|false||isosorbide mononitratenull|isosorbide|Drug|false|false||isosorbide
null|isosorbide|Drug|false|false||isosorbidenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|nitroglycerin|Drug|false|false||nitroglycerin
null|nitroglycerin|Drug|false|false||nitroglycerinnull|Sublingual Tablet|Drug|false|false||Tablet, Sublingualnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Sublingual Route of Administration|Finding|false|false||Sublingual
null|Sublingual (intended site)|Finding|false|false||Sublingualnull|Sublingual location|Modifier|false|false||Sublingualnull|Receptors, Antigen, B-Cell|Drug|false|false||Sig
null|Receptors, Antigen, B-Cell|Drug|false|false||Signull|Receptors, Antigen, B-Cell|Finding|false|false||Signull|Short insular gyrus|Anatomy|false|false||Signull|Surveillance Implementation Group|Entity|false|false||Sig
null|Staphylococcus intermedius group|Entity|false|false||Signull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Sublingual Route of Administration|Finding|false|false||Sublingual
null|Sublingual (intended site)|Finding|false|false||Sublingualnull|Sublingual location|Modifier|false|false||Sublingualnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|insulin glargine|Drug|false|false||insulin glargine
null|insulin glargine|Drug|false|false||insulin glargine
null|insulin glargine|Drug|false|false||insulin glarginenull|insulin, regular, human|Drug|false|false||insulin
null|Insulin [EPC]|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulinnull|INS gene|Finding|false|false||insulinnull|Insulin measurement|Procedure|false|false||insulinnull|insulin glargine|Drug|false|false||glargine
null|insulin glargine|Drug|false|false||glargine
null|insulin glargine|Drug|false|false||glarginenull|Unit per Milliliter|LabModifier|false|false||unit/mLnull|Storage Unit|Device|false|false||unit
null|Unit device|Device|false|false||unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||unit
null|Unit of Measure|LabModifier|false|false||unit
null|Unit|LabModifier|false|false||unit
null|Enzyme Unit|LabModifier|false|false||unitnull|per milliliter|LabModifier|false|false||/mLnull|Solution Dosage Form|Drug|false|false||Solution
null|Solutions|Drug|false|false||Solution
null|Pharmaceutical Solutions|Drug|false|false||Solutionnull|Resolution|Finding|false|false||Solutionnull|Unit - NCI Thesaurus Property|LabModifier|false|false||units
null|Unit of Measure|LabModifier|false|false||units
null|Unit|LabModifier|false|false||unitsnull|Subcutaneous Route of Administration|Finding|false|false||Subcutaneousnull|subcutaneous|Modifier|false|false||Subcutaneousnull|Once a day, at bedtime|Time|false|false||at bedtimenull|Once a day, at bedtime|Time|false|false||bedtime
null|Bedtime (qualifier value)|Time|false|false||bedtimenull|insulin lispro|Drug|false|false||insulin lispro
null|insulin lispro|Drug|false|false||insulin lispro
null|insulin lispro|Drug|false|false||insulin lispronull|insulin, regular, human|Drug|false|false||insulin
null|Insulin [EPC]|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulinnull|INS gene|Finding|false|false||insulinnull|Insulin measurement|Procedure|false|false||insulinnull|insulin lispro|Drug|false|false||lispro
null|insulin lispro|Drug|false|false||lispro
null|insulin lispro|Drug|false|false||lispronull|Unit per Milliliter|LabModifier|false|false||unit/mLnull|Storage Unit|Device|false|false||unit
null|Unit device|Device|false|false||unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||unit
null|Unit of Measure|LabModifier|false|false||unit
null|Unit|LabModifier|false|false||unit
null|Enzyme Unit|LabModifier|false|false||unitnull|per milliliter|LabModifier|false|false||/mLnull|Solution Dosage Form|Drug|false|false||Solution
null|Solutions|Drug|false|false||Solution
null|Pharmaceutical Solutions|Drug|false|false||Solutionnull|Resolution|Finding|false|false||Solutionnull|sliding scale|Procedure|false|false||Sliding scalenull|Sliding|Finding|false|false||Slidingnull|Scale, LOINC Axis 5|Finding|false|false||scale
null|Base Number|Finding|false|false||scale
null|Scale - rank|Finding|false|false||scalenull|Integumentary scale|Anatomy|false|false||scalenull|Weight measurement scales|Device|false|false||scalenull|Scaling|Event|false|false||scalenull|Unit - NCI Thesaurus Property|LabModifier|false|false||units
null|Unit of Measure|LabModifier|false|false||units
null|Unit|LabModifier|false|false||unitsnull|insulin, regular, human|Drug|false|false||insulin
null|Insulin [EPC]|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulinnull|INS gene|Finding|false|false||insulinnull|Insulin measurement|Procedure|false|false||insulinnull|Subcutaneous Route of Administration|Finding|false|false||Subcutaneousnull|subcutaneous|Modifier|false|false||Subcutaneousnull|Three times daily|Time|false|false||three times a daynull|Thrice|LabModifier|false|false||three timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Transaction counts and value totals - provider|Finding|false|false||provider
null|Provider|Finding|false|false||providernull|albuterol sulfate|Drug|false|false||albuterol sulfate
null|albuterol sulfate|Drug|false|false||albuterol sulfatenull|albuterol|Drug|false|false||albuterol
null|albuterol|Drug|false|false||albuterolnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfate
null|Sulfates, Inorganic|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfatenull|mcg/actuation|LabModifier|false|false||mcg/actuationnull|microgram|LabModifier|false|false||mcgnull|Actuation (unit of presentation)|LabModifier|false|false||actuationnull|Facial Hemiatrophy|Disorder|false|false||HFAnull|High frequency audiometry|Procedure|false|false||HFAnull|Inhalers, Aerosol|Device|false|false||Aerosol Inhalernull|Aerosol Dose Form|Drug|false|false||Aerosolnull|Aerosols|Device|false|false||Aerosolnull|Inhaler (unit of presentation)|Finding|false|false||Inhalernull|Inhaler|Device|false|false||Inhalernull|Inhaler Dosing Unit|LabModifier|false|false||Inhalernull|Puff Dosing Unit|LabModifier|false|false||Puff
null|Picofarad|LabModifier|false|false||Puffnull|Inhalation Route of Administration|Finding|false|false||Inhalation
null|Inspiration (function)|Finding|false|false||Inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||Inhalationnull|Hour|Time|false|false||hoursnull|Dyspnea|Finding|false|false||SOBnull|Wheezing|Finding|false|false||wheezingnull|fluticasone|Drug|false|false||fluticasone
null|fluticasone|Drug|false|false||fluticasonenull|mcg/actuation|LabModifier|false|false||mcg/actuationnull|microgram|LabModifier|false|false||mcgnull|Actuation (unit of presentation)|LabModifier|false|false||actuationnull|Aerosol Dose Form|Drug|false|false||Aerosolnull|Aerosols|Device|false|false||Aerosolnull|Puff Dosing Unit|LabModifier|false|false||Puff
null|Picofarad|LabModifier|false|false||Puffnull|Inhalation Route of Administration|Finding|false|false||Inhalation
null|Inspiration (function)|Finding|false|false||Inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||Inhalationnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|2 times|Finding|false|false||2 timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|pantoprazole|Drug|false|false||pantoprazole
null|pantoprazole|Drug|false|false||pantoprazolenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Delayed Release Dosage Form|Drug|false|false||Delayed Releasenull|Views delayed|Attribute|false|false||Delayednull|Deferred|Time|false|false||Delayednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Delayed Release Dosage Form|Drug|false|false||Delayed Releasenull|Views delayed|Attribute|false|false||Delayednull|Deferred|Time|false|false||Delayednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Every twelve hours|Time|false|false||Q12Hnull|12 hours (qualifier value)|Time|false|false||12 hoursnull|Hour|Time|false|false||hoursnull|acetaminophen / oxycodone|Drug|false|false||oxycodone-acetaminophennull|oxycodone|Drug|false|false||oxycodone
null|oxycodone|Drug|false|false||oxycodonenull|Oxycodone measurement|Procedure|false|false||oxycodonenull|Acetaminophen [EPC]|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophennull|Acetaminophen measurement|Procedure|false|false||acetaminophennull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Every eight hours|Time|false|false||Q8Hnull|8 Hours|Time|false|false||8 hoursnull|Hour|Time|false|false||hoursnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|cholecalciferol|Drug|false|false||cholecalciferol (vitamin D3)
null|cholecalciferol|Drug|false|false||cholecalciferol (vitamin D3)
null|cholecalciferol|Drug|false|false||cholecalciferol (vitamin D3)null|cholecalciferol|Drug|false|false||cholecalciferol
null|cholecalciferol|Drug|false|false||cholecalciferol
null|cholecalciferol|Drug|false|false||cholecalciferolnull|vitamin D3|Drug|false|false||vitamin D3
null|vitamin D3|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitaminnull|Storage Unit|Device|false|false||unit
null|Unit device|Device|false|false||unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||unit
null|Unit of Measure|LabModifier|false|false||unit
null|Unit|LabModifier|false|false||unit
null|Enzyme Unit|LabModifier|false|false||unitnull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|metronidazole|Drug|false|false||metronidazole
null|metronidazole|Drug|false|false||metronidazolenull|Lotion|Drug|false|false||Lotionnull|HL7 Version 2.5 - Application|Finding|false|false||application
null|Application Document|Finding|false|false||application
null|Computer Application|Finding|false|false||application
null|Regulatory Application|Finding|false|false||application
null|Apply|Finding|false|false||applicationnull|Application procedure|Procedure|false|false||applicationnull|Application - unit of product usage|LabModifier|false|false||applicationnull|Topical Dosage Form|Drug|false|false||Topicalnull|Topical Route of Administration|Finding|false|false||Topicalnull|Topical surface|Modifier|false|false||Topicalnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|null|Attribute|false|false||Primary diagnosisnull|Principal diagnosis|Modifier|false|false||Primary diagnosisnull|True primary (qualifier value)|Time|false|false||Primarynull|Primary|Modifier|false|false||Primarynull|Diagnosis Classification - Diagnosis|Finding|false|false||diagnosis
null|diagnosis aspects|Finding|false|false||diagnosisnull|Diagnosis|Procedure|false|false||diagnosisnull|null|Attribute|false|false||diagnosisnull|Atypical chest pain|Finding|false|false||Atypical chest painnull|atypia morphology|Finding|false|false||Atypicalnull|Atypical|Modifier|false|false||Atypicalnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Secondary diagnosis|Finding|false|false||Secondary diagnosisnull|null|Attribute|false|false||Secondary diagnosisnull|Neoplasm Metastasis|Disorder|false|false||Secondarynull|metastatic qualifier|Finding|false|false||Secondarynull|Secondary to|Modifier|false|false||Secondarynull|second (number)|LabModifier|false|false||Secondarynull|Diagnosis Classification - Diagnosis|Finding|false|false||diagnosis
null|diagnosis aspects|Finding|false|false||diagnosisnull|Diagnosis|Procedure|false|false||diagnosisnull|null|Attribute|false|false||diagnosisnull|Coronary Artery Disease|Disorder|false|false||Coronary artery disease
null|Coronary Arteriosclerosis|Disorder|false|false||Coronary artery diseasenull|Coronary artery|Anatomy|false|false||Coronary arterynull|Heart|Anatomy|false|false||Coronarynull|Coronary|Modifier|false|false||Coronarynull|Arteriopathic disease|Disorder|false|false||artery diseasenull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Disease|Disorder|false|false||diseasenull|Hypertensive disease|Disorder|false|false||Hypertensionnull|Hyperlipidemia|Disorder|false|false||Hyperlipidemia
null|Hyperlipoproteinemias|Disorder|false|false||Hyperlipidemianull|Serum lipids high (finding)|Finding|false|false||Hyperlipidemianull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Type 2 Diabetes Mellitusnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Type 2 Diabetesnull|Type 2|Finding|false|false||Type 2null|Type - ParameterizedDataType|Finding|false|false||Type
null|SGCG gene|Finding|false|false||Typenull|null|Modifier|false|false||Typenull|Diabetes Mellitus|Disorder|false|false||Diabetes Mellitusnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Diabetes
null|Diabetes|Disorder|false|false||Diabetes
null|Diabetes Mellitus|Disorder|false|false||Diabetesnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Disease|Disorder|false|false||Conditionnull|Logical Condition|Finding|false|false||Conditionnull|null|Attribute|false|false||Conditionnull|Condition|Modifier|false|false||Conditionnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|Discharge instructions|Finding|false|false||Discharge Instructionsnull|hospital discharge instructions (treatment)|Procedure|false|false||Discharge Instructionsnull|null|Attribute|false|false||Discharge Instructionsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|Production Class Code - Pleasure|Finding|false|false||pleasure
null|pleasurable emotion|Finding|false|false||pleasurenull|Pleasure - Animals raised for recreation|Entity|false|false||pleasurenull|care of - AddressPartType|Finding|false|false||care ofnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Hospitalization|Procedure|false|false||hospitalizationnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Nuclear (incident type)|Modifier|false|false||nuclear
null|Nuclear (nucleus)|Modifier|false|false||nuclearnull|Stress bismuth subsalicylate|Drug|false|false||stress
null|Stress bismuth subsalicylate|Drug|false|false||stressnull|Stress|Finding|false|false||stressnull|W stress|Attribute|false|false||stressnull|Tests (qualifier value)|Finding|false|false||test
null|Testing|Finding|false|false||testnull|Laboratory Procedures|Procedure|false|false||testnull|Test - temporal region|Anatomy|false|false||testnull|Test Result|Lab|false|false||testnull|Test Dosing Unit|LabModifier|false|false||testnull|Observation Interpretation - Abnormal|Finding|false|false||abnormal
null|Abnormal|Finding|false|false||abnormalnull|Cardiac attachment|Finding|false|false||cardiacnull|Heart|Anatomy|false|false||cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||cardiacnull|Catheterization|Procedure|false|false||catheterizationnull|Partial Blockage within Medical Device|Finding|false|false||blockage
null|Blockage (obstruction - finding)|Finding|false|false||blockage
null|null|Finding|false|false||blockagenull|Structure of circumflex branch of left coronary artery|Anatomy|false|false||left circumflex coronary arterynull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Structure of circumflex branch of left coronary artery|Anatomy|false|false||circumflex coronary arterynull|Circumflex|Modifier|false|false||circumflexnull|Coronary artery|Anatomy|false|false||coronary arterynull|Heart|Anatomy|false|false||coronarynull|Coronary|Modifier|false|false||coronarynull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Malignant neoplasm of heart|Disorder|false|false||heart
null|benign neoplasm of heart|Disorder|false|false||heartnull|HEART PROBLEM|Finding|false|false||heartnull|Chest>Heart|Anatomy|false|false||heart
null|Heart|Anatomy|false|false||heartnull|Blood Vessel|Anatomy|false|false||vesselsnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Following|Time|false|false||following
null|Status post|Time|false|false||followingnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Potassium supplement|Drug|false|false||potassium supplement
null|Potassium supplement|Drug|false|false||potassium supplementnull|Potassium supplement|Drug|false|false||potassium
null|Dietary Potassium|Drug|false|false||potassium
null|potassium|Drug|false|false||potassium
null|potassium|Drug|false|false||potassium
null|potassium|Drug|false|false||potassium
null|Potassium Drug Class|Drug|false|false||potassium
null|Potassium supplement|Drug|false|false||potassiumnull|Potassium metabolic function|Finding|false|false||potassiumnull|Potassium measurement|Procedure|false|false||potassiumnull|Dietary Supplements|Drug|false|false||supplementnull|Supplement - Diet Code Specification Type|Finding|false|false||supplement
null|Supplement|Finding|false|false||supplement
null|Supplement (document)|Finding|false|false||supplementnull|Potassium Drug Class|Drug|false|false||potassium
null|Dietary Potassium|Drug|false|false||potassium
null|potassium|Drug|false|false||potassium
null|potassium|Drug|false|false||potassium
null|potassium|Drug|false|false||potassium
null|Potassium supplement|Drug|false|false||potassium
null|Potassium supplement|Drug|false|false||potassiumnull|Potassium metabolic function|Finding|false|false||potassiumnull|Potassium measurement|Procedure|false|false||potassiumnull|Levels (qualifier value)|Modifier|false|false||levelsnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|atorvastatin|Drug|false|false||atorvastatin
null|atorvastatin|Drug|false|false||atorvastatinnull|Lipitor|Drug|false|false||lipitor
null|Lipitor|Drug|false|false||lipitornull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Daily|Time|false|false||dailynull|lisinopril|Drug|false|false||lisinopril
null|lisinopril|Drug|false|false||lisinoprilnull|Lasix|Drug|false|false||lasix
null|Lasix|Drug|false|false||lasixnull|furosemide|Drug|false|false||furosemide
null|furosemide|Drug|false|false||furosemidenull|Primary Care Physicians|Subject|false|false||primary care physician
null|Primary care provider|Subject|false|false||primary care physiciannull|Location Service Code - Primary Care|Finding|false|false||primary carenull|Primary Health Care|Procedure|false|false||primary carenull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|null|Attribute|false|false||physiciannull|Physicians|Subject|false|false||physiciannull|Repeat Object|Finding|false|false||repeat
null|Repeat|Finding|false|false||repeatnull|Repeat Pattern|Time|false|false||repeatnull|Primary Care Physicians|Subject|false|false||primary care physician
null|Primary care provider|Subject|false|false||primary care physiciannull|Location Service Code - Primary Care|Finding|false|false||primary carenull|Primary Health Care|Procedure|false|false||primary carenull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|null|Attribute|false|false||physiciannull|Physicians|Subject|false|false||physiciannull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Appointments|Event|false|false||appointmentsnull|Appointments|Event|false|false||appointmentsnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions