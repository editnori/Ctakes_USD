 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|48,57|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|48,57|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|48,62|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|82,91|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|82,91|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|82,91|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|82,91|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|82,91|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|82,96|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|114,119|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|114,119|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|114,119|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|138,141|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|138,141|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|138,141|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|138,141|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|138,141|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|149,156|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|149,156|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|Allergies|185,190|false|false|false|C0749139|sulfa|Sulfa
Event|Event|Allergies|185,190|false|false|false|||Sulfa
Drug|Antibiotic|Allergies|192,203|false|false|false|C0038760;C0599503;C3536763|Sulfonamide Anti-Infective Agents;Sulfonamide [EPC];Sulfonamides|Sulfonamide
Drug|Organic Chemical|Allergies|192,203|false|false|false|C0038760;C0599503;C3536763|Sulfonamide Anti-Infective Agents;Sulfonamide [EPC];Sulfonamides|Sulfonamide
Drug|Pharmacologic Substance|Allergies|192,203|false|false|false|C0038760;C0599503;C3536763|Sulfonamide Anti-Infective Agents;Sulfonamide [EPC];Sulfonamides|Sulfonamide
Drug|Antibiotic|Allergies|204,215|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|Antibiotics
Event|Event|Allergies|204,215|false|false|false|||Antibiotics
Disorder|Injury or Poisoning|Allergies|219,230|false|false|false|C0161486;C2876539|Poisoning by penicillin;Poisoning by, adverse effect of and underdosing of penicillins|Penicillins
Drug|Antibiotic|Allergies|219,230|false|false|false|C0030842|penicillins|Penicillins
Drug|Organic Chemical|Allergies|219,230|false|false|false|C0030842|penicillins|Penicillins
Event|Event|Allergies|219,230|false|false|false|||Penicillins
Finding|Pathologic Function|Allergies|219,230|false|false|false|C0413443|Adverse reaction to penicillins|Penicillins
Event|Event|Allergies|233,242|false|false|false|||Attending
Finding|Functional Concept|Allergies|233,242|false|false|false|C1999232|Attending (action)|Attending
Anatomy|Body Location or Region|Chief Complaint|268,272|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|Chief Complaint|268,272|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|Chief Complaint|268,272|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Finding|Sign or Symptom|Chief Complaint|268,277|false|false|false|C0007859|Neck Pain|neck pain
Attribute|Clinical Attribute|Chief Complaint|273,277|false|false|false|C2598155||pain
Event|Event|Chief Complaint|273,277|false|false|false|||pain
Finding|Functional Concept|Chief Complaint|273,277|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Chief Complaint|273,277|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Chief Complaint|282,286|false|false|false|C0085639|Falls|fall
Finding|Classification|Chief Complaint|289,294|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|295,303|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|295,303|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|307,325|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|316,325|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|316,325|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|316,325|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|316,325|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|316,325|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|Chief Complaint|340,349|true|false|false|||Admission
Procedure|Health Care Activity|Chief Complaint|340,349|true|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Finding|Finding|History of Present Illness|384,388|false|false|false|C1706180|Male Gender|male
Event|Event|History of Present Illness|389,400|false|false|false|||transferred
Finding|Idea or Concept|History of Present Illness|414,422|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|History of Present Illness|428,438|false|false|false|||evaluation
Finding|Idea or Concept|History of Present Illness|428,438|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|History of Present Illness|428,438|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Anatomy|Body Location or Region|History of Present Illness|442,450|false|false|false|C0027530|Neck|cervical
Disorder|Injury or Poisoning|History of Present Illness|455,463|false|false|false|C0016658|Fracture|fracture
Event|Event|History of Present Illness|455,463|false|false|false|||fracture
Finding|Body Substance|History of Present Illness|475,482|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|475,482|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|475,482|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|488,498|false|false|false|||attempting
Event|Event|History of Present Illness|502,505|false|false|false|||use
Event|Event|History of Present Illness|545,552|false|false|false|||hitting
Finding|Finding|History of Present Illness|545,552|false|false|false|C0596020|Does hit (finding)|hitting
Anatomy|Body Location or Region|History of Present Illness|570,574|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|570,574|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|History of Present Illness|570,574|false|false|false|C0362076|Problems with head|head
Event|Event|History of Present Illness|570,574|false|false|false|||head
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|570,574|false|false|false|C0876917|Procedure on head|head
Event|Event|History of Present Illness|589,593|true|false|false|||loss
Finding|Finding|History of Present Illness|589,593|true|false|false|C5890125|Loss (adaptation)|loss
Finding|Finding|History of Present Illness|589,610|true|false|false|C0041657|Unconscious State|loss of consciousness
Event|Event|History of Present Illness|597,610|true|false|false|||consciousness
Finding|Finding|History of Present Illness|597,610|true|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|consciousness
Finding|Mental Process|History of Present Illness|597,610|true|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|consciousness
Finding|Body Substance|History of Present Illness|617,624|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|617,624|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|617,624|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|625,634|false|false|false|||complains
Event|Event|History of Present Illness|638,646|false|false|false|||headache
Finding|Sign or Symptom|History of Present Illness|638,646|false|false|false|C0018681|Headache|headache
Anatomy|Body Location or Region|History of Present Illness|651,655|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|History of Present Illness|651,655|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|History of Present Illness|651,655|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Finding|Sign or Symptom|History of Present Illness|651,660|false|false|false|C0007859|Neck Pain|neck pain
Attribute|Clinical Attribute|History of Present Illness|656,660|false|false|false|C2598155||pain
Event|Event|History of Present Illness|656,660|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|656,660|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|656,660|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Idea or Concept|History of Present Illness|675,683|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Body Substance|History of Present Illness|688,695|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|688,695|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|688,695|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Anatomy|Body Location or Region|History of Present Illness|704,708|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|704,708|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|History of Present Illness|704,708|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|704,708|false|false|false|C0876917|Procedure on head|head
Disorder|Injury or Poisoning|History of Present Illness|704,719|false|false|false|C0856548|Laceration of head|head laceration
Disorder|Injury or Poisoning|History of Present Illness|709,719|false|false|false|C0043246|Laceration|laceration
Event|Event|History of Present Illness|709,719|false|false|false|||laceration
Event|Event|History of Present Illness|720,727|false|false|false|||stapled
Procedure|Diagnostic Procedure|History of Present Illness|731,738|false|false|false|C0040405|X-Ray Computed Tomography|CT scan
Event|Event|History of Present Illness|734,738|false|false|false|||scan
Procedure|Diagnostic Procedure|History of Present Illness|734,738|false|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Event|Event|History of Present Illness|744,755|false|false|false|||demonstrate
Disorder|Injury or Poisoning|History of Present Illness|760,768|false|false|false|C0016658|Fracture|fracture
Event|Event|History of Present Illness|760,768|false|false|false|||fracture
Finding|Body Substance|History of Present Illness|774,781|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|774,781|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|774,781|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|782,788|true|false|false|||denies
Event|Event|History of Present Illness|793,801|true|false|false|||numbness
Finding|Finding|History of Present Illness|793,801|true|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|History of Present Illness|793,801|true|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Disorder|Disease or Syndrome|History of Present Illness|804,812|true|false|false|C0030554|Paresthesia|tingling
Event|Event|History of Present Illness|804,812|true|false|false|||tingling
Finding|Sign or Symptom|History of Present Illness|804,812|true|false|false|C2242996|Has tingling sensation|tingling
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|820,824|true|false|false|C0446516|Upper arm|arms
Attribute|Clinical Attribute|History of Present Illness|820,824|true|false|false|C5782111||arms
Disorder|Neoplastic Process|History of Present Illness|820,824|true|false|false|C0206655|Alveolar rhabdomyosarcoma|arms
Finding|Gene or Genome|History of Present Illness|820,824|true|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Finding|Intellectual Product|History of Present Illness|820,824|true|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|828,832|false|false|false|C1140621|Leg|legs
Attribute|Clinical Attribute|History of Present Illness|828,832|false|false|false|C5781420||legs
Event|Event|History of Present Illness|837,845|true|false|false|||weakness
Finding|Sign or Symptom|History of Present Illness|837,845|true|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|853,857|true|false|false|C0446516|Upper arm|arms
Attribute|Clinical Attribute|History of Present Illness|853,857|true|false|false|C5782111||arms
Disorder|Neoplastic Process|History of Present Illness|853,857|true|false|false|C0206655|Alveolar rhabdomyosarcoma|arms
Finding|Gene or Genome|History of Present Illness|853,857|true|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Finding|Intellectual Product|History of Present Illness|853,857|true|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|861,865|true|false|false|C1140621|Leg|legs
Attribute|Clinical Attribute|History of Present Illness|861,865|true|false|false|C5781420||legs
Event|Event|History of Present Illness|868,874|true|false|false|||Denies
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|879,884|true|false|false|C0021853|Intestines|bowel
Disorder|Disease or Syndrome|History of Present Illness|879,897|true|false|false|C0015732|Fecal Incontinence|bowel incontinence
Disorder|Disease or Syndrome|History of Present Illness|885,897|true|false|false|C0021167|Incontinence|incontinence
Event|Event|History of Present Illness|885,897|true|false|false|||incontinence
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|901,908|true|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|History of Present Illness|901,908|true|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|901,908|true|false|false|C0872388|Procedures on bladder|bladder
Finding|Functional Concept|History of Present Illness|901,918|true|false|false|C0080274|Urinary Retention|bladder retention
Attribute|Clinical Attribute|History of Present Illness|909,918|true|false|false|C1318143|Retention - dental|retention
Event|Event|History of Present Illness|909,918|true|false|false|||retention
Finding|Cell Function|History of Present Illness|909,918|true|false|false|C0035280;C0080274;C0333117;C1753315|Retention (Psychology);Retention of content;Urinary Retention;cellular entity retention|retention
Finding|Functional Concept|History of Present Illness|909,918|true|false|false|C0035280;C0080274;C0333117;C1753315|Retention (Psychology);Retention of content;Urinary Retention;cellular entity retention|retention
Finding|Mental Process|History of Present Illness|909,918|true|false|false|C0035280;C0080274;C0333117;C1753315|Retention (Psychology);Retention of content;Urinary Retention;cellular entity retention|retention
Attribute|Clinical Attribute|History of Present Illness|931,941|true|false|false|C2926599||anesthesia
Drug|Pharmacologic Substance|History of Present Illness|931,941|true|false|false|C4049933|Anesthesia substance|anesthesia
Event|Event|History of Present Illness|931,941|true|false|false|||anesthesia
Finding|Finding|History of Present Illness|931,941|true|false|false|C0278134;C2219802|Absence of sensation|anesthesia
Finding|Sign or Symptom|History of Present Illness|931,941|true|false|false|C0278134;C2219802|Absence of sensation|anesthesia
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|931,941|true|false|false|C0002903;C0002912|Anesthesia procedures;Dental anesthesia|anesthesia
Event|Event|History of Present Illness|943,949|true|false|false|||Denies
Anatomy|Body Location or Region|History of Present Illness|954,959|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|954,959|true|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|954,964|true|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|954,964|true|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|960,964|true|false|false|C2598155||pain
Event|Event|History of Present Illness|960,964|true|false|false|||pain
Finding|Functional Concept|History of Present Illness|960,964|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|960,964|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|966,975|true|false|false|||shortness
Attribute|Clinical Attribute|History of Present Illness|966,985|true|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|History of Present Illness|966,985|true|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|History of Present Illness|979,985|true|false|false|C0225386|Breath|breath
Anatomy|Body Location or Region|History of Present Illness|990,999|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|History of Present Illness|990,1004|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|History of Present Illness|1000,1004|false|false|false|C2598155||pain
Event|Event|History of Present Illness|1000,1004|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|1000,1004|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1000,1004|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Past Medical History|1034,1037|false|false|false|||PMH
Finding|Finding|Past Medical History|1034,1037|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|PMH
Event|Event|Past Medical History|1042,1045|false|false|false|||fib
Finding|Gene or Genome|Past Medical History|1042,1045|false|false|false|C1414538|FBL gene|fib
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1047,1052|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|Past Medical History|1047,1052|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|Past Medical History|1047,1052|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Finding|Finding|Past Medical History|1047,1052|false|false|false|C0750873|COLON PROBLEM|colon
Disorder|Neoplastic Process|Past Medical History|1047,1055|false|true|false|C0007102|Malignant tumor of colon|colon ca
Event|Event|Past Medical History|1053,1055|false|false|false|||ca
Disorder|Disease or Syndrome|Past Medical History|1057,1060|false|false|false|C0020538|Hypertensive disease|htn
Event|Event|Past Medical History|1057,1060|false|false|false|||htn
Disorder|Disease or Syndrome|Past Medical History|1062,1066|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|copd
Drug|Pharmacologic Substance|Past Medical History|1062,1066|false|false|false|C1647218|COPD pharmacologic substance|copd
Event|Event|Past Medical History|1062,1066|false|false|false|||copd
Finding|Gene or Genome|Past Medical History|1062,1066|false|false|false|C1412502|ARCN1 gene|copd
Disorder|Congenital Abnormality|Past Medical History|1070,1073|false|false|false|C0026760|Multiple Epiphyseal Dysplasia|MED
Event|Event|Past Medical History|1070,1073|false|false|false|||MED
Finding|Gene or Genome|Past Medical History|1070,1073|false|false|false|C1413596;C1413597;C1419866;C1456376;C1549978;C4321267;C5781216|COL9A2 gene;COL9A3 gene;COMP gene;COMP wt Allele;Master of Education;SCN8A gene;SCN8A wt Allele|MED
Finding|Intellectual Product|Past Medical History|1070,1073|false|false|false|C1413596;C1413597;C1419866;C1456376;C1549978;C4321267;C5781216|COL9A2 gene;COL9A3 gene;COMP gene;COMP wt Allele;Master of Education;SCN8A gene;SCN8A wt Allele|MED
Drug|Hazardous or Poisonous Substance|Past Medical History|1075,1083|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|Past Medical History|1075,1083|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|Past Medical History|1075,1083|false|false|false|C0043031|warfarin|warfarin
Event|Event|Past Medical History|1075,1083|false|false|false|||warfarin
Drug|Organic Chemical|Past Medical History|1085,1096|false|false|false|C0002144|allopurinol|allopurinol
Drug|Pharmacologic Substance|Past Medical History|1085,1096|false|false|false|C0002144|allopurinol|allopurinol
Event|Event|Past Medical History|1085,1096|false|false|false|||allopurinol
Drug|Amino Acid, Peptide, or Protein|Past Medical History|1098,1104|false|false|false|C0678172|Asacol|asacol
Drug|Pharmacologic Substance|Past Medical History|1098,1104|false|false|false|C0678172|Asacol|asacol
Event|Event|Past Medical History|1098,1104|false|false|false|||asacol
Event|Event|Past Medical History|1108,1111|false|false|false|||ALL
Drug|Organic Chemical|Past Medical History|1113,1116|false|false|false|C0033017|Pregnenolone Carbonitrile|pcn
Drug|Pharmacologic Substance|Past Medical History|1113,1116|false|false|false|C0033017|Pregnenolone Carbonitrile|pcn
Event|Event|Past Medical History|1113,1116|false|false|false|||pcn
Finding|Gene or Genome|Past Medical History|1113,1116|false|false|false|C1418643;C1826553;C4050150|PCNT gene;PLEC gene;PLEC wt Allele|pcn
Drug|Pharmacologic Substance|Past Medical History|1118,1123|false|false|false|C0749139|sulfa|sulfa
Event|Event|Past Medical History|1118,1123|false|false|false|||sulfa
Event|Event|General Exam|1185,1191|false|false|false|||collar
Event|Activity|General Exam|1195,1200|false|false|false|C1882509|put - instruction imperative|place
Event|Event|General Exam|1195,1200|false|false|false|||place
Finding|Functional Concept|General Exam|1195,1200|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|General Exam|1195,1200|false|false|false|C1533810||place
Drug|Amino Acid, Peptide, or Protein|General Exam|1216,1219|false|false|false|C1366678;C1433371;C4049852|L-Type Amino Acid Transporter;LAT protein, human;ORC3 protein, human|lat
Drug|Biologically Active Substance|General Exam|1216,1219|false|false|false|C1366678;C1433371;C4049852|L-Type Amino Acid Transporter;LAT protein, human;ORC3 protein, human|lat
Drug|Immunologic Factor|General Exam|1216,1219|false|false|false|C1366678;C1433371;C4049852|L-Type Amino Acid Transporter;LAT protein, human;ORC3 protein, human|lat
Finding|Gene or Genome|General Exam|1216,1219|false|false|false|C1335085;C1425844;C1705279;C2240043|LAT gene;ORC3 gene;ORC3 wt Allele;SPNS1 gene|lat
Anatomy|Body Part, Organ, or Organ Component|General Exam|1220,1223|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|General Exam|1220,1223|false|false|false|C3495676|Anorectal Malformations|arm
Event|Event|General Exam|1220,1223|false|false|false|||arm
Finding|Gene or Genome|General Exam|1220,1223|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|General Exam|1220,1223|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|General Exam|1220,1223|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|General Exam|1220,1223|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Anatomy|Body Part, Organ, or Organ Component|General Exam|1227,1232|false|false|false|C0040067|Thumb structure|thumb
Anatomy|Body Part, Organ, or Organ Component|General Exam|1249,1255|false|false|false|C0016129;C0851278;C4299059|Fingers;Fingers not including thumb;Upper extremity>Finger|finger
Disorder|Congenital Abnormality|General Exam|1258,1261|false|false|false|C0026760|Multiple Epiphyseal Dysplasia|med
Finding|Gene or Genome|General Exam|1258,1261|false|false|false|C1413596;C1413597;C1419866;C1456376;C1549978;C4321267;C5781216|COL9A2 gene;COL9A3 gene;COMP gene;COMP wt Allele;Master of Education;SCN8A gene;SCN8A wt Allele|med
Finding|Intellectual Product|General Exam|1258,1261|false|false|false|C1413596;C1413597;C1419866;C1456376;C1549978;C4321267;C5781216|COL9A2 gene;COL9A3 gene;COMP gene;COMP wt Allele;Master of Education;SCN8A gene;SCN8A wt Allele|med
Anatomy|Body Part, Organ, or Organ Component|General Exam|1262,1265|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|General Exam|1262,1265|false|false|false|C3495676|Anorectal Malformations|arm
Event|Event|General Exam|1262,1265|false|false|false|||arm
Finding|Gene or Genome|General Exam|1262,1265|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|General Exam|1262,1265|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|General Exam|1262,1265|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|General Exam|1262,1265|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Finding|Finding|General Exam|1280,1286|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Finding|General Exam|1294,1300|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Finding|General Exam|1308,1314|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|General Exam|1322,1328|false|false|false|||intact
Finding|Finding|General Exam|1322,1328|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Finding|General Exam|1342,1348|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Finding|General Exam|1356,1362|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Finding|General Exam|1370,1376|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|General Exam|1384,1390|false|false|false|||intact
Finding|Finding|General Exam|1384,1390|false|false|false|C1554187|Gender Status - Intact|intact
Anatomy|Body Location or Region|General Exam|1399,1404|false|false|false|C0225442;C0460005;C1523842|Trunk of elephant;Trunk structure;dendritic shaft|Trunk
Anatomy|Body Part, Organ, or Organ Component|General Exam|1399,1404|false|false|false|C0225442;C0460005;C1523842|Trunk of elephant;Trunk structure;dendritic shaft|Trunk
Anatomy|Cell Component|General Exam|1399,1404|false|false|false|C0225442;C0460005;C1523842|Trunk of elephant;Trunk structure;dendritic shaft|Trunk
Event|Event|General Exam|1406,1412|false|false|false|||intact
Finding|Finding|General Exam|1406,1412|false|false|false|C1554187|Gender Status - Intact|intact
Anatomy|Body Location or Region|General Exam|1449,1454|false|false|false|C0018246;C0816951;C4266533|Inguinal part of abdomen;Inguinal region;Pelvis>Groin|Groin
Anatomy|Body Location or Region|General Exam|1456,1460|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|Knee
Anatomy|Body Part, Organ, or Organ Component|General Exam|1456,1460|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|Knee
Anatomy|Body Space or Junction|General Exam|1456,1460|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|Knee
Procedure|Diagnostic Procedure|General Exam|1456,1460|false|false|false|C0562271|Examination of knee joint|Knee
Disorder|Congenital Abnormality|General Exam|1466,1469|false|false|false|C0026760|Multiple Epiphyseal Dysplasia|Med
Finding|Gene or Genome|General Exam|1466,1469|false|false|false|C1413596;C1413597;C1419866;C1456376;C1549978;C4321267;C5781216|COL9A2 gene;COL9A3 gene;COMP gene;COMP wt Allele;Master of Education;SCN8A gene;SCN8A wt Allele|Med
Finding|Intellectual Product|General Exam|1466,1469|false|false|false|C1413596;C1413597;C1419866;C1456376;C1549978;C4321267;C5781216|COL9A2 gene;COL9A3 gene;COMP gene;COMP wt Allele;Master of Education;SCN8A gene;SCN8A wt Allele|Med
Anatomy|Body Location or Region|General Exam|1470,1474|false|false|false|C0230445;C1305418|Structure of calf of leg|Calf
Anatomy|Body Part, Organ, or Organ Component|General Exam|1470,1474|false|false|false|C0230445;C1305418|Structure of calf of leg|Calf
Anatomy|Body Part, Organ, or Organ Component|General Exam|1477,1480|false|false|false|C0228547|Clava structure (body structure)|Grt
Anatomy|Body Part, Organ, or Organ Component|General Exam|1481,1484|false|false|false|C0040357;C4299090|Lower extremity>Toes;Toes|Toe
Anatomy|Body Part, Organ, or Organ Component|General Exam|1490,1493|false|false|false|C0040357;C4299090|Lower extremity>Toes;Toes|Toe
Anatomy|Body Location or Region|General Exam|1501,1506|false|false|false|C0039866;C4299091|Lower extremity>Thigh;Thigh structure|Thigh
Event|Event|General Exam|1599,1604|false|false|false|||Motor
Finding|Functional Concept|General Exam|1599,1604|false|false|false|C1513492|motor movement|Motor
Anatomy|Body Part, Organ, or Organ Component|General Exam|1615,1618|false|false|false|C0175372;C3495985|Structure of inferior brachium of corpora quadrigemina;nucleus of the brachium of the inferior colliculus|Bic
Drug|Organic Chemical|General Exam|1615,1618|false|false|false|C0063382|imidazole mustard|Bic
Drug|Pharmacologic Substance|General Exam|1615,1618|false|false|false|C0063382|imidazole mustard|Bic
Finding|Gene or Genome|General Exam|1615,1618|false|false|false|C1537811;C2681931|MIR155 gene;MIR155HG gene|Bic
Procedure|Therapeutic or Preventive Procedure|General Exam|1615,1618|false|false|false|C5202575|BIC Regimen|Bic
Finding|Gene or Genome|General Exam|1628,1631|false|false|false|C0814229;C3891460|TRI-AAT9-1 gene;Temptation and Restraint Inventory|Tri
Finding|Intellectual Product|General Exam|1628,1631|false|false|false|C0814229;C3891460|TRI-AAT9-1 gene;Temptation and Restraint Inventory|Tri
Finding|Finding|General Exam|1840,1848|false|false|false|C0034935|Babinski Reflex|Babinski
Event|Event|General Exam|1851,1859|false|false|false|||negative
Finding|Classification|General Exam|1851,1859|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|General Exam|1851,1859|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|General Exam|1851,1859|false|false|false|C5237010|Expression Negative|negative
Event|Event|General Exam|1861,1867|false|false|false|||Clonus
Finding|Sign or Symptom|General Exam|1861,1867|false|false|false|C0009024|Clonus|Clonus
Event|Event|General Exam|1873,1880|true|false|false|||present
Finding|Finding|General Exam|1873,1880|true|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|General Exam|1873,1880|true|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Body Substance|Hospital Course|1910,1917|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|1910,1917|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|1910,1917|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|1922,1930|false|false|false|||admitted
Finding|Finding|Hospital Course|1946,1953|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Finding|Functional Concept|Hospital Course|1946,1953|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Finding|Idea or Concept|Hospital Course|1946,1953|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Procedure|Therapeutic or Preventive Procedure|Hospital Course|1946,1953|false|false|false|C0543467|Operative Surgical Procedures|Surgery
Event|Occupational Activity|Hospital Course|1954,1961|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|Hospital Course|1954,1961|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|Hospital Course|1967,1978|false|false|false|||observation
Finding|Finding|Hospital Course|1967,1978|false|false|false|C0478530;C1548358;C1554188;C5890437|Examination and observation for unspecified reason;Observation (finding)|observation
Finding|Idea or Concept|Hospital Course|1967,1978|false|false|false|C0478530;C1548358;C1554188;C5890437|Examination and observation for unspecified reason;Observation (finding)|observation
Procedure|Diagnostic Procedure|Hospital Course|1967,1978|false|false|false|C0302523;C0700325;C1964257|Observation - diagnostic procedure;Observation in research;Patient observation|observation
Procedure|Health Care Activity|Hospital Course|1967,1978|false|false|false|C0302523;C0700325;C1964257|Observation - diagnostic procedure;Observation in research;Patient observation|observation
Procedure|Research Activity|Hospital Course|1967,1978|false|false|false|C0302523;C0700325;C1964257|Observation - diagnostic procedure;Observation in research;Patient observation|observation
Disorder|Injury or Poisoning|Hospital Course|1990,1998|false|false|false|C0016658|Fracture|fracture
Event|Event|Hospital Course|1990,1998|false|false|false|||fracture
Event|Event|Hospital Course|2001,2005|false|false|false|||TEDs
Event|Event|Hospital Course|2022,2026|false|false|false|||used
Disorder|Disease or Syndrome|Hospital Course|2032,2049|false|false|false|C0589110|Postoperative deep vein thrombosis|postoperative DVT
Anatomy|Body Location or Region|Hospital Course|2046,2049|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Hospital Course|2046,2049|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Hospital Course|2046,2049|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|Hospital Course|2046,2049|false|false|false|||DVT
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2046,2061|false|false|false|C0853245|DVT prophylaxis|DVT prophylaxis
Event|Event|Hospital Course|2050,2061|false|false|false|||prophylaxis
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2050,2061|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Drug|Food|Hospital Course|2064,2068|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|Diet
Event|Event|Hospital Course|2064,2068|false|false|false|||Diet
Finding|Functional Concept|Hospital Course|2064,2068|false|false|false|C1549512|diet - supply|Diet
Procedure|Health Care Activity|Hospital Course|2064,2068|false|false|false|C0012159|Diet therapy|Diet
Event|Event|Hospital Course|2073,2081|false|false|false|||advanced
Event|Event|Hospital Course|2085,2094|false|false|false|||tolerated
Finding|Body Substance|Hospital Course|2102,2109|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|2102,2109|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|2102,2109|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|2114,2123|false|false|false|||tolerated
Anatomy|Body Space or Junction|Hospital Course|2124,2128|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|2124,2128|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|2124,2128|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|2124,2128|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Sign or Symptom|Hospital Course|2124,2133|false|false|false|C0221776|Oral pain|oral pain
Attribute|Clinical Attribute|Hospital Course|2129,2133|false|false|false|C2598155||pain
Event|Event|Hospital Course|2129,2133|false|false|false|||pain
Finding|Functional Concept|Hospital Course|2129,2133|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|2129,2133|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Pharmacologic Substance|Hospital Course|2134,2144|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Hospital Course|2134,2144|false|false|false|||medication
Finding|Intellectual Product|Hospital Course|2134,2144|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Finding|Finding|Hospital Course|2146,2154|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|Hospital Course|2146,2154|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|Hospital Course|2146,2154|false|false|false|C0031809|Physical Examination|Physical
Finding|Intellectual Product|Hospital Course|2146,2162|false|false|false|C1547999|Diagnostic Service Section ID - Physical Therapy|Physical therapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2146,2162|false|false|false|C0949766|Physical therapy|Physical therapy
Event|Event|Hospital Course|2155,2162|false|false|false|||therapy
Finding|Finding|Hospital Course|2155,2162|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|Hospital Course|2155,2162|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2155,2162|false|false|false|C0087111|Therapeutic procedure|therapy
Event|Event|Hospital Course|2168,2177|false|false|false|||consulted
Event|Event|Hospital Course|2182,2194|false|false|false|||mobilization
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2182,2194|false|false|false|C0185112;C2080791|Mobilization (procedure);physical therapy mobilization (treatment)|mobilization
Event|Event|Hospital Course|2195,2198|false|false|false|||OOB
Event|Event|Hospital Course|2202,2210|false|false|false|||ambulate
Finding|Finding|Hospital Course|2202,2210|false|false|false|C4036205|Ambulate|ambulate
Event|Event|Hospital Course|2216,2224|false|false|false|||remained
Event|Event|Hospital Course|2226,2238|false|false|false|||hypertensive
Finding|Finding|Hospital Course|2226,2238|false|false|false|C0857121|Hypertensive (finding)|hypertensive
Drug|Pharmacologic Substance|Hospital Course|2257,2265|false|false|false|C0013227|Pharmaceutical Preparations|Medicine
Procedure|Health Care Activity|Hospital Course|2257,2273|false|false|false|C0746478|MEDICINE CONSULT|Medicine consult
Event|Event|Hospital Course|2266,2273|false|false|false|||consult
Procedure|Health Care Activity|Hospital Course|2266,2273|false|false|false|C0009818|Consultation|consult
Event|Event|Hospital Course|2274,2285|false|false|false|||appreciated
Event|Event|Hospital Course|2289,2293|false|false|false|||felt
Event|Event|Hospital Course|2308,2316|false|false|false|||standing
Event|Event|Hospital Course|2319,2330|false|false|false|||recommended
Finding|Gene or Genome|Hospital Course|2331,2334|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Pharmacologic Substance|Hospital Course|2335,2352|false|false|false|C0003364|Antihypertensive Agents|antihypertensives
Event|Event|Hospital Course|2335,2352|false|false|false|||antihypertensives
Event|Event|Hospital Course|2358,2367|false|false|false|||cautioned
Event|Event|Hospital Course|2385,2393|false|false|false|||pressure
Finding|Finding|Hospital Course|2385,2393|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|Hospital Course|2385,2393|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|Hospital Course|2385,2393|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|Hospital Course|2385,2393|false|false|false|C0033095||pressure
Finding|Finding|Hospital Course|2394,2401|false|false|false|C4036057|Too low|too low
Event|Event|Hospital Course|2398,2401|false|false|false|||low
Finding|Finding|Hospital Course|2398,2401|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Hospital Course|2398,2401|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Finding|Hospital Course|2402,2413|false|false|false|C4036056|Too quickly|too quickly
Finding|Idea or Concept|Hospital Course|2417,2425|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|Hospital Course|2417,2432|false|false|false|C0488549||Hospital course
Finding|Finding|Hospital Course|2417,2432|false|false|false|C0489547|Hospital course|Hospital course
Event|Event|Hospital Course|2426,2432|false|false|false|||course
Event|Event|Hospital Course|2447,2459|false|false|false|||unremarkable
Finding|Idea or Concept|Hospital Course|2469,2472|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|2469,2472|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|2477,2486|false|false|false|||discharge
Finding|Body Substance|Hospital Course|2477,2486|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|2477,2486|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|2477,2486|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|2477,2486|false|false|false|C0030685|Patient Discharge|discharge
Finding|Body Substance|Hospital Course|2491,2498|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|2491,2498|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|2491,2498|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|2503,2511|false|false|false|||afebrile
Finding|Finding|Hospital Course|2503,2511|false|false|false|C0277797|Apyrexial|afebrile
Event|Event|Hospital Course|2517,2523|false|false|false|||stable
Finding|Intellectual Product|Hospital Course|2517,2523|false|false|false|C1547311|Patient Condition Code - Stable|stable
Drug|Food|Hospital Course|2524,2529|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|vital
Attribute|Clinical Attribute|Hospital Course|2524,2535|false|false|false|C0488614;C0518766|Vital signs|vital signs
Procedure|Health Care Activity|Hospital Course|2524,2535|false|false|false|C0150404|Taking vital signs|vital signs
Event|Event|Hospital Course|2530,2535|false|false|false|||signs
Finding|Finding|Hospital Course|2530,2535|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Hospital Course|2530,2535|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Event|Event|Hospital Course|2538,2549|false|false|false|||comfortable
Finding|Finding|Hospital Course|2538,2549|false|false|false|C5546696|Feeling comfortable|comfortable
Anatomy|Body Space or Junction|Hospital Course|2553,2557|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|2553,2557|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|2553,2557|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|2553,2557|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Sign or Symptom|Hospital Course|2553,2562|false|false|false|C0221776|Oral pain|oral pain
Attribute|Clinical Attribute|Hospital Course|2558,2562|false|false|false|C2598155||pain
Event|Event|Hospital Course|2558,2562|false|false|false|||pain
Finding|Functional Concept|Hospital Course|2558,2562|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|2558,2562|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Hospital Course|2558,2570|false|false|false|C5548091|Demonstrates adequate pain control|pain control
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2558,2570|false|false|false|C0002766;C1304888|Pain control;Pain management (procedure)|pain control
Drug|Organic Chemical|Hospital Course|2563,2570|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|Hospital Course|2563,2570|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|Hospital Course|2563,2570|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Event|Event|Hospital Course|2563,2570|false|false|false|||control
Finding|Conceptual Entity|Hospital Course|2563,2570|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|Hospital Course|2563,2570|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|Hospital Course|2563,2570|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Event|Event|Hospital Course|2575,2585|false|false|false|||tolerating
Finding|Daily or Recreational Activity|Hospital Course|2588,2600|false|false|false|C0184625||regular diet
Drug|Food|Hospital Course|2596,2600|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|Hospital Course|2596,2600|false|false|false|||diet
Finding|Functional Concept|Hospital Course|2596,2600|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|Hospital Course|2596,2600|false|false|false|C0012159|Diet therapy|diet
Event|Event|Hospital Course|2605,2614|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|2605,2614|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|2605,2614|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|2605,2614|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|2605,2614|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|2605,2626|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|2615,2626|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|2615,2626|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|2615,2626|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|2615,2626|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|2631,2644|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|2631,2644|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Hospital Course|2631,2644|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|2631,2644|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|Hospital Course|2659,2662|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|2663,2667|false|false|false|C2598155||pain
Event|Event|Hospital Course|2663,2667|false|false|false|||pain
Finding|Functional Concept|Hospital Course|2663,2667|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|2663,2667|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|2669,2673|false|false|false|||temp
Finding|Gene or Genome|Hospital Course|2669,2673|false|false|false|C1823816|C1orf210 gene|temp
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2669,2673|false|false|false|C0279848|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|temp
Event|Event|Hospital Course|2682,2690|false|false|false|||headache
Finding|Sign or Symptom|Hospital Course|2682,2690|false|false|false|C0018681|Headache|headache
Drug|Organic Chemical|Hospital Course|2695,2706|false|false|false|C0002144|allopurinol|Allopurinol
Drug|Pharmacologic Substance|Hospital Course|2695,2706|false|false|false|C0002144|allopurinol|Allopurinol
Drug|Organic Chemical|Hospital Course|2727,2737|false|false|false|C0127615|mesalamine|Mesalamine
Drug|Pharmacologic Substance|Hospital Course|2727,2737|false|false|false|C0127615|mesalamine|Mesalamine
Event|Event|Hospital Course|2752,2755|false|false|false|||TID
Drug|Organic Chemical|Hospital Course|2760,2770|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|Hospital Course|2760,2770|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|Hospital Course|2760,2779|false|false|false|C0700548|metoprolol tartrate|Metoprolol Tartrate
Drug|Pharmacologic Substance|Hospital Course|2760,2779|false|false|false|C0700548|metoprolol tartrate|Metoprolol Tartrate
Drug|Organic Chemical|Hospital Course|2771,2779|false|false|false|C0039328;C0144544|Tartrates;tartrate|Tartrate
Drug|Pharmacologic Substance|Hospital Course|2771,2779|false|false|false|C0039328;C0144544|Tartrates;tartrate|Tartrate
Event|Event|Hospital Course|2771,2779|false|false|false|||Tartrate
Disorder|Mental or Behavioral Dysfunction|Hospital Course|2789,2792|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|2789,2792|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|2789,2792|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|2789,2792|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|2789,2792|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|2797,2807|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Pharmacologic Substance|Hospital Course|2797,2807|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Hazardous or Poisonous Substance|Hospital Course|2827,2835|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|Hospital Course|2827,2835|false|false|false|C0043031|warfarin|Warfarin
Drug|Pharmacologic Substance|Hospital Course|2827,2835|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|Hospital Course|2854,2863|false|false|false|C0030049|oxycodone|OxycoDONE
Drug|Pharmacologic Substance|Hospital Course|2854,2863|false|false|false|C0030049|oxycodone|OxycoDONE
Event|Event|Hospital Course|2854,2863|false|false|false|||OxycoDONE
Procedure|Laboratory Procedure|Hospital Course|2854,2863|false|false|false|C0524222|Oxycodone measurement|OxycoDONE
Finding|Idea or Concept|Hospital Course|2865,2874|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Finding|Intellectual Product|Hospital Course|2865,2874|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Drug|Biomedical or Dental Material|Hospital Course|2865,2882|false|false|false|C1708470|Immediate Release Dosage Form|Immediate Release
Event|Event|Hospital Course|2875,2882|false|false|false|||Release
Finding|Functional Concept|Hospital Course|2875,2882|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|2875,2882|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2875,2882|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Finding|Gene or Genome|Hospital Course|2901,2904|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|2905,2909|false|false|false|C2598155||pain
Event|Event|Hospital Course|2905,2909|false|false|false|||pain
Finding|Functional Concept|Hospital Course|2905,2909|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|2905,2909|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|2914,2922|false|false|false|C0012010|diazepam|Diazepam
Drug|Pharmacologic Substance|Hospital Course|2914,2922|false|false|false|C0012010|diazepam|Diazepam
Finding|Gene or Genome|Hospital Course|2936,2939|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|2940,2946|false|false|false|||spasms
Finding|Sign or Symptom|Hospital Course|2940,2946|false|false|false|C0037763|Spasm|spasms
Event|Event|Hospital Course|2951,2960|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|2951,2960|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|2951,2960|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|2951,2960|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|2951,2960|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|2951,2972|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|2951,2972|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|2961,2972|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|2961,2972|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|2961,2972|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|Hospital Course|2974,2978|false|false|false|||Home
Finding|Idea or Concept|Hospital Course|2974,2978|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|2974,2978|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|2974,2978|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|Hospital Course|2984,2991|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|Hospital Course|2984,2991|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|Hospital Course|2994,3002|false|false|false|||Facility
Finding|Intellectual Product|Hospital Course|2994,3002|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|Hospital Course|3010,3019|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|3010,3019|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|3010,3019|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|3010,3019|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|3010,3019|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|3010,3029|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|3020,3029|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|3020,3029|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|3020,3029|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|3020,3029|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|3020,3029|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Injury or Poisoning|Hospital Course|3034,3042|false|false|false|C0016658|Fracture|fracture
Event|Event|Hospital Course|3034,3042|false|false|false|||fracture
Finding|Mental Process|Discharge Condition|3066,3072|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|3066,3079|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|3066,3079|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|3073,3079|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|3073,3079|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|3081,3086|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|3081,3086|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|3091,3099|false|false|false|||coherent
Finding|Finding|Discharge Condition|3091,3099|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|3101,3106|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|3101,3123|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|3101,3123|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|3110,3123|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|3110,3123|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|3110,3123|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|3125,3130|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|3125,3130|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|3125,3130|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|3125,3130|false|false|false|||Alert
Finding|Finding|Discharge Condition|3125,3130|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|3125,3130|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|3125,3130|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|3135,3146|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|3135,3146|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|3148,3156|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|3148,3156|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|3148,3156|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|3157,3163|false|false|false|C5889824||Status
Event|Event|Discharge Condition|3157,3163|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|3157,3163|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|3165,3175|false|false|false|||Ambulatory
Finding|Functional Concept|Discharge Condition|3165,3175|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|3165,3175|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|3165,3175|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|3165,3175|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|3178,3189|false|false|false|||Independent
Finding|Finding|Discharge Condition|3178,3189|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Condition|3178,3189|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Event|Event|Discharge Instructions|3226,3235|false|false|false|||undergone
Event|Activity|Discharge Instructions|3250,3259|false|false|false|C3241922|Operation Activity|operation
Event|Event|Discharge Instructions|3250,3259|false|false|false|||operation
Procedure|Machine Activity|Discharge Instructions|3250,3259|false|false|false|C0543467;C1880161|Computer Operation;Operative Surgical Procedures|operation
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|3250,3259|false|false|false|C0543467;C1880161|Computer Operation;Operative Surgical Procedures|operation
Disorder|Disease or Syndrome|Discharge Instructions|3261,3269|false|false|false|C0751437|Adenohypophyseal Diseases|Anterior
Anatomy|Body Location or Region|Discharge Instructions|3270,3278|false|false|false|C0027530|Neck|Cervical
Event|Event|Discharge Instructions|3280,3293|false|false|false|||Decompression
Finding|Functional Concept|Discharge Instructions|3280,3293|false|false|false|C1965697|Decompression - action (qualifier value)|Decompression
Phenomenon|Phenomenon or Process|Discharge Instructions|3280,3293|false|false|false|C0011117|external decompression|Decompression
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|3280,3293|false|false|false|C0021153;C1829459|Decompression;Decompressive incision|Decompression
Event|Event|Discharge Instructions|3298,3304|false|false|false|||Fusion
Finding|Functional Concept|Discharge Instructions|3298,3304|false|false|false|C0332466|Fused structure|Fusion
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|3298,3304|false|false|false|C1293131|Fusion procedure|Fusion
Event|Activity|Discharge Instructions|3328,3337|false|false|false|C3241922|Operation Activity|operation
Event|Event|Discharge Instructions|3328,3337|false|false|false|||operation
Procedure|Machine Activity|Discharge Instructions|3328,3337|false|false|false|C0543467;C1880161|Computer Operation;Operative Surgical Procedures|operation
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|3328,3337|false|false|false|C0543467;C1880161|Computer Operation;Operative Surgical Procedures|operation
Event|Activity|Discharge Instructions|3340,3348|false|false|false|C0441655|Activities|Activity
Event|Event|Discharge Instructions|3340,3348|false|false|false|||Activity
Finding|Daily or Recreational Activity|Discharge Instructions|3340,3348|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Instructions|3340,3348|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Event|Event|Discharge Instructions|3365,3369|true|false|false|||lift
Procedure|Laboratory Procedure|Discharge Instructions|3394,3397|true|false|false|C3161851|liquid-based cytology (procedure)|lbs
Event|Event|Discharge Instructions|3429,3440|false|false|false|||comfortable
Finding|Finding|Discharge Instructions|3429,3440|false|false|false|C5546696|Feeling comfortable|comfortable
Event|Event|Discharge Instructions|3455,3458|true|false|false|||sit
Anatomy|Cell Component|Discharge Instructions|3464,3467|true|false|false|C1166663|actomyosin contractile ring|car
Disorder|Disease or Syndrome|Discharge Instructions|3464,3467|true|false|false|C0406810|Carney Complex|car
Drug|Amino Acid, Peptide, or Protein|Discharge Instructions|3464,3467|true|false|false|C3539542;C4039583;C5890846|Chimeric antigen receptor;Coxsackievirus and Adenovirus Receptor, human;Extracellular Calcium-Sensing Receptor, Human|car
Drug|Biologically Active Substance|Discharge Instructions|3464,3467|true|false|false|C3539542;C4039583;C5890846|Chimeric antigen receptor;Coxsackievirus and Adenovirus Receptor, human;Extracellular Calcium-Sensing Receptor, Human|car
Drug|Immunologic Factor|Discharge Instructions|3464,3467|true|false|false|C3539542;C4039583;C5890846|Chimeric antigen receptor;Coxsackievirus and Adenovirus Receptor, human;Extracellular Calcium-Sensing Receptor, Human|car
Finding|Gene or Genome|Discharge Instructions|3464,3467|true|false|false|C1413828;C1417827;C1420354;C1547285;C1706434;C1858724;C2239319;C3273602;C3540475;C3811749;C4039583;C5890846;C5890847;C5960871|CASR wt Allele;CXADR gene;CXADR wt Allele;CXADRP1 gene;Car - Mode of Arrival Code;Caronte Gene;Chimeric antigen receptor;Extracellular Calcium-Sensing Receptor, Human;NR1I3 gene;NR1I3 wt Allele;PRKAR1A wt Allele;SPG7 gene;SPG7 wt Allele;TRIM13 wt Allele|car
Finding|Intellectual Product|Discharge Instructions|3464,3467|true|false|false|C1413828;C1417827;C1420354;C1547285;C1706434;C1858724;C2239319;C3273602;C3540475;C3811749;C4039583;C5890846;C5890847;C5960871|CASR wt Allele;CXADR gene;CXADR wt Allele;CXADRP1 gene;Car - Mode of Arrival Code;Caronte Gene;Chimeric antigen receptor;Extracellular Calcium-Sensing Receptor, Human;NR1I3 gene;NR1I3 wt Allele;PRKAR1A wt Allele;SPG7 gene;SPG7 wt Allele;TRIM13 wt Allele|car
Finding|Receptor|Discharge Instructions|3464,3467|true|false|false|C1413828;C1417827;C1420354;C1547285;C1706434;C1858724;C2239319;C3273602;C3540475;C3811749;C4039583;C5890846;C5890847;C5960871|CASR wt Allele;CXADR gene;CXADR wt Allele;CXADRP1 gene;Car - Mode of Arrival Code;Caronte Gene;Chimeric antigen receptor;Extracellular Calcium-Sensing Receptor, Human;NR1I3 gene;NR1I3 wt Allele;PRKAR1A wt Allele;SPG7 gene;SPG7 wt Allele;TRIM13 wt Allele|car
Event|Event|Discharge Instructions|3472,3477|true|false|false|||chair
Event|Event|Discharge Instructions|3528,3535|true|false|false|||walking
Event|Event|Discharge Instructions|3546,3560|false|false|false|||Rehabilitation
Finding|Finding|Discharge Instructions|3546,3560|false|false|false|C0007237;C0034992|Encounter due to care involving use of rehabilitation procedures;Rehabilitation aspects|Rehabilitation
Finding|Functional Concept|Discharge Instructions|3546,3560|false|false|false|C0007237;C0034992|Encounter due to care involving use of rehabilitation procedures;Rehabilitation aspects|Rehabilitation
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|3546,3560|false|false|false|C0034991|Rehabilitation therapy|Rehabilitation
Finding|Finding|Discharge Instructions|3562,3570|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|Discharge Instructions|3562,3570|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|Discharge Instructions|3562,3570|false|false|false|C0031809|Physical Examination|Physical
Finding|Intellectual Product|Discharge Instructions|3562,3578|false|false|false|C1547999|Diagnostic Service Section ID - Physical Therapy|Physical Therapy
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|3562,3578|false|false|false|C0949766|Physical therapy|Physical Therapy
Event|Event|Discharge Instructions|3571,3578|false|false|false|||Therapy
Finding|Finding|Discharge Instructions|3571,3578|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|Therapy
Finding|Functional Concept|Discharge Instructions|3571,3578|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|Therapy
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|3571,3578|false|false|false|C0087111|Therapeutic procedure|Therapy
Finding|Finding|Discharge Instructions|3584,3591|false|false|false|C4035626|3 times|3 times
Disorder|Disease or Syndrome|Discharge Instructions|3586,3591|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Event|Event|Discharge Instructions|3586,3591|false|false|false|||times
Finding|Idea or Concept|Discharge Instructions|3594,3597|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Discharge Instructions|3594,3597|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Discharge Instructions|3618,3622|false|false|false|||walk
Finding|Daily or Recreational Activity|Discharge Instructions|3618,3622|false|false|false|C0080331|Walking (function)|walk
Event|Event|Discharge Instructions|3643,3647|false|false|false|||part
Finding|Idea or Concept|Discharge Instructions|3643,3647|false|false|false|C1552020|Role Class - part|part
Event|Activity|Discharge Instructions|3656,3664|false|false|false|C0237820||recovery
Event|Event|Discharge Instructions|3656,3664|false|false|false|||recovery
Finding|Organism Function|Discharge Instructions|3656,3664|false|false|false|C2004454|Recovery - healing process|recovery
Event|Event|Discharge Instructions|3675,3679|false|false|false|||walk
Finding|Finding|Discharge Instructions|3683,3687|false|false|false|C4281574|Much|much
Event|Event|Discharge Instructions|3700,3708|false|false|false|||tolerate
Finding|Conceptual Entity|Discharge Instructions|3723,3732|false|false|false|C0231448;C1880641|Extension;Telephone Extension Number|Extension
Finding|Functional Concept|Discharge Instructions|3723,3732|false|false|false|C0231448;C1880641|Extension;Telephone Extension Number|Extension
Event|Event|Discharge Instructions|3733,3741|false|false|false|||Exercise
Finding|Daily or Recreational Activity|Discharge Instructions|3733,3741|false|false|false|C0015259|Exercise|Exercise
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|3733,3741|false|false|false|C1522704|Exercise Pain Management|Exercise
Finding|Idea or Concept|Discharge Instructions|3760,3763|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Discharge Instructions|3760,3763|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Discharge Instructions|3769,3777|false|false|false|||xercises
Event|Event|Discharge Instructions|3781,3791|false|false|false|||instructed
Attribute|Clinical Attribute|Discharge Instructions|3795,3805|false|false|false|C2598159||Swallowing
Event|Event|Discharge Instructions|3795,3805|false|false|false|||Swallowing
Finding|Finding|Discharge Instructions|3795,3805|false|false|false|C0011167;C0740170;C4281783|Deglutition;Does swallow;Swallowing G-code|Swallowing
Finding|Intellectual Product|Discharge Instructions|3795,3805|false|false|false|C0011167;C0740170;C4281783|Deglutition;Does swallow;Swallowing G-code|Swallowing
Finding|Organism Function|Discharge Instructions|3795,3805|false|false|false|C0011167;C0740170;C4281783|Deglutition;Does swallow;Swallowing G-code|Swallowing
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|3795,3805|false|false|false|C3665547|outcomes otolaryngology swallowing (treatment)|Swallowing
Finding|Finding|Discharge Instructions|3807,3817|true|false|false|C1299586|Has difficulty doing (qualifier value)|Difficulty
Disorder|Disease or Syndrome|Discharge Instructions|3807,3828|true|false|false|C0011168|Deglutition Disorders|Difficulty swallowing
Attribute|Clinical Attribute|Discharge Instructions|3818,3828|true|false|false|C2598159||swallowing
Event|Event|Discharge Instructions|3818,3828|true|false|false|||swallowing
Finding|Finding|Discharge Instructions|3818,3828|true|false|false|C0011167;C0740170;C4281783|Deglutition;Does swallow;Swallowing G-code|swallowing
Finding|Intellectual Product|Discharge Instructions|3818,3828|true|false|false|C0011167;C0740170;C4281783|Deglutition;Does swallow;Swallowing G-code|swallowing
Finding|Organism Function|Discharge Instructions|3818,3828|true|false|false|C0011167;C0740170;C4281783|Deglutition;Does swallow;Swallowing G-code|swallowing
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|3818,3828|true|false|false|C3665547|outcomes otolaryngology swallowing (treatment)|swallowing
Event|Event|Discharge Instructions|3836,3844|true|false|false|||uncommon
Event|Event|Discharge Instructions|3857,3861|true|false|false|||type
Finding|Gene or Genome|Discharge Instructions|3857,3861|true|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Intellectual Product|Discharge Instructions|3857,3861|true|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Event|Event|Discharge Instructions|3865,3872|true|false|false|||surgery
Finding|Finding|Discharge Instructions|3865,3872|true|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Discharge Instructions|3865,3872|true|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Discharge Instructions|3865,3872|true|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|3865,3872|true|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Event|Discharge Instructions|3886,3893|false|false|false|||resolve
Finding|Finding|Discharge Instructions|3899,3903|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Discharge Instructions|3899,3903|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Discharge Instructions|3899,3903|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Disorder|Injury or Poisoning|Discharge Instructions|3925,3930|false|false|false|C0005658|bite injury|bites
Event|Event|Discharge Instructions|3925,3930|false|false|false|||bites
Event|Event|Discharge Instructions|3935,3938|false|false|false|||eat
Event|Event|Discharge Instructions|3948,3956|false|false|false|||Removing
Event|Event|Discharge Instructions|3961,3967|false|false|false|||collar
Event|Event|Discharge Instructions|3974,3980|false|false|false|||eating
Event|Event|Discharge Instructions|3989,3996|false|false|false|||helpful
Event|Event|Discharge Instructions|4015,4020|false|false|false|||limit
Event|Event|Discharge Instructions|4026,4034|false|false|false|||movement
Finding|Organism Function|Discharge Instructions|4026,4034|false|false|false|C0026649|Movement|movement
Anatomy|Body Location or Region|Discharge Instructions|4044,4048|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|Discharge Instructions|4044,4048|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|Discharge Instructions|4044,4048|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Event|Event|Discharge Instructions|4056,4062|false|false|false|||remove
Event|Event|Discharge Instructions|4068,4074|false|false|false|||collar
Event|Event|Discharge Instructions|4081,4087|false|false|false|||eating
Anatomy|Body Location or Region|Discharge Instructions|4091,4099|false|false|false|C0027530|Neck|Cervical
Anatomy|Body Location or Region|Discharge Instructions|4109,4113|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|Discharge Instructions|4109,4113|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|Discharge Instructions|4109,4113|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|Discharge Instructions|4114,4119|false|false|false|||Brace
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|4114,4119|false|false|false|C1828220|Application of brace (procedure)|Brace
Event|Event|Discharge Instructions|4125,4129|false|false|false|||need
Event|Event|Discharge Instructions|4133,4137|false|false|false|||wear
Event|Event|Discharge Instructions|4142,4147|false|false|false|||brace
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|4142,4147|false|false|false|C1828220|Application of brace (procedure)|brace
Disorder|Disease or Syndrome|Discharge Instructions|4156,4161|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Event|Event|Discharge Instructions|4156,4161|false|false|false|||times
Event|Event|Discharge Instructions|4173,4179|false|false|false|||follow
Finding|Functional Concept|Discharge Instructions|4173,4179|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|Discharge Instructions|4173,4179|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|Discharge Instructions|4173,4182|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|Discharge Instructions|4173,4182|false|false|false|C1522577|follow-up|follow-up
Event|Activity|Discharge Instructions|4183,4194|false|false|false|C0003629|Appointments|appointment
Event|Event|Discharge Instructions|4183,4194|false|false|false|||appointment
Event|Event|Discharge Instructions|4233,4239|false|false|false|||remove
Event|Event|Discharge Instructions|4254,4258|false|false|false|||take
Finding|Daily or Recreational Activity|Discharge Instructions|4254,4267|false|false|false|C2937301|take a shower|take a shower
Event|Event|Discharge Instructions|4261,4267|false|false|false|||shower
Event|Event|Discharge Instructions|4270,4275|false|false|false|||Limit
Event|Event|Discharge Instructions|4282,4288|false|false|false|||motion
Phenomenon|Natural Phenomenon or Process|Discharge Instructions|4282,4288|false|false|false|C0026597|Motion|motion
Anatomy|Body Location or Region|Discharge Instructions|4297,4301|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|Discharge Instructions|4297,4301|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|Discharge Instructions|4297,4301|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Event|Activity|Discharge Instructions|4327,4332|false|false|false|C1882509|put - instruction imperative|Place
Event|Event|Discharge Instructions|4327,4332|false|false|false|||Place
Finding|Functional Concept|Discharge Instructions|4327,4332|false|false|false|C1704765|Place - dosing instruction imperative|Place
Procedure|Health Care Activity|Discharge Instructions|4327,4332|false|false|false|C1533810||Place
Event|Event|Discharge Instructions|4345,4349|false|false|false|||back
Anatomy|Body Location or Region|Discharge Instructions|4358,4362|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|Discharge Instructions|4358,4362|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|Discharge Instructions|4358,4362|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Disorder|Injury or Poisoning|Discharge Instructions|4395,4400|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|Wound
Event|Event|Discharge Instructions|4395,4400|false|false|false|||Wound
Finding|Body Substance|Discharge Instructions|4395,4400|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|Wound
Finding|Functional Concept|Discharge Instructions|4395,4400|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|Wound
Finding|Intellectual Product|Discharge Instructions|4395,4400|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|Wound
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|4395,4405|false|false|false|C0886052;C1272654|Wound care management;wound care|Wound Care
Event|Activity|Discharge Instructions|4401,4405|false|false|false|C1947933|care activity|Care
Event|Event|Discharge Instructions|4401,4405|false|false|false|||Care
Finding|Finding|Discharge Instructions|4401,4405|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Discharge Instructions|4401,4405|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Disorder|Injury or Poisoning|Discharge Instructions|4415,4425|false|false|false|C0043246|Laceration|laceration
Event|Event|Discharge Instructions|4415,4425|false|false|false|||laceration
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|4429,4434|false|false|false|C0036270|Scalp structure|scalp
Event|Event|Discharge Instructions|4439,4447|false|false|false|||drainage
Finding|Body Substance|Discharge Instructions|4439,4447|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|Discharge Instructions|4439,4447|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|4439,4447|false|false|false|C0013103|Drainage procedure|drainage
Disorder|Disease or Syndrome|Discharge Instructions|4448,4455|false|false|false|C0041834|Erythema|redness
Event|Event|Discharge Instructions|4448,4455|false|false|false|||redness
Finding|Finding|Discharge Instructions|4448,4455|false|false|false|C0332575|Redness|redness
Disorder|Disease or Syndrome|Discharge Instructions|4464,4467|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|Discharge Instructions|4464,4467|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|Discharge Instructions|4464,4467|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|Discharge Instructions|4464,4467|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|Discharge Instructions|4464,4467|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|Discharge Instructions|4464,4467|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|Discharge Instructions|4464,4467|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|Discharge Instructions|4464,4467|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|Discharge Instructions|4464,4467|false|false|false|||PCP
Finding|Gene or Genome|Discharge Instructions|4464,4467|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|Discharge Instructions|4464,4467|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|Discharge Instructions|4472,4476|false|false|false|||take
Event|Event|Discharge Instructions|4483,4490|false|false|false|||staples
Event|Event|Discharge Instructions|4509,4515|false|false|false|||resume
Event|Event|Discharge Instructions|4516,4522|false|false|false|||taking
Finding|Idea or Concept|Discharge Instructions|4535,4539|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Discharge Instructions|4535,4539|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Discharge Instructions|4535,4539|false|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|Discharge Instructions|4540,4551|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|4540,4551|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|4540,4551|false|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|4540,4551|false|false|false|C4284232|Medications|medications
Finding|Functional Concept|Discharge Instructions|4580,4590|false|false|false|C1524062|Additional|Additional
Attribute|Clinical Attribute|Discharge Instructions|4591,4602|false|false|true|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Discharge Instructions|4591,4602|false|false|true|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Discharge Instructions|4591,4602|false|false|false|||Medications
Finding|Intellectual Product|Discharge Instructions|4591,4602|false|false|true|C4284232|Medications|Medications
Drug|Organic Chemical|Discharge Instructions|4606,4613|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|Discharge Instructions|4606,4613|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|Discharge Instructions|4606,4613|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Event|Event|Discharge Instructions|4606,4613|false|false|false|||control
Finding|Conceptual Entity|Discharge Instructions|4606,4613|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|Discharge Instructions|4606,4613|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|Discharge Instructions|4606,4613|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Attribute|Clinical Attribute|Discharge Instructions|4620,4624|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|4620,4624|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|4620,4624|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|4620,4624|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Discharge Instructions|4634,4639|false|false|false|||allow
Event|Event|Discharge Instructions|4653,4659|false|false|false|||refill
Finding|Idea or Concept|Discharge Instructions|4653,4659|false|false|false|C0807726|refill|refill
Drug|Hazardous or Poisonous Substance|Discharge Instructions|4663,4671|false|false|false|C0027415|Narcotics|narcotic
Drug|Pharmacologic Substance|Discharge Instructions|4663,4671|false|false|false|C0027415|Narcotics|narcotic
Event|Event|Discharge Instructions|4663,4671|false|false|false|||narcotic
Attribute|Clinical Attribute|Discharge Instructions|4673,4686|false|false|false|C2741652||prescriptions
Event|Event|Discharge Instructions|4673,4686|false|false|false|||prescriptions
Procedure|Health Care Activity|Discharge Instructions|4673,4686|false|false|false|C0033080|Prescription (procedure)|prescriptions
Disorder|Disease or Syndrome|Discharge Instructions|4691,4695|false|false|false|C0270724|Infantile Neuroaxonal Dystrophy|plan
Event|Event|Discharge Instructions|4691,4695|false|false|false|||plan
Finding|Functional Concept|Discharge Instructions|4691,4695|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Intellectual Product|Discharge Instructions|4691,4695|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Mental Process|Discharge Instructions|4691,4695|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Event|Event|Discharge Instructions|4729,4735|false|false|false|||mailed
Event|Event|Discharge Instructions|4745,4749|false|false|false|||home
Finding|Idea or Concept|Discharge Instructions|4745,4749|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Discharge Instructions|4745,4749|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Discharge Instructions|4745,4749|false|false|false|C1553498|home health encounter|home
Event|Event|Discharge Instructions|4753,4757|false|false|false|||pick
Event|Event|Discharge Instructions|4809,4816|true|false|false|||allowed
Event|Event|Discharge Instructions|4820,4824|true|false|false|||call
Drug|Hazardous or Poisonous Substance|Discharge Instructions|4828,4836|true|false|false|C0027415|Narcotics|narcotic
Drug|Pharmacologic Substance|Discharge Instructions|4828,4836|true|false|false|C0027415|Narcotics|narcotic
Event|Event|Discharge Instructions|4828,4836|true|false|false|||narcotic
Drug|Organic Chemical|Discharge Instructions|4838,4847|true|false|false|C0722364|Oxycontin|oxycontin
Drug|Pharmacologic Substance|Discharge Instructions|4838,4847|true|false|false|C0722364|Oxycontin|oxycontin
Event|Event|Discharge Instructions|4838,4847|true|false|false|||oxycontin
Drug|Organic Chemical|Discharge Instructions|4849,4858|false|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|Discharge Instructions|4849,4858|false|false|false|C0030049|oxycodone|oxycodone
Event|Event|Discharge Instructions|4849,4858|false|false|false|||oxycodone
Procedure|Laboratory Procedure|Discharge Instructions|4849,4858|false|false|false|C0524222|Oxycodone measurement|oxycodone
Drug|Organic Chemical|Discharge Instructions|4861,4869|false|false|false|C0086787|Percocet|percocet
Drug|Pharmacologic Substance|Discharge Instructions|4861,4869|false|false|false|C0086787|Percocet|percocet
Event|Event|Discharge Instructions|4861,4869|false|false|false|||percocet
Attribute|Clinical Attribute|Discharge Instructions|4871,4884|false|false|false|C2741652||prescriptions
Event|Event|Discharge Instructions|4871,4884|false|false|false|||prescriptions
Procedure|Health Care Activity|Discharge Instructions|4871,4884|false|false|false|C0033080|Prescription (procedure)|prescriptions
Event|Event|Discharge Instructions|4892,4900|false|false|false|||pharmacy
Finding|Intellectual Product|Discharge Instructions|4892,4900|false|false|false|C1547997;C3244303|Diagnostic Service Section ID - Pharmacy;Pharmacy domain|pharmacy
Procedure|Health Care Activity|Discharge Instructions|4892,4900|false|false|false|C0031321|Pharmaceutical Services|pharmacy
Finding|Functional Concept|Discharge Instructions|4907,4915|false|false|false|C0332287;C1883712|Add - instruction imperative;In addition to|addition
Event|Event|Discharge Instructions|4930,4937|false|false|false|||allowed
Event|Event|Discharge Instructions|4941,4946|false|false|false|||write
Attribute|Clinical Attribute|Discharge Instructions|4951,4955|false|false|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|4951,4955|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|4951,4955|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|Discharge Instructions|4956,4967|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|4956,4967|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|4956,4967|false|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|4956,4967|false|false|false|C4284232|Medications|medications
Event|Event|Discharge Instructions|4998,5005|false|false|false|||surgery
Finding|Finding|Discharge Instructions|4998,5005|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Discharge Instructions|4998,5005|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Discharge Instructions|4998,5005|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|4998,5005|false|false|false|C0543467|Operative Surgical Procedures|surgery
Finding|Functional Concept|Discharge Instructions|5009,5015|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|Follow
Finding|Intellectual Product|Discharge Instructions|5009,5015|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|Follow
Finding|Finding|Discharge Instructions|5009,5018|false|false|false|C0589120|Follow-up status|Follow up
Procedure|Health Care Activity|Discharge Instructions|5009,5018|false|false|false|C1522577|follow-up|Follow up
Event|Event|Discharge Instructions|5016,5018|false|false|false|||up
Event|Event|Discharge Instructions|5028,5032|false|false|false|||Call
Event|Event|Discharge Instructions|5037,5043|false|false|false|||office
Finding|Idea or Concept|Discharge Instructions|5037,5043|false|false|false|C1549636|Address type - Office|office
Event|Activity|Discharge Instructions|5060,5071|false|false|false|C0003629|Appointments|appointment
Event|Event|Discharge Instructions|5060,5071|false|false|false|||appointment
Finding|Idea or Concept|Discharge Instructions|5104,5107|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Discharge Instructions|5104,5107|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Activity|Discharge Instructions|5116,5125|false|false|false|C3241922|Operation Activity|operation
Event|Event|Discharge Instructions|5116,5125|false|false|false|||operation
Procedure|Machine Activity|Discharge Instructions|5116,5125|false|false|false|C0543467;C1880161|Computer Operation;Operative Surgical Procedures|operation
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|5116,5125|false|false|false|C0543467;C1880161|Computer Operation;Operative Surgical Procedures|operation
Finding|Intellectual Product|Discharge Instructions|5172,5176|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|Discharge Instructions|5177,5182|false|false|false|||visit
Finding|Social Behavior|Discharge Instructions|5177,5182|false|false|false|C0545082|Visit|visit
Event|Event|Discharge Instructions|5191,5196|false|false|false|||check
Anatomy|Body Location or Region|Discharge Instructions|5202,5210|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Discharge Instructions|5202,5210|false|false|false|C0332803|Surgical wound|incision
Event|Event|Discharge Instructions|5202,5210|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|5202,5210|false|false|false|C0184898|Surgical incisions|incision
Drug|Biomedical or Dental Material|Discharge Instructions|5217,5225|true|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|Discharge Instructions|5217,5225|true|false|false|||baseline
Finding|Idea or Concept|Discharge Instructions|5217,5225|true|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Phenomenon|Natural Phenomenon or Process|Discharge Instructions|5227,5233|true|false|false|C0043309|Roentgen Rays|x rays
Procedure|Diagnostic Procedure|Discharge Instructions|5227,5233|true|false|false|C1306645|Plain x-ray|x rays
Event|Event|Discharge Instructions|5229,5233|true|false|false|||rays
Phenomenon|Natural Phenomenon or Process|Discharge Instructions|5229,5233|true|false|false|C0851346|Radiation|rays
Event|Event|Discharge Instructions|5238,5244|true|false|false|||answer
Event|Event|Discharge Instructions|5249,5258|true|false|false|||questions
Finding|Intellectual Product|Discharge Instructions|5269,5273|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|Discharge Instructions|5274,5277|false|false|false|||see
Finding|Idea or Concept|Discharge Instructions|5302,5305|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Discharge Instructions|5302,5305|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Activity|Discharge Instructions|5313,5322|false|false|false|C3241922|Operation Activity|operation
Event|Event|Discharge Instructions|5313,5322|false|false|false|||operation
Procedure|Machine Activity|Discharge Instructions|5313,5322|false|false|false|C0543467;C1880161|Computer Operation;Operative Surgical Procedures|operation
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|5313,5322|false|false|false|C0543467;C1880161|Computer Operation;Operative Surgical Procedures|operation
Finding|Finding|Discharge Instructions|5333,5337|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Discharge Instructions|5333,5337|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Discharge Instructions|5333,5337|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Discharge Instructions|5346,5357|false|false|false|C0750501|most likely|most likely
Finding|Finding|Discharge Instructions|5351,5357|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Discharge Instructions|5351,5357|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|Discharge Instructions|5358,5364|false|false|false|||obtain
Attribute|Clinical Attribute|Discharge Instructions|5365,5372|false|false|false|C1525443|W flexion|Flexion
Event|Event|Discharge Instructions|5365,5372|false|false|false|||Flexion
Finding|Organ or Tissue Function|Discharge Instructions|5365,5372|false|false|false|C0231452||Flexion
Finding|Conceptual Entity|Discharge Instructions|5373,5382|false|false|false|C0231448;C1880641|Extension;Telephone Extension Number|Extension
Finding|Functional Concept|Discharge Instructions|5373,5382|false|false|false|C0231448;C1880641|Extension;Telephone Extension Number|Extension
Drug|Pharmacologic Substance|Discharge Instructions|5383,5389|false|false|false|C0885876|X-rays, Homeopathic Preparations|X-rays
Event|Event|Discharge Instructions|5383,5389|false|false|false|||X-rays
Phenomenon|Natural Phenomenon or Process|Discharge Instructions|5383,5389|false|false|false|C0043309|Roentgen Rays|X-rays
Procedure|Diagnostic Procedure|Discharge Instructions|5383,5389|false|false|false|C0043299;C1306645|Diagnostic radiologic examination;Plain x-ray|X-rays
Finding|Intellectual Product|Discharge Instructions|5395,5400|false|false|false|C4050225|Often - answer to question|often
Event|Event|Discharge Instructions|5401,5405|false|false|false|||able
Finding|Finding|Discharge Instructions|5401,5405|false|false|false|C1299581|Able (qualifier value)|able
Event|Event|Discharge Instructions|5409,5414|false|false|false|||place
Disorder|Disease or Syndrome|Discharge Instructions|5424,5428|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|Discharge Instructions|5451,5455|false|false|false|||wean
Finding|Intellectual Product|Discharge Instructions|5471,5475|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|Discharge Instructions|5487,5491|false|false|false|||call
Event|Event|Discharge Instructions|5496,5502|false|false|false|||office
Finding|Idea or Concept|Discharge Instructions|5496,5502|false|false|false|C1549636|Address type - Office|office
Event|Event|Discharge Instructions|5517,5522|false|false|false|||fever
Finding|Finding|Discharge Instructions|5517,5522|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|Discharge Instructions|5517,5522|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|Discharge Instructions|5529,5536|false|false|false|||degrees
Finding|Intellectual Product|Discharge Instructions|5529,5536|false|false|false|C0542560|Academic degree|degrees
Event|Event|Discharge Instructions|5550,5558|true|false|false|||drainage
Finding|Body Substance|Discharge Instructions|5550,5558|true|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|Discharge Instructions|5550,5558|true|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|5550,5558|true|false|false|C0013103|Drainage procedure|drainage
Disorder|Injury or Poisoning|Discharge Instructions|5569,5574|true|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Event|Event|Discharge Instructions|5569,5574|true|false|false|||wound
Finding|Body Substance|Discharge Instructions|5569,5574|true|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|Discharge Instructions|5569,5574|true|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|Discharge Instructions|5569,5574|true|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Event|Event|Discharge Instructions|5588,5597|true|false|false|||questions
Event|Event|Discharge Instructions|5600,5608|false|false|false|||Physical
Finding|Finding|Discharge Instructions|5600,5608|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|Discharge Instructions|5600,5608|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|Discharge Instructions|5600,5608|false|false|false|C0031809|Physical Examination|Physical
Finding|Intellectual Product|Discharge Instructions|5600,5616|false|false|false|C1547999|Diagnostic Service Section ID - Physical Therapy|Physical Therapy
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|5600,5616|false|false|false|C0949766|Physical therapy|Physical Therapy
Event|Event|Discharge Instructions|5609,5616|false|false|false|||Therapy
Finding|Finding|Discharge Instructions|5609,5616|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|Therapy
Finding|Functional Concept|Discharge Instructions|5609,5616|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|Therapy
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|5609,5616|false|false|false|C0087111|Therapeutic procedure|Therapy
Event|Activity|Discharge Instructions|5618,5626|false|false|false|C0441655|Activities|activity
Event|Event|Discharge Instructions|5618,5626|false|false|false|||activity
Finding|Daily or Recreational Activity|Discharge Instructions|5618,5626|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Finding|Finding|Discharge Instructions|5618,5626|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Event|Event|Discharge Instructions|5630,5639|false|false|false|||tolerated
Finding|Finding|Discharge Instructions|5649,5658|false|false|false|C0682295|Full-time employment (finding)|full time
Event|Event|Discharge Instructions|5654,5658|false|false|false|||time
Finding|Finding|Discharge Instructions|5654,5658|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Discharge Instructions|5654,5658|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Discharge Instructions|5654,5658|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|Discharge Instructions|5676,5679|true|false|false|||use
Finding|Functional Concept|Discharge Instructions|5680,5690|true|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|ambulatory
Finding|Idea or Concept|Discharge Instructions|5680,5690|true|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|ambulatory
Finding|Intellectual Product|Discharge Instructions|5680,5690|true|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|ambulatory
Procedure|Health Care Activity|Discharge Instructions|5680,5690|true|false|false|C1561560|ambulatory encounter|ambulatory
Event|Event|Discharge Instructions|5701,5708|true|false|false|||devices
Event|Event|Discharge Instructions|5713,5719|true|false|false|||safety
Phenomenon|Human-caused Phenomenon or Process|Discharge Instructions|5713,5719|true|true|false|C0036043|Safety|safety
Disorder|Disease or Syndrome|Discharge Instructions|5724,5731|true|false|false|C0011119|Decompression Sickness|bending
Event|Event|Discharge Instructions|5724,5731|true|false|false|||bending
Finding|Finding|Discharge Instructions|5724,5731|true|false|false|C0700231;C2584296|Bending - Changing basic body position;Does bend|bending
Finding|Physiologic Function|Discharge Instructions|5724,5731|true|false|false|C0700231;C2584296|Bending - Changing basic body position;Does bend|bending
Event|Event|Discharge Instructions|5732,5740|true|false|false|||twisting
Finding|Pathologic Function|Discharge Instructions|5732,5740|true|false|false|C0040480;C1265748|Musculoskeletal torsion (function);Torsion (malposition)|twisting
Finding|Physiologic Function|Discharge Instructions|5732,5740|true|false|false|C0040480;C1265748|Musculoskeletal torsion (function);Torsion (malposition)|twisting
Event|Event|Discharge Instructions|5745,5752|true|false|false|||lifting
Event|Event|Discharge Instructions|5759,5768|false|false|false|||Treatment
Finding|Conceptual Entity|Discharge Instructions|5759,5768|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|Treatment
Finding|Functional Concept|Discharge Instructions|5759,5768|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|Treatment
Procedure|Health Care Activity|Discharge Instructions|5759,5768|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|Treatment
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|5759,5768|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|Treatment
Finding|Intellectual Product|Discharge Instructions|5769,5778|false|false|false|C3898838;C4321352|Frequency;How Often|Frequency
Drug|Hazardous or Poisonous Substance|Discharge Instructions|5780,5787|false|false|false|C0728873|Monitor brand of insecticide|monitor
Drug|Organic Chemical|Discharge Instructions|5780,5787|false|false|false|C0728873|Monitor brand of insecticide|monitor
Anatomy|Body System|Discharge Instructions|5788,5792|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|Discharge Instructions|5788,5792|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|Discharge Instructions|5788,5792|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Event|Event|Discharge Instructions|5788,5792|false|false|false|||skin
Finding|Body Substance|Discharge Instructions|5788,5792|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|Discharge Instructions|5788,5792|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Anatomy|Body Location or Region|Discharge Instructions|5796,5800|false|false|false|C0008114|Chin|chin
Procedure|Health Care Activity|Discharge Instructions|5796,5800|false|false|false|C2226982|examination of chin|chin
Anatomy|Body Location or Region|Discharge Instructions|5805,5817|false|false|false|C0230005|Occipital region|back of head
Anatomy|Body Location or Region|Discharge Instructions|5813,5817|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|5813,5817|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|Discharge Instructions|5813,5817|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|5813,5817|false|false|false|C0876917|Procedure on head|head
Disorder|Acquired Abnormality|Discharge Instructions|5822,5831|false|false|false|C1265875|Disintegration (morphologic abnormality)|breakdown
Event|Event|Discharge Instructions|5822,5831|false|false|false|||breakdown
Finding|Organism Function|Discharge Instructions|5822,5831|false|false|false|C0699900|Catabolism|breakdown
Event|Event|Discharge Instructions|5837,5843|false|false|false|||collar
Procedure|Health Care Activity|Discharge Instructions|5846,5854|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|5855,5867|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|5855,5867|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|5855,5867|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

