CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Known|Modifier|false|false||Knownnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Adverse reaction to drug|Finding|true|false||Adverse Drug Reactionsnull|Adverse reaction to drug|Finding|true|false||Drug Reactionsnull|Pharmaceutical Preparations|Drug|false|false||Drug
null|Pharmacologic Substance|Drug|false|false||Drugnull|Drug problem|Finding|false|false||Drugnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Chief complaint (finding)|Finding|false|false||Chief Complaintnull|Complaint (finding)|Finding|false|false||Complaintnull|null|Attribute|false|false||Complaintnull|Patient Outcome - Worsening|Finding|false|false||Worseningnull|Worsening (qualifier value)|Modifier|false|false||Worseningnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false||ABDnull|ABD (body structure)|Anatomy|false|false||ABD
null|Abdomen|Anatomy|false|false||ABDnull|Pathological Dilatation|Finding|false|false||distension
null|Distention|Finding|false|false||distensionnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Paracentesis|Procedure|false|false||Paracentesisnull|History of present illness (finding)|Finding|false|false||History of Present Illnessnull|null|Attribute|false|false||History of Present Illnessnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Present illness|Finding|false|false||Present Illnessnull|Present|Finding|false|false||Present
null|Presentation|Finding|false|false||Presentnull|Illness (finding)|Finding|false|false||Illnessnull|hepatitis C virus|Disorder|false|false||HCV
null|Hepatitis C|Disorder|false|false||HCVnull|Liver Cirrhosis|Disorder|false|false||cirrhosis
null|Cirrhosis|Disorder|false|false||cirrhosisnull|Ascites|Disorder|false|false||ascitesnull|Peritoneal Effusion|Finding|false|false||ascitesnull|HIV Vaccine|Drug|false|false||hiv
null|HIV Vaccine|Drug|false|false||hivnull|HIV Infections|Disorder|false|false||hiv
null|HIV|Disorder|false|false||hivnull|artesunate|Drug|false|false||ART
null|artesunate|Drug|false|false||ARTnull|AGRP wt Allele|Finding|false|false||ART
null|AGRP gene|Finding|false|false||ARTnull|Assisted Reproductive Technologies|Procedure|false|false||ART
null|Antiretroviral therapy|Procedure|false|false||ARTnull|Artwork|Device|false|false||ARTnull|Arts|Subject|false|false||ARTnull|intravenous drug use|Finding|false|false||IVDUnull|Intravenous drug user|Subject|false|false||IVDUnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|6-pyruvoyl-tetrahydropterin synthase deficiency|Disorder|false|false||PTSD
null|Post-Traumatic Stress Disorder|Disorder|false|false||PTSDnull|Patient Outcome - Worsening|Finding|false|false||worseningnull|Worsening (qualifier value)|Modifier|false|false||worseningnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false||abdnull|ABD (body structure)|Anatomy|false|false||abd
null|Abdomen|Anatomy|false|false||abdnull|Pathological Dilatation|Finding|false|false||distension
null|Distention|Finding|false|false||distensionnull|Past Week|Time|false|false||past weeknull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|subscriber - self|Finding|false|false||self
null|Self|Finding|false|false||selfnull|Lasix|Drug|false|false||lasix
null|Lasix|Drug|false|false||lasixnull|week|Time|false|false||weeksnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|More|LabModifier|false|false||morenull|Chemicals|Drug|false|false||chemicalsnull|Document Confidentiality Status - Restricted|Finding|false|false||restricted
null|Confidentiality - restricted|Finding|false|false||restricted
null|Confidentiality code - Restricted|Finding|false|false||restricted
null|Restricted|Finding|false|false||restrictednull|Diet|Drug|false|false||dietsnull|Past Week|Time|false|false||past weeknull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Patient Outcome - Worsening|Finding|false|false||worseningnull|Worsening (qualifier value)|Modifier|false|false||worseningnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false||abdnull|ABD (body structure)|Anatomy|false|false||abd
null|Abdomen|Anatomy|false|false||abdnull|Pathological Dilatation|Finding|false|false||distension
null|Distention|Finding|false|false||distensionnull|Discomfort|Finding|false|false||discomfortnull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Dyspnea|Finding|false|false||SOBnull|sleeping upright or using specific number of extra pillows (orthopnea)|Finding|false|false||orthopnea
null|Orthopnea|Finding|false|false||orthopneanull|Dysuria|Finding|false|false||dysurianull|Food Poisoning|Disorder|false|false||food poisoningnull|Food allergenic extracts|Drug|false|false||food
null|Food|Drug|false|false||food
null|Food allergenic extracts|Drug|false|false||foodnull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|Lopes Gorlin syndrome|Disorder|false|false||stalenull|Topical Cake|Drug|false|false||cake
null|Cake|Drug|false|false||cakenull|Minangkabau Language|Entity|false|false||minnull|Minute of time|Time|false|false||minnull|Minimum|Modifier|false|false||minnull|Minute Unit of Plane Angle|LabModifier|false|false||min
null|minim|LabModifier|false|false||minnull|Postprandial Period|Time|false|false||after foodnull|Food allergenic extracts|Drug|false|false||food
null|Food|Drug|false|false||food
null|Food allergenic extracts|Drug|false|false||foodnull|Ingestion|Phenomenon|false|false||ingestionnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Recent|Time|false|false||recentnull|Illness (finding)|Finding|false|false||illnessnull|Illness (finding)|Finding|false|false||sicknull|Contacts|Procedure|false|false||contactsnull|Gingival Hemorrhage|Finding|false|false||gum bleedingnull|Gum as an ingredient|Drug|false|false||gum
null|Gum Dose Form|Drug|false|false||gumnull|OTULIN wt Allele|Finding|false|false||gum
null|OTULIN gene|Finding|false|false||gumnull|Gingiva|Anatomy|false|false||gumnull|Gum - unit of product usage|LabModifier|false|false||gum
null|Gum Dosing Unit|LabModifier|false|false||gumnull|Hemorrhage|Finding|false|false||bleedingnull|examination of teeth|Procedure|false|false||teethnull|Head>Teeth|Anatomy|false|false||teeth
null|Tooth structure|Anatomy|false|false||teethnull|Recent|Time|false|false||recentnull|week|Time|false|false||weeksnull|Increased tendency to bruise|Finding|true|false||easy bruisingnull|Easy|Finding|false|false||easynull|Contusions|Disorder|true|false||bruisingnull|reported bruising (history)|Finding|true|false||bruisingnull|Melena|Finding|true|false||melenanull|Hematochezia|Disorder|true|false||BRBPRnull|Hemoptysis|Finding|false|false||hemoptysisnull|Hematuria|Disorder|false|false||hematurianull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false||abdnull|ABD (body structure)|Anatomy|false|false||abd
null|Abdomen|Anatomy|false|false||abdnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Further|Modifier|false|false||furthernull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Report (document)|Finding|false|false||reportnull|Reporting|Procedure|false|false||reportnull|null|Attribute|false|false||reportnull|Behavior Rating Inventory of Executive Function|Finding|false|false||brief
null|BRIEF Health Literacy Screening Tool|Finding|false|false||briefnull|Brief|Time|false|false||briefnull|Shortened|Modifier|false|false||briefnull|Menstruation|Finding|false|false||periodnull|Clinical Trial Period|Procedure|false|false||periodnull|per period (qualifier value)|Time|false|false||period
null|Time periods|Time|false|false||periodnull|Transaction counts and value totals - Period|LabModifier|false|false||periodnull|Confusion|Disorder|false|false||confusionnull|Clouded consciousness|Finding|false|false||confusionnull|Ultrasonic|Finding|true|false||ultrasoundnull|Urological ultrasound|Procedure|true|false||ultrasound
null|Ultrasonography|Procedure|true|false||ultrasoundnull|ultrasound device|Device|true|false||ultrasoundnull|Ultrasonic Shockwave|Phenomenon|true|false||ultrasound
null|Ultrasonics (sound)|Phenomenon|true|false||ultrasoundnull|Recent|Time|false|false||recentnull|Drug usage|Disorder|true|false||drug usenull|Encounter due to drug use|Finding|true|false||drug use
null|Drug use history|Finding|true|false||drug usenull|Pharmaceutical Preparations|Drug|true|false||drug
null|Pharmacologic Substance|Drug|true|false||drugnull|Drug problem|Finding|true|false||drugnull|Use - dosing instruction imperative|Finding|false|false||use
null|utilization qualifier|Finding|false|false||use
null|Usage|Finding|false|false||usenull|Alcohols|Drug|false|false||alcohol
null|Alcohols|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcoholnull|Alcohol - Recreational Drug Use Code|Finding|false|false||alcoholnull|Confusion|Disorder|false|false||confusednull|Precaution Code - Confused|Finding|false|false||confused
null|Clouded consciousness|Finding|false|false||confusednull|Forgetful|Finding|false|false||forgetfulnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Initial (abbreviation)|Finding|false|false||initialnull|Initially|Time|false|false||initialnull|Firstly|Modifier|false|false||initialnull|Laboratory test finding|Lab|false|false||Labsnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||ASTnull|Atypical Spitz Nevus|Disorder|false|false||ASTnull|SLC17A5 wt Allele|Finding|false|false||AST
null|SLC17A5 gene|Finding|false|false||AST
null|GOT1 gene|Finding|false|false||ASTnull|Asterion|Anatomy|false|false||ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Leukocytes|Anatomy|false|false||WBCnull|Blood Platelets|Anatomy|false|false||plateletnull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|hepatitis C virus|Disorder|false|false||HCV
null|Hepatitis C|Disorder|false|false||HCVnull|Liver Cirrhosis|Disorder|false|false||Cirrhosis
null|Cirrhosis|Disorder|false|false||Cirrhosisnull|Medical History|Finding|true|false||history ofnull|History of present illness (finding)|Finding|true|false||history
null|History of previous events|Finding|true|false||history
null|Historical aspects qualifier|Finding|true|false||history
null|Medical History|Finding|true|false||history
null|Concept History|Finding|true|false||historynull|History|Subject|false|false||historynull|Abnormal cervical smear|Finding|true|false||abnormal Pap smearsnull|Observation Interpretation - Abnormal|Finding|true|false||abnormal
null|Abnormal|Finding|true|false||abnormalnull|Pap smear|Procedure|true|false||Pap smearsnull|alpha 2-plasmin inhibitor-plasmin complex|Drug|true|false||Pap
null|alpha 2-plasmin inhibitor-plasmin complex|Drug|true|false||Pap
null|ACPP protein, human|Drug|true|false||Pap
null|ACPP protein, human|Drug|true|false||Papnull|null|Finding|true|false||Pap
null|PAPOLA wt Allele|Finding|true|false||Pap
null|PDAP1 gene|Finding|true|false||Pap
null|TUSC2 wt Allele|Finding|true|false||Pap
null|ASAP1 wt Allele|Finding|true|false||Pap
null|ACP3 wt Allele|Finding|true|false||Pap
null|Pulmonary artery pressure|Finding|true|false||Pap
null|TUSC2 gene|Finding|true|false||Pap
null|ASAP2 gene|Finding|true|false||Pap
null|ASAP1 gene|Finding|true|false||Pap
null|REG3A gene|Finding|true|false||Pap
null|PITUITARY ADENOMA PREDISPOSITION|Finding|true|false||Pap
null|PAPOLA gene|Finding|true|false||Pap
null|ACP3 gene|Finding|true|false||Pap
null|REG3A wt Allele|Finding|true|false||Pap
null|MRPS30 gene|Finding|true|false||Papnull|pars anterior of the paramedian lobule|Anatomy|false|false||Papnull|Papiamento language|Entity|true|false||Papnull|Smear test|Procedure|true|false||smearsnull|Physiologic calcification|Finding|false|false||calcification
null|Calcification|Finding|false|false||calcification
null|Calcinosis|Finding|false|false||calcificationnull|Calcified (qualifier value)|Modifier|false|false||calcificationnull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||breastnull|Breast problem|Finding|false|false||breastnull|Procedures on breast|Procedure|false|false||breastnull|Breast|Anatomy|false|false||breastnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Benign|Modifier|false|false||benignnull|HIV Infections|Disorder|false|false||HIV diseasenull|HIV Vaccine|Drug|false|false||HIV
null|HIV Vaccine|Drug|false|false||HIVnull|HIV Infections|Disorder|false|false||HIV
null|HIV|Disorder|false|false||HIVnull|Disease|Disorder|false|false||diseasenull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Past history of|Finding|false|false||Past history ofnull|Past history of|Finding|false|false||Past historynull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Location characteristic ID - Smoking|Finding|false|false||smoking
null|Smoking|Finding|false|false||smoking
null|Tobacco smoking behavior|Finding|false|false||smokingnull|Skin lesion|Disorder|false|false||skin lesionnull|Skin and subcutaneous tissue disorders|Disorder|false|false||skin
null|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||skinnull|Skin Specimen Source Code|Finding|false|false||skin
null|Skin Specimen|Finding|false|false||skinnull|Skin, Human|Anatomy|false|false||skin
null|Skin|Anatomy|false|false||skinnull|Lesion|Finding|false|false||lesion
null|null|Finding|false|false||lesionnull|Malignant neoplasm of skin|Disorder|false|false||skin cancernull|Skin and subcutaneous tissue disorders|Disorder|false|false||skin
null|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||skinnull|Skin Specimen Source Code|Finding|false|false||skin
null|Skin Specimen|Finding|false|false||skinnull|Skin, Human|Anatomy|false|false||skin
null|Skin|Anatomy|false|false||skinnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Patient-Reported|Finding|false|false||patient reportnull|Report source - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Relationship modifier - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Report (document)|Finding|false|false||reportnull|Reporting|Procedure|false|false||reportnull|null|Attribute|false|false||reportnull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|removal technique|Procedure|false|false||removal
null|Excision|Procedure|false|false||removal
null|Extraction|Procedure|false|false||removalnull|Removing (action)|Event|false|false||removalnull|Skin lesion|Disorder|false|false||skin lesionnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false||skinnull|Skin Specimen Source Code|Finding|false|false||skin
null|Skin Specimen|Finding|false|false||skinnull|Skin, Human|Anatomy|false|false||skin
null|Skin|Anatomy|false|false||skinnull|Lesion|Finding|false|false||lesion
null|null|Finding|false|false||lesionnull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Lesion|Finding|false|false||lesion
null|null|Finding|false|false||lesionnull|Forehead|Anatomy|false|false||foreheadnull|Purple|Modifier|false|false||purplenull|Abnormal color|Finding|false|false||discolorationnull|Sarcoma|Disorder|false|false||sarcoma
null|Malignant neoplasm of soft tissue|Disorder|false|false||sarcomanull|Pending - Allergy Clinical Status|Finding|false|false||pending
null|Pending - referral status|Finding|false|false||pendingnull|Pending - status|Time|false|false||pendingnull|pending - ManagedParticipationStatus|Modifier|false|false||pending
null|pending - RoleStatus|Modifier|false|false||pending
null|Pending - Day type|Modifier|false|false||pendingnull|Hypoechoic|Finding|false|false||hypoechoicnull|Lesion|Finding|false|false||lesion
null|null|Finding|false|false||lesionnull|Ultrasonic|Finding|false|false||ultrasoundnull|Urological ultrasound|Procedure|false|false||ultrasound
null|Ultrasonography|Procedure|false|false||ultrasoundnull|ultrasound device|Device|false|false||ultrasoundnull|Ultrasonic Shockwave|Phenomenon|false|false||ultrasound
null|Ultrasonics (sound)|Phenomenon|false|false||ultrasoundnull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Dysplasia of anus|Disorder|false|false||dysplasia of anusnull|Dysplasia|Disorder|false|false||dysplasianull|Anus Diseases|Disorder|false|false||anusnull|Procedure on anus|Procedure|false|false||anusnull|Anus|Anatomy|false|false||anusnull|Bipolar affective disorder, currently manic, mild|Disorder|false|false||Bipolar affective disorder, currently manic, mildnull|MAJOR AFFECTIVE DISORDER 4|Disorder|false|false||Bipolar affective disorder
null|MAJOR AFFECTIVE DISORDER 9|Disorder|false|false||Bipolar affective disorder
null|Bipolar Disorder|Disorder|false|false||Bipolar affective disorder
null|MAJOR AFFECTIVE DISORDER 2|Disorder|false|false||Bipolar affective disorder
null|MAJOR AFFECTIVE DISORDER 1|Disorder|false|false||Bipolar affective disorder
null|MAJOR AFFECTIVE DISORDER 8|Disorder|false|false||Bipolar affective disorder
null|MAJOR AFFECTIVE DISORDER 6|Disorder|false|false||Bipolar affective disorder
null|MAJOR AFFECTIVE DISORDER 7|Disorder|false|false||Bipolar affective disordernull|Bipolar|Modifier|false|false||Bipolarnull|Mood Disorders|Disorder|false|false||affective disordernull|Disease|Disorder|false|false||disordernull|Current (present time)|Time|false|false||currentlynull|Manic|Disorder|false|false||manicnull|Manic mood|Finding|false|false||manicnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Post-Traumatic Stress Disorder|Disorder|false|false||PTSD
null|6-pyruvoyl-tetrahydropterin synthase deficiency|Disorder|false|false||PTSDnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|cocaine|Drug|true|false||cocaine
null|cocaine|Drug|true|false||cocaine
null|cocaine|Drug|true|false||cocaine
null|cocaine|Drug|true|false||cocainenull|Poisoning by cocaine|Disorder|true|false||cocainenull|Cocaine measurement|Procedure|true|false||cocainenull|heroin|Drug|true|false||heroin
null|heroin|Drug|true|false||heroin
null|heroin|Drug|true|false||heroinnull|Poisoning by heroin|Disorder|true|false||heroinnull|Use - dosing instruction imperative|Finding|false|false||use
null|utilization qualifier|Finding|false|false||use
null|Usage|Finding|false|false||usenull|Social and personal history|Finding|false|false||Social History
null|Social History|Finding|false|false||Social Historynull|Social|Finding|false|false||Socialnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Family Medical History|Finding|false|false||Family Historynull|Entity Name Part Type - family|Finding|false|false||Family
null|Last Name|Finding|false|false||Family
null|Living Arrangement - Family|Finding|false|false||Family
null|Family (taxonomic)|Finding|false|false||Family
null|Family Collection|Finding|false|false||Familynull|Family|Subject|false|false||Familynull|History of present illness (finding)|Finding|false|true||History
null|History of previous events|Finding|false|true||History
null|Historical aspects qualifier|Finding|false|true||History
null|Medical History|Finding|false|true||History
null|Concept History|Finding|false|true||Historynull|History|Subject|false|false||Historynull|Total|Modifier|false|false||totalnull|Sibling|Subject|false|false||siblingsnull|Brother - courtesy title|Finding|false|false||brother
null|Relationship - Brother|Finding|false|false||brothernull|Brothers|Subject|false|false||brothernull|Touch Perception|Finding|false|false||touch
null|Touch sensation|Finding|false|false||touchnull|Therapeutic Touch|Procedure|false|false||touchnull|Tactile|Modifier|false|false||touchnull|Awareness|Finding|true|false||awarenull|Known|Modifier|false|false||knownnull|Liver diseases|Disorder|false|false||liver disease
null|Hepatobiliary Disorder|Disorder|false|false||liver diseasenull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Disease|Disorder|false|false||diseasenull|ErbB Receptors|Drug|false|false||her family
null|ErbB Receptors|Drug|false|false||her familynull|ErbB Receptors|Finding|false|false||her familynull|Entity Name Part Type - family|Finding|false|false||family
null|Last Name|Finding|false|false||family
null|Living Arrangement - Family|Finding|false|false||family
null|Family (taxonomic)|Finding|false|false||family
null|Family Collection|Finding|false|false||familynull|Family|Subject|false|false||familynull|Last|Modifier|false|false||lastnull|alcohol consumption (history)|Finding|false|false||alcohol consumption
null|Alcohol consumption|Finding|false|false||alcohol consumptionnull|Alcohols|Drug|false|false||alcohol
null|Alcohols|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcoholnull|Alcohol - Recreational Drug Use Code|Finding|false|false||alcoholnull|Consumption-archaic term for TB|Disorder|false|false||consumptionnull|biologic consumption|Finding|false|false||consumptionnull|Consumption of goods|Event|false|false||consumptionnull|Drink (dietary substance)|Drug|false|false||drinknull|month|Time|false|false||monthsnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|Regular|Modifier|false|false||regularnull|alcohol consumption (history)|Finding|false|false||alcohol consumption
null|Alcohol consumption|Finding|false|false||alcohol consumptionnull|Alcohols|Drug|false|false||alcohol
null|Alcohols|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcoholnull|Alcohol - Recreational Drug Use Code|Finding|false|false||alcoholnull|Consumption-archaic term for TB|Disorder|false|false||consumptionnull|biologic consumption|Finding|false|false||consumptionnull|Consumption of goods|Event|false|false||consumptionnull|Last|Modifier|false|false||Lastnull|Drug usage|Disorder|false|false||drug usenull|Encounter due to drug use|Finding|false|false||drug use
null|Drug use history|Finding|false|false||drug usenull|Pharmaceutical Preparations|Drug|false|false||drug
null|Pharmacologic Substance|Drug|false|false||drugnull|Drug problem|Finding|false|false||drugnull|Use - dosing instruction imperative|Finding|false|false||use
null|utilization qualifier|Finding|false|false||use
null|Usage|Finding|false|false||usenull|year|Time|false|false||yearsnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|Couple (action)|Finding|false|false||couplenull|Couples (persons)|Subject|false|false||couplenull|year|Time|false|false||yearsnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Generalnull|General medical service|Procedure|false|false||Generalnull|Generalized|Modifier|false|false||Generalnull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|HEENT|Anatomy|false|false||HEENTnull|cetrimonium bromide|Drug|false|false||CTABnull|Anicteric|Finding|false|false||anictericnull|Scleral Diseases|Disorder|false|false||scleranull|examination of sclera|Procedure|false|false||scleranull|Sclera|Anatomy|false|false||scleranull|Remote control command - Clear|Finding|false|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Passive joint movement of neck (finding)|Finding|false|false||Neck
null|Neck problem|Finding|false|false||Necknull|dendritic spine neck|Anatomy|false|false||Neck
null|Neck|Anatomy|false|false||Necknull|Supple|Finding|false|false||supplenull|Leukocyte adhesion deficiency type 1|Disorder|true|false||LAD
null|Leukocyte adhesion deficiency|Disorder|true|false||LADnull|ITGB2 wt Allele|Finding|true|false||LAD
null|DLD gene|Finding|true|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false||LADnull|Ladino Language|Entity|true|false||LADnull|Lung|Anatomy|false|false||Lungsnull|cetrimonium bromide|Drug|false|false||CTAbnull|Prolonged|Time|false|false||prolongednull|Expiration, Respiratory|Finding|false|false||expiratorynull|Phase|Time|false|false||phasenull|Malignant neoplasm of abdomen|Disorder|false|false||Abdomennull|Abdomen problem|Finding|false|false||Abdomennull|Abdomen|Anatomy|false|false||Abdomen
null|Abdominal Cavity|Anatomy|false|false||Abdomennull|Dilated|Finding|false|false||distendednull|Distended|Modifier|false|false||distendednull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Diffuse|Modifier|false|false||diffusenull|Emotional tenderness|Finding|false|false||tenderness
null|Sore to touch|Finding|false|false||tendernessnull|Flank (surface region)|Anatomy|false|false||flanknull|Dullness|Finding|false|false||dullnessnull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Malignant neoplasm of spleen|Disorder|false|false||spleennull|Spleen problem|Finding|false|false||spleennull|Procedures on Spleen|Procedure|false|false||spleennull|Abdomen>Spleen|Anatomy|false|false||spleen
null|Spleen|Anatomy|false|false||spleennull|Graph Edge|Finding|false|false||edgenull|Along edge (qualifier value)|Modifier|false|false||edgenull|Pathological Dilatation|Finding|false|false||distension
null|Distention|Finding|false|false||distensionnull|Hereditary Multiple Exostoses|Disorder|false|false||Extnull|EXT1 wt Allele|Finding|false|false||Ext
null|EXT1 gene|Finding|false|false||Extnull|Clubbing|Disorder|false|false||clubbingnull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|abscisic aldehyde oxidase activity|Finding|false|false||AAO3null|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|Mental Recall|Finding|false|false||recallnull|Recall (activity)|Event|false|false||recallnull|3 times|Finding|false|false||3 timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Minute of time|Time|false|false||minutesnull|Minute Unit of Plane Angle|LabModifier|false|false||minutes
null|Minute (diminutive)|LabModifier|false|false||minutes
null|Small|LabModifier|false|false||minutesnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|physical examination (physical finding)|Finding|false|false||PHYSICAL EXAMINATIONnull|Physical Examination|Procedure|false|false||PHYSICAL EXAMINATIONnull|physical examination (physical finding)|Finding|false|false||PHYSICAL
null|Physical|Finding|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||EXAMINATION
null|Medical Examination|Procedure|false|false||EXAMINATIONnull|Examination|Event|false|false||EXAMINATIONnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Generalnull|General medical service|Procedure|false|false||Generalnull|Generalized|Modifier|false|false||Generalnull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|HEENT|Anatomy|false|false||HEENTnull|Anicteric|Finding|false|false||anictericnull|Scleral Diseases|Disorder|false|false||scleranull|examination of sclera|Procedure|false|false||scleranull|Sclera|Anatomy|false|false||scleranull|Remote control command - Clear|Finding|false|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Passive joint movement of neck (finding)|Finding|false|false||Neck
null|Neck problem|Finding|false|false||Necknull|dendritic spine neck|Anatomy|false|false||Neck
null|Neck|Anatomy|false|false||Necknull|Supple|Finding|false|false||supplenull|Leukocyte adhesion deficiency type 1|Disorder|true|false||LAD
null|Leukocyte adhesion deficiency|Disorder|true|false||LADnull|ITGB2 wt Allele|Finding|true|false||LAD
null|DLD gene|Finding|true|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false||LADnull|Ladino Language|Entity|true|false||LADnull|Lung|Anatomy|false|false||Lungsnull|cetrimonium bromide|Drug|false|false||CTAbnull|Prolonged|Time|false|false||prolongednull|Expiration, Respiratory|Finding|false|false||expiratorynull|Phase|Time|false|false||phasenull|Malignant neoplasm of abdomen|Disorder|false|false||Abdomennull|Abdomen problem|Finding|false|false||Abdomennull|Abdomen|Anatomy|false|false||Abdomen
null|Abdominal Cavity|Anatomy|false|false||Abdomennull|Dilated|Finding|false|false||distendednull|Distended|Modifier|false|false||distendednull|Admission Level of Care Code - Improved|Finding|false|false||improved
null|Improved - answer to question|Finding|false|false||improved
null|Improved|Finding|false|false||improvednull|Better|Modifier|false|false||improvednull|thiamine triphosphorate|Drug|false|false||TTP
null|ZFP36 protein, human|Drug|false|false||TTP
null|ZFP36 protein, human|Drug|false|false||TTP
null|thiamine triphosphorate|Drug|false|false||TTPnull|Congenital Thrombotic Thrombocytopenic Purpura|Disorder|false|false||TTP
null|Purpura, Thrombotic Thrombocytopenic|Disorder|false|false||TTPnull|ZFP36 wt Allele|Finding|false|false||TTP
null|ZFP36 gene|Finding|false|false||TTP
null|ADAMTS13 gene|Finding|false|false||TTPnull|Time to Progression|Time|false|false||TTPnull|Structure of right upper quadrant of abdomen|Anatomy|false|false||RUQnull|RUQ - Right upper quadrant|Modifier|false|false||RUQnull|Hereditary Multiple Exostoses|Disorder|false|false||Extnull|EXT1 wt Allele|Finding|false|false||Ext
null|EXT1 gene|Finding|false|false||Extnull|Clubbing|Disorder|false|false||clubbingnull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|abscisic aldehyde oxidase activity|Finding|false|false||AAO3null|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Mandibular right central incisor mesial prosthesis|Device|false|false||25PMnull|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSEnull|Glucose measurement|Procedure|false|false||GLUCOSEnull|Glucose^1.5H post dose glucagon|Lab|false|false||GLUCOSEnull|urea|Drug|false|false||UREA
null|urea|Drug|false|false||UREA
null|urea|Drug|false|false||UREAnull|Urea measurement|Procedure|false|false||UREAnull|Sodium supplements|Drug|false|false||SODIUM
null|sodium|Drug|false|false||SODIUM
null|sodium|Drug|false|false||SODIUM
null|Sodium Drug Class|Drug|false|false||SODIUMnull|Sodium metabolic function|Finding|false|false||SODIUMnull|Sodium measurement|Procedure|false|false||SODIUMnull|Potassium Drug Class|Drug|false|false||POTASSIUM
null|Dietary Potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|Potassium supplement|Drug|false|false||POTASSIUM
null|Potassium supplement|Drug|false|false||POTASSIUMnull|Potassium metabolic function|Finding|false|false||POTASSIUMnull|Potassium measurement|Procedure|false|false||POTASSIUMnull|chloride ion|Drug|false|false||CHLORIDE
null|Chlorides|Drug|false|false||CHLORIDEnull|Chloride metabolic function|Finding|false|false||CHLORIDEnull|Chloride measurement|Procedure|false|false||CHLORIDEnull|Total|Modifier|false|false||TOTALnull|carbon dioxide|Drug|false|false||CO2
null|carbon dioxide|Drug|false|false||CO2null|MT-CO2 gene|Finding|false|false||CO2
null|null|Finding|false|false||CO2
null|C2 wt Allele|Finding|false|false||CO2null|blood anion gap (lab test)|Procedure|false|false||ANION GAP
null|Anion gap measurement|Procedure|false|false||ANION GAPnull|Anion Gap|Attribute|false|false||ANION GAPnull|Anion gap result|Lab|false|false||ANION GAPnull|Anions|Drug|false|false||ANIONnull|Ras GTPase-Activating Protein 1, Human|Drug|false|false||GAP
null|Ras GTPase-Activating Protein 1, Human|Drug|false|false||GAP
null|GTPase-Activating Proteins|Drug|false|false||GAP
null|GTPase-Activating Proteins|Drug|false|false||GAPnull|RASA1 wt Allele|Finding|false|false||GAP
null|RASA1 gene|Finding|false|false||GAPnull|Gap (space)|Modifier|false|false||GAPnull|Mandibular right central incisor mesial prosthesis|Device|false|false||25PMnull|Mandibular right central incisor mesial prosthesis|Device|false|false||25PMnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGPT - Glutamate pyruvate transaminase|Drug|false|false||SGPT
null|SGPT - Glutamate pyruvate transaminase|Drug|false|false||SGPTnull|GPT gene|Finding|false|false||SGPTnull|Serum Alanine Transaminase Test|Procedure|false|false||SGPTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||ASTnull|Atypical Spitz Nevus|Disorder|false|false||ASTnull|SLC17A5 wt Allele|Finding|false|false||AST
null|SLC17A5 gene|Finding|false|false||AST
null|GOT1 gene|Finding|false|false||ASTnull|Asterion|Anatomy|false|false||ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||SGOT
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||SGOTnull|GOT1 gene|Finding|false|false||SGOTnull|Aspartate aminotransferase measurement|Procedure|false|false||SGOTnull|Alkaline Phosphatase|Drug|false|false||ALK PHOS
null|Alkaline Phosphatase|Drug|false|false||ALK PHOSnull|Alkaline phosphatase measurement|Procedure|false|false||ALK PHOSnull|ALK protein, human|Drug|false|false||ALK
null|ALK protein, human|Drug|false|false||ALKnull|ALK protein, human|Finding|false|false||ALK
null|ALK gene|Finding|false|false||ALK
null|ALK wt Allele|Finding|false|false||ALKnull|Phos <Photinae>|Entity|false|false||PHOSnull|Mandibular right central incisor mesial prosthesis|Device|false|false||25PMnull|lipase|Drug|false|false||LIPASE
null|lipase|Drug|false|false||LIPASE
null|lipase|Drug|false|false||LIPASEnull|Lipase measurement|Procedure|false|false||LIPASEnull|Mandibular right central incisor mesial prosthesis|Device|false|false||25PMnull|Albumin|Drug|false|false||ALBUMIN
null|Albumins|Drug|false|false||ALBUMIN
null|Albumins|Drug|false|false||ALBUMIN
null|Albumin|Drug|false|false||ALBUMINnull|Albumin metabolic function|Finding|false|false||ALBUMIN
null|ALB gene|Finding|false|false||ALBUMINnull|Albumin measurement|Procedure|false|false||ALBUMINnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||HGB
null|Hemoglobin|Drug|false|false||HGBnull|CYGB gene|Finding|false|false||HGBnull|Hemoglobin concentration|Lab|false|false||HGBnull|Hemopoietic stem cell transplant|Procedure|false|false||HCT
null|Hematocrit Measurement|Procedure|false|false||HCTnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Lymph|Finding|false|false||LYMPHSnull|Monos|Drug|false|false||MONOS
null|Mono-S|Drug|false|false||MONOS
null|Monos|Drug|false|false||MONOSnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||EOS
null|Familial eosinophilia|Disorder|false|false||EOSnull|PRSS33 gene|Finding|false|false||EOS
null|IKZF4 gene|Finding|false|false||EOSnull|Eos <Loriini>|Entity|false|false||EOSnull|Mandibular right central incisor mesial prosthesis|Device|false|false||25PMnull|Primed lymphocyte test|Procedure|false|false||PLTnull|Count Dosing Unit|LabModifier|false|false||COUNT
null|Count|LabModifier|false|false||COUNTnull|Mandibular right central incisor mesial prosthesis|Device|false|false||25PMnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Mandibular right central incisor mesial prosthesis|Device|false|false||25PMnull|Plain chest X-ray|Procedure|false|false||CXRnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Cardiovascular disease+Pulmonary disease|Disorder|false|false||cardiopulmonarynull|Cardiopulmonary|Anatomy|false|false||cardiopulmonarynull|Process Pharmacologic Substance|Drug|true|false||processnull|Process (qualifier value)|Finding|true|false||processnull|bony process|Anatomy|false|false||processnull|Process|Phenomenon|true|false||processnull|patient appearance regarding mental status exam|Procedure|false|false||appearancenull|null|Attribute|false|false||appearancenull|Personal appearance|Subject|false|false||appearancenull|Appearance|Modifier|false|false||appearancenull|Kind of quantity - Appearance|LabModifier|false|false||appearancenull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Consistent with|Finding|false|false||compatible withnull|Compatible|Modifier|false|false||compatible withnull|Consistent with|Finding|false|false||compatiblenull|Compatible|Modifier|false|false||compatiblenull|Liver Cirrhosis|Disorder|false|false||cirrhosis
null|Cirrhosis|Disorder|false|false||cirrhosisnull|Aspects of signs|Finding|false|false||Signs
null|Physical findings|Finding|false|false||Signsnull|Manufactured sign|Device|false|false||Signsnull|Hepatic|Anatomy|false|false||portalnull|Hypertensive disease|Disorder|false|false||hypertensionnull|Small amount|LabModifier|false|false||small amountnull|Small|LabModifier|false|false||smallnull|Amount class - Amount|Finding|false|false||amountnull|Quantity|LabModifier|false|false||amountnull|Ascites|Disorder|false|false||ascitesnull|Peritoneal Effusion|Finding|false|false||ascitesnull|Splenomegaly|Finding|false|false||splenomegalynull|Cholelithiasis|Disorder|false|false||Cholelithiasisnull|Legal patent|Finding|false|false||Patentnull|Open|Modifier|false|false||Patentnull|Portal vein structure|Anatomy|false|false||portal veinsnull|Hepatic|Anatomy|false|false||portalnull|Procedure on vein|Procedure|false|false||veinsnull|Veins|Anatomy|false|false||veinsnull|Flow|Phenomenon|false|false||flownull|Diagnostic agents|Drug|false|false||Diagnosticnull|Location Service Code - Diagnostic|Finding|false|false||Diagnostic
null|Diagnostic|Finding|false|false||Diagnosticnull|Diagnostic dental procedure|Procedure|false|false||Diagnostic
null|Diagnosis|Procedure|false|false||Diagnosticnull|Parity|Finding|false|false||paranull|Para (Brazil)|Entity|false|false||paranull|Unsuccessful|Modifier|false|false||unsuccessfulnull|Floor (anatomic)|Anatomy|false|false||floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false||abdnull|ABD (body structure)|Anatomy|false|false||abd
null|Abdomen|Anatomy|false|false||abdnull|Pathological Dilatation|Finding|false|false||distension
null|Distention|Finding|false|false||distensionnull|Discomfort|Finding|false|false||discomfortnull|BRIEF Health Literacy Screening Tool|Finding|false|false||Brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||Briefnull|Brief|Time|false|false||Briefnull|Shortened|Modifier|false|false||Briefnull|Hospital course|Finding|false|false||Hospital Coursenull|null|Attribute|false|false||Hospital Coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||Coursenull|hepatitis C virus|Disorder|false|false||HCV
null|Hepatitis C|Disorder|false|false||HCVnull|Liver Cirrhosis|Disorder|false|false||cirrhosis
null|Cirrhosis|Disorder|false|false||cirrhosisnull|Ascites|Disorder|false|false||ascitesnull|Peritoneal Effusion|Finding|false|false||ascitesnull|HIV Vaccine|Drug|false|false||hiv
null|HIV Vaccine|Drug|false|false||hivnull|HIV Infections|Disorder|false|false||hiv
null|HIV|Disorder|false|false||hivnull|artesunate|Drug|false|false||ART
null|artesunate|Drug|false|false||ARTnull|AGRP wt Allele|Finding|false|false||ART
null|AGRP gene|Finding|false|false||ARTnull|Assisted Reproductive Technologies|Procedure|false|false||ART
null|Antiretroviral therapy|Procedure|false|false||ARTnull|Artwork|Device|false|false||ARTnull|Arts|Subject|false|false||ARTnull|intravenous drug use|Finding|false|false||IVDUnull|Intravenous drug user|Subject|false|false||IVDUnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|6-pyruvoyl-tetrahydropterin synthase deficiency|Disorder|false|false||PTSD
null|Post-Traumatic Stress Disorder|Disorder|false|false||PTSDnull|Patient Outcome - Worsening|Finding|false|false||worseningnull|Worsening (qualifier value)|Modifier|false|false||worseningnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false||abdnull|ABD (body structure)|Anatomy|false|false||abd
null|Abdomen|Anatomy|false|false||abdnull|Pathological Dilatation|Finding|false|false||distension
null|Distention|Finding|false|false||distensionnull|Past Week|Time|false|false||past weeknull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Confusion|Disorder|false|false||confusionnull|Clouded consciousness|Finding|false|false||confusionnull|Ascites|Disorder|false|false||Ascitesnull|Peritoneal Effusion|Finding|false|false||Ascitesnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false||abdnull|ABD (body structure)|Anatomy|false|false||abd
null|Abdomen|Anatomy|false|false||abdnull|Pathological Dilatation|Finding|false|false||distension
null|Distention|Finding|false|false||distensionnull|Discomfort|Finding|false|false||discomfortnull|Last|Modifier|false|false||lastnull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Hepatic|Anatomy|false|false||portalnull|Hypertensive disease|Disorder|false|false||HTNnull|Liver diseases|Disorder|false|false||liver disease
null|Hepatobiliary Disorder|Disorder|false|false||liver diseasenull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Disease|Disorder|false|false||diseasenull|Ascitic Fluid|Finding|false|false||ascitic fluidnull|Ascitic|Modifier|false|false||asciticnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Availability of|Finding|false|false||availablenull|Night time|Time|false|false||nightnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Congestive heart failure|Disorder|false|false||heart failure
null|Heart failure|Disorder|false|false||heart failurenull|Malignant neoplasm of heart|Disorder|false|false||heart
null|benign neoplasm of heart|Disorder|false|false||heartnull|HEART PROBLEM|Finding|false|false||heartnull|Chest>Heart|Anatomy|false|false||heart
null|Heart|Anatomy|false|false||heartnull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Multiple Epiphyseal Dysplasia|Disorder|false|false||mednull|Master of Education|Finding|false|false||med
null|COMP wt Allele|Finding|false|false||med
null|COL9A3 gene|Finding|false|false||med
null|SCN8A wt Allele|Finding|false|false||med
null|COL9A2 gene|Finding|false|false||med
null|COMP gene|Finding|false|false||med
null|SCN8A gene|Finding|false|false||mednull|Lacking|Modifier|false|false||lacknull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Restricted|Finding|false|false||restrictionnull|Androgen Binding Protein|Drug|true|false||SBP
null|Androgen Binding Protein|Drug|true|false||SBPnull|CCHCR1 wt Allele|Finding|true|false||SBP
null|SHBG wt Allele|Finding|true|false||SBPnull|Systolic blood pressure measurement|Procedure|true|false||SBPnull|Systolic Pressure|Attribute|true|false||SBPnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Diuretics|Drug|false|false||diureticsnull|furosemide|Drug|false|false||Furosemide
null|furosemide|Drug|false|false||Furosemidenull|Daily|Time|false|false||DAILYnull|spironolactone|Drug|false|false||Spironolactone
null|spironolactone|Drug|false|false||Spironolactonenull|Daily|Time|false|false||DAILYnull|Usual|Modifier|false|false||usualnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Plain chest X-ray|Procedure|false|false||CXRnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Urine culture|Procedure|true|false||Urine culturenull|Portion of urine|Finding|false|false||Urine
null|null|Finding|false|false||Urine
null|Urine|Finding|false|false||Urine
null|In Urine|Finding|false|false||Urine
null|Urine specimen|Finding|false|false||Urinenull|Blood culture|Procedure|false|false||culture bloodnull|Culture Dose Form|Drug|false|false||culturenull|Culture (Anthropological)|Finding|false|false||culture
null|Cultural aspects|Finding|false|false||culturenull|Microbial culture (procedure)|Procedure|false|false||culture
null|Laboratory culture|Procedure|false|false||culturenull|Blood culture negative|Lab|false|false||blood culture negativenull|Blood culture|Procedure|false|false||blood culturenull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Culture negative|Lab|false|false||culture negativenull|Culture Dose Form|Drug|false|false||culturenull|Culture (Anthropological)|Finding|false|false||culture
null|Cultural aspects|Finding|false|false||culturenull|Microbial culture (procedure)|Procedure|false|false||culture
null|Laboratory culture|Procedure|false|false||culturenull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Hypervolemia (finding)|Finding|false|false||excess fluid
null|Edema|Finding|false|false||excess fluidnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Table Frame - above|Finding|false|false||abovenull|Upper|Modifier|false|false||abovenull|GDC Regimen Terminology|Finding|false|false||regimennull|Treatment Protocols|Procedure|false|false||regimennull|Electrical Current|Phenomenon|false|false||currentnull|Current (present time)|Time|false|false||currentnull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Liver brand of Vitamin B 12|Drug|false|false||Liver
null|liver extract|Drug|false|false||Liver
null|liver extract|Drug|false|false||Liver
null|Liver brand of Vitamin B 12|Drug|false|false||Liver
null|Liver brand of Vitamin B 12|Drug|false|false||Livernull|Benign neoplasm of liver|Disorder|false|false||Liver
null|Liver diseases|Disorder|false|false||Livernull|Liver problem|Finding|false|false||Livernull|Procedures on liver|Procedure|false|false||Livernull|Abdomen>Liver|Anatomy|false|false||Liver
null|null|Anatomy|false|false||Liver
null|Liver|Anatomy|false|false||Livernull|Clinic|Device|false|false||clinic
null|Ambulatory Care Facilities|Device|false|false||clinicnull|Clinic|Entity|false|false||clinic
null|Ambulatory Care Facilities|Entity|false|false||clinicnull|Patient location type - Clinic|Modifier|false|false||clinic
null|Person location type - Clinic|Modifier|false|false||clinicnull|Schedule (document)|Finding|false|false||schedulenull|Scheduling (procedure)|Procedure|false|false||schedulenull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Screening - procedure intent|Finding|false|false||screening
null|Special screening finding|Finding|false|false||screening
null|Aspects of disease screening|Finding|false|false||screeningnull|research subject screening|Procedure|false|false||screening
null|Disease Screening|Procedure|false|false||screening
null|Screening|Procedure|false|false||screening
null|Screening for cancer|Procedure|false|false||screening
null|Screening procedure|Procedure|false|false||screeningnull|Esophagogastroduodenoscopy|Procedure|false|false||EGDnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Accurate (qualifier value)|Modifier|false|false||accuratenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|furosemide|Drug|false|false||Furosemide
null|furosemide|Drug|false|false||Furosemidenull|Daily|Time|false|false||DAILYnull|spironolactone|Drug|false|false||Spironolactone
null|spironolactone|Drug|false|false||Spironolactonenull|Daily|Time|false|false||DAILYnull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|Inhaler (unit of presentation)|Finding|false|false||Inhalernull|Inhaler|Device|false|false||Inhalernull|Inhaler Dosing Unit|LabModifier|false|false||Inhalernull|Puff Dosing Unit|LabModifier|false|false||PUFF
null|Picofarad|LabModifier|false|false||PUFFnull|Every four hours|Time|false|false||Q4Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Wheezing|Finding|false|false||wheezingnull|Dyspnea|Finding|false|false||SOBnull|raltegravir|Drug|false|false||Raltegravir
null|raltegravir|Drug|false|false||Raltegravirnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Emtricitabine- and tenofovir-containing product|Drug|false|false||Emtricitabine-Tenofovir
null|Emtricitabine- and tenofovir-containing product|Drug|false|false||Emtricitabine-Tenofovirnull|emtricitabine|Drug|false|false||Emtricitabine
null|emtricitabine|Drug|false|false||Emtricitabinenull|tenofovir|Drug|false|false||Tenofovir
null|tenofovir|Drug|false|false||Tenofovirnull|Truvada|Drug|false|false||Truvada
null|Truvada|Drug|false|false||Truvadanull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|Daily|Time|false|false||DAILYnull|Nicotine Transdermal Patch|Drug|false|false||Nicotine Patchnull|nicotine|Drug|false|false||Nicotine
null|nicotine|Drug|false|false||Nicotinenull|Patch - Extended Release Film|Drug|false|false||Patch
null|Human patch material|Drug|false|false||Patch
null|Body tissue patch material|Drug|false|false||Patchnull|Plaque (lesion)|Finding|false|false||Patchnull|Patch Dosage Form|Device|false|false||Patch
null|Surgical patch|Device|false|false||Patchnull|Patch (unit of presentation)|LabModifier|false|false||Patch
null|Patch Dosing Unit|LabModifier|false|false||Patchnull|Daily|Time|false|false||DAILYnull|ipratropium bromide|Drug|false|false||Ipratropium Bromide
null|ipratropium bromide|Drug|false|false||Ipratropium Bromidenull|ipratropium|Drug|false|false||Ipratropium
null|ipratropium|Drug|false|false||Ipratropiumnull|Bromides|Drug|false|false||Bromidenull|Bromides measurement|Procedure|false|false||Bromidenull|NEB protein, human|Drug|false|false||Neb
null|NEB protein, human|Drug|false|false||Neb
null|Nebulizer solution|Drug|false|false||Nebnull|NEB gene|Finding|false|false||Neb
null|mitotic nuclear membrane disassembly|Finding|false|false||Nebnull|NEB protein, human|Drug|false|false||NEB
null|NEB protein, human|Drug|false|false||NEB
null|Nebulizer solution|Drug|false|false||NEBnull|NEB gene|Finding|false|false||NEB
null|mitotic nuclear membrane disassembly|Finding|false|false||NEBnull|Every six hours|Time|false|false||Q6Hnull|Dyspnea|Finding|false|false||SOBnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|Inhaler (unit of presentation)|Finding|false|false||Inhalernull|Inhaler|Device|false|false||Inhalernull|Inhaler Dosing Unit|LabModifier|false|false||Inhalernull|Puff Dosing Unit|LabModifier|false|false||PUFF
null|Picofarad|LabModifier|false|false||PUFFnull|Every four hours|Time|false|false||Q4Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Wheezing|Finding|false|false||wheezingnull|Dyspnea|Finding|false|false||SOBnull|Emtricitabine- and tenofovir-containing product|Drug|false|false||Emtricitabine-Tenofovir
null|Emtricitabine- and tenofovir-containing product|Drug|false|false||Emtricitabine-Tenofovirnull|emtricitabine|Drug|false|false||Emtricitabine
null|emtricitabine|Drug|false|false||Emtricitabinenull|tenofovir|Drug|false|false||Tenofovir
null|tenofovir|Drug|false|false||Tenofovirnull|Truvada|Drug|false|false||Truvada
null|Truvada|Drug|false|false||Truvadanull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|Daily|Time|false|false||DAILYnull|furosemide|Drug|false|false||Furosemide
null|furosemide|Drug|false|false||Furosemidenull|Daily|Time|false|false||DAILYnull|furosemide|Drug|false|false||furosemide
null|furosemide|Drug|false|false||furosemidenull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Daily|Time|false|false||Dailynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|ipratropium bromide|Drug|false|false||Ipratropium Bromide
null|ipratropium bromide|Drug|false|false||Ipratropium Bromidenull|ipratropium|Drug|false|false||Ipratropium
null|ipratropium|Drug|false|false||Ipratropiumnull|Bromides|Drug|false|false||Bromidenull|Bromides measurement|Procedure|false|false||Bromidenull|NEB protein, human|Drug|false|false||Neb
null|NEB protein, human|Drug|false|false||Neb
null|Nebulizer solution|Drug|false|false||Nebnull|NEB gene|Finding|false|false||Neb
null|mitotic nuclear membrane disassembly|Finding|false|false||Nebnull|NEB protein, human|Drug|false|false||NEB
null|NEB protein, human|Drug|false|false||NEB
null|Nebulizer solution|Drug|false|false||NEBnull|NEB gene|Finding|false|false||NEB
null|mitotic nuclear membrane disassembly|Finding|false|false||NEBnull|Every six hours|Time|false|false||Q6Hnull|Dyspnea|Finding|false|false||SOBnull|Nicotine Transdermal Patch|Drug|false|false||Nicotine Patchnull|nicotine|Drug|false|false||Nicotine
null|nicotine|Drug|false|false||Nicotinenull|Patch - Extended Release Film|Drug|false|false||Patch
null|Human patch material|Drug|false|false||Patch
null|Body tissue patch material|Drug|false|false||Patchnull|Plaque (lesion)|Finding|false|false||Patchnull|Patch Dosage Form|Device|false|false||Patch
null|Surgical patch|Device|false|false||Patchnull|Patch (unit of presentation)|LabModifier|false|false||Patch
null|Patch Dosing Unit|LabModifier|false|false||Patchnull|Daily|Time|false|false||DAILYnull|raltegravir|Drug|false|false||Raltegravir
null|raltegravir|Drug|false|false||Raltegravirnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|spironolactone|Drug|false|false||Spironolactone
null|spironolactone|Drug|false|false||Spironolactonenull|Daily|Time|false|false||DAILYnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Ascites|Disorder|false|false||Ascitesnull|Peritoneal Effusion|Finding|false|false||Ascitesnull|Hepatic|Anatomy|false|false||Portalnull|Hypertensive disease|Disorder|false|false||HTNnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Disease|Disorder|false|false||Conditionnull|Logical Condition|Finding|false|false||Conditionnull|null|Attribute|false|false||Conditionnull|Condition|Modifier|false|false||Conditionnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|Discharge instructions|Finding|false|false||Discharge Instructionsnull|hospital discharge instructions (treatment)|Procedure|false|false||Discharge Instructionsnull|null|Attribute|false|false||Discharge Instructionsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|FBXW7-AS1 gene|Finding|false|false||Dearnull|Production Class Code - Pleasure|Finding|false|false||pleasure
null|pleasurable emotion|Finding|false|false||pleasurenull|Pleasure - Animals raised for recreation|Entity|false|false||pleasurenull|care of - AddressPartType|Finding|false|false||care ofnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Abdominal Pain|Finding|false|false||stomach pain
null|Stomach ache|Finding|false|false||stomach painnull|Neoplasm of uncertain or unknown behavior of stomach|Disorder|false|false||stomach
null|Stomach Diseases|Disorder|false|false||stomach
null|Benign neoplasm of stomach|Disorder|false|false||stomach
null|Carcinoma in situ of stomach|Disorder|false|false||stomachnull|Stomach problem|Finding|false|false||stomachnull|Procedure on stomach|Procedure|false|false||stomachnull|Stomach structure|Anatomy|false|false||stomach
null|Abdomen>Stomach|Anatomy|false|false||stomach
null|Stomach|Anatomy|false|false||stomachnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Patient Outcome - Worsening|Finding|false|false||worseningnull|Worsening (qualifier value)|Modifier|false|false||worseningnull|Pathological Dilatation|Finding|false|false||distension
null|Distention|Finding|false|false||distensionnull|Paracentesis|Procedure|false|false||paracentesisnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Belly of skeletal muscle|Anatomy|false|false||bellynull|Bellis <Bellidinae>|Entity|false|false||bellynull|Lasix|Drug|false|false||Lasix
null|Lasix|Drug|false|false||Lasixnull|Aldactone|Drug|false|false||Aldactone
null|Aldactone|Drug|false|false||Aldactonenull|Help document|Finding|false|false||helpnull|Assisted (qualifier value)|Modifier|false|false||helpnull|Hypervolemia (finding)|Finding|false|false||excess fluid
null|Edema|Finding|false|false||excess fluidnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Still|Disorder|false|false||stillnull|Belly of skeletal muscle|Anatomy|false|false||bellynull|Bellis <Bellidinae>|Entity|false|false||bellynull|Different|Modifier|false|false||differentnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Lasix|Drug|false|false||lasix
null|Lasix|Drug|false|false||lasixnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Daily|Time|false|false||dailynull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Low sodium diet|Procedure|false|false||low salt dietnull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Sodium Chloride, Dietary|Drug|false|false||salt
null|sodium chloride|Drug|false|false||salt
null|Salts|Drug|false|false||saltnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Clinic|Device|false|false||clinic
null|Ambulatory Care Facilities|Device|false|false||clinicnull|Clinic|Entity|false|false||clinic
null|Ambulatory Care Facilities|Entity|false|false||clinicnull|Patient location type - Clinic|Modifier|false|false||clinic
null|Person location type - Clinic|Modifier|false|false||clinicnull|Consent Type - Colonoscopy|Procedure|false|false||colonoscopy
null|colonoscopy|Procedure|false|false||colonoscopynull|Esophagogastroduodenoscopy|Procedure|false|false||EGDnull|Course|Time|false|false||coursenull|Always - AcknowledgementCondition|Finding|false|false||always
null|All of the Time|Finding|false|false||alwaysnull|Always (frequency)|Time|false|false||alwaysnull|Vitelliform Macular Dystrophy|Disorder|false|false||bestnull|BEST1 wt Allele|Finding|false|false||best
null|BEST1 gene|Finding|false|false||bestnull|best (quality)|Modifier|false|false||bestnull|Team|Subject|false|false||Teamnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions