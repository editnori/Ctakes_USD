 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|49,58|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|49,58|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|49,63|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|83,92|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|83,92|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|83,92|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|83,92|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|83,92|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|83,97|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|115,120|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|115,120|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|115,120|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|139,142|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|139,142|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|139,142|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|139,142|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|139,142|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|150,157|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|150,157|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|159,167|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|170,179|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|170,179|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|170,179|false|false|false|C0020517|Hypersensitivity|Allergies
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|182,193|false|false|false|C0161486;C2876539|Poisoning by penicillin;Poisoning by, adverse effect of and underdosing of penicillins|Penicillins
Drug|Antibiotic|SIMPLE_SEGMENT|182,193|false|false|false|C0030842|penicillins|Penicillins
Drug|Organic Chemical|SIMPLE_SEGMENT|182,193|false|false|false|C0030842|penicillins|Penicillins
Event|Event|SIMPLE_SEGMENT|182,193|false|false|false|||Penicillins
Finding|Pathologic Function|SIMPLE_SEGMENT|182,193|false|false|false|C0413443|Adverse reaction to penicillins|Penicillins
Drug|Organic Chemical|SIMPLE_SEGMENT|196,204|false|false|false|C0699512|Dilantin|Dilantin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|196,204|false|false|false|C0699512|Dilantin|Dilantin
Event|Event|SIMPLE_SEGMENT|211,220|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|211,220|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|229,244|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|235,244|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|235,244|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|235,244|false|false|false|C5441521|Complaint (finding)|Complaint
Event|Event|SIMPLE_SEGMENT|246,254|false|false|false|||diarrhea
Finding|Finding|SIMPLE_SEGMENT|246,254|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|246,254|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Classification|SIMPLE_SEGMENT|257,262|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|263,271|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|263,271|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|275,293|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|284,293|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|284,293|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|284,293|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|284,293|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|284,293|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|SIMPLE_SEGMENT|303,310|true|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|303,310|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|303,310|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|303,310|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|303,313|true|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|303,329|true|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|303,329|true|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|314,321|true|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|314,321|true|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|314,329|true|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|322,329|true|false|false|C0221423|Illness (finding)|Illness
Finding|Functional Concept|SIMPLE_SEGMENT|358,365|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|SIMPLE_SEGMENT|358,365|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|SIMPLE_SEGMENT|358,365|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|358,365|false|false|false|C0199168|Medical service|medical
Finding|Finding|SIMPLE_SEGMENT|358,373|false|false|false|C0262926|Medical History|medical history
Event|Event|SIMPLE_SEGMENT|366,373|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|366,373|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|366,373|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|366,373|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|387,396|false|false|false|C0022107;C2700617|Irritability - emotion;Irritable Mood|irritable
Finding|Mental Process|SIMPLE_SEGMENT|387,396|false|false|false|C0022107;C2700617|Irritability - emotion;Irritable Mood|irritable
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|387,402|false|false|false|C0022104|Irritable Bowel Syndrome|irritable bowel
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|387,411|false|false|false|C0022104|Irritable Bowel Syndrome|irritable bowel syndrome
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|397,402|false|false|false|C0021853|Intestines|bowel
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|403,411|false|false|false|C0039082|Syndrome|syndrome
Event|Event|SIMPLE_SEGMENT|403,411|false|false|false|||syndrome
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|416,424|false|false|false|C0011265;C0497327|Dementia;Presenile dementia|dementia
Event|Event|SIMPLE_SEGMENT|416,424|false|false|false|||dementia
Event|Event|SIMPLE_SEGMENT|432,439|true|false|false|||reports
Event|Event|SIMPLE_SEGMENT|443,451|true|false|false|||problems
Finding|Idea or Concept|SIMPLE_SEGMENT|443,451|true|false|false|C1546466|Problems - What subject filter|problems
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|461,467|true|false|false|C0021853|Intestines|bowels
Finding|Intellectual Product|SIMPLE_SEGMENT|494,499|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Intellectual Product|SIMPLE_SEGMENT|494,505|false|false|false|C1272517|Sudden onset (contextual qualifier) (qualifier value)|acute onset
Event|Event|SIMPLE_SEGMENT|500,505|false|false|false|||onset
Event|Event|SIMPLE_SEGMENT|509,517|false|false|false|||diarrhea
Finding|Finding|SIMPLE_SEGMENT|509,517|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|509,517|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Event|Event|SIMPLE_SEGMENT|546,551|false|false|false|C0441471|Event|event
Event|Event|SIMPLE_SEGMENT|570,576|true|false|false|||travel
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|570,576|true|false|false|C0040802|travel|travel
Procedure|Health Care Activity|SIMPLE_SEGMENT|570,576|true|false|false|C1555670|travel charge|travel
Finding|Sign or Symptom|SIMPLE_SEGMENT|580,584|true|false|false|C0221423|Illness (finding)|sick
Event|Event|SIMPLE_SEGMENT|585,593|true|false|false|||contacts
Procedure|Health Care Activity|SIMPLE_SEGMENT|585,593|true|false|false|C4036459|Contacts|contacts
Event|Event|SIMPLE_SEGMENT|602,605|false|false|false|||eat
Drug|Food|SIMPLE_SEGMENT|607,618|false|false|false|C0452959|Corned beef|corned beef
Drug|Food|SIMPLE_SEGMENT|614,618|false|false|false|C0452849;C2267224;C2362309;C2702424|Beef (dietary);Beef Antigen;Beef preparation;beef allergenic extract|beef
Drug|Immunologic Factor|SIMPLE_SEGMENT|614,618|false|false|false|C0452849;C2267224;C2362309;C2702424|Beef (dietary);Beef Antigen;Beef preparation;beef allergenic extract|beef
Drug|Organic Chemical|SIMPLE_SEGMENT|614,618|false|false|false|C0452849;C2267224;C2362309;C2702424|Beef (dietary);Beef Antigen;Beef preparation;beef allergenic extract|beef
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|614,618|false|false|false|C0452849;C2267224;C2362309;C2702424|Beef (dietary);Beef Antigen;Beef preparation;beef allergenic extract|beef
Event|Event|SIMPLE_SEGMENT|614,618|false|false|false|||beef
Drug|Food|SIMPLE_SEGMENT|623,630|false|false|false|C0006619;C1095889;C2740612|cabbage allergenic extract;cabbage preparation|cabbage
Drug|Immunologic Factor|SIMPLE_SEGMENT|623,630|false|false|false|C0006619;C1095889;C2740612|cabbage allergenic extract;cabbage preparation|cabbage
Drug|Organic Chemical|SIMPLE_SEGMENT|623,630|false|false|false|C0006619;C1095889;C2740612|cabbage allergenic extract;cabbage preparation|cabbage
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|623,630|false|false|false|C0006619;C1095889;C2740612|cabbage allergenic extract;cabbage preparation|cabbage
Event|Event|SIMPLE_SEGMENT|623,630|false|false|false|||cabbage
Finding|Idea or Concept|SIMPLE_SEGMENT|638,643|false|false|false|C1550012|Local Remote Control State - Local|local
Event|Event|SIMPLE_SEGMENT|678,683|false|false|false|||noted
Attribute|Clinical Attribute|SIMPLE_SEGMENT|684,690|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|684,690|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|684,690|false|false|false|C0027497|Nausea|nausea
Event|Event|SIMPLE_SEGMENT|721,730|false|false|false|||vomitting
Finding|Sign or Symptom|SIMPLE_SEGMENT|741,756|false|false|false|C0239182|Watery diarrhoea|watery diarrhea
Event|Event|SIMPLE_SEGMENT|748,756|false|false|false|||diarrhea
Finding|Finding|SIMPLE_SEGMENT|748,756|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|748,756|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Event|Event|SIMPLE_SEGMENT|770,775|true|false|false|||fever
Finding|Finding|SIMPLE_SEGMENT|770,775|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|770,775|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Anatomy|Body Location or Region|SIMPLE_SEGMENT|777,786|true|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|SIMPLE_SEGMENT|777,795|true|false|false|C0000729|Abdominal Cramps|abdominal cramping
Event|Event|SIMPLE_SEGMENT|787,795|true|false|false|||cramping
Finding|Sign or Symptom|SIMPLE_SEGMENT|787,795|true|false|false|C0026821|Muscle Cramp|cramping
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|800,805|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|800,805|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|800,805|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Body Substance|SIMPLE_SEGMENT|813,818|false|false|false|C0015733|Feces|stool
Finding|Finding|SIMPLE_SEGMENT|832,836|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|832,836|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|832,836|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Attribute|Clinical Attribute|SIMPLE_SEGMENT|841,847|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|841,847|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|841,847|false|false|false|C0027497|Nausea|nausea
Event|Event|SIMPLE_SEGMENT|863,871|false|false|false|||improved
Event|Event|SIMPLE_SEGMENT|881,889|true|false|false|||diarrhea
Finding|Finding|SIMPLE_SEGMENT|881,889|true|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|881,889|true|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Event|Event|SIMPLE_SEGMENT|898,906|true|false|false|||improved
Drug|Organic Chemical|SIMPLE_SEGMENT|915,922|true|true|false|C0591635|Imodium|Imodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|915,922|true|true|false|C0591635|Imodium|Imodium
Event|Event|SIMPLE_SEGMENT|915,922|true|false|false|||Imodium
Event|Event|SIMPLE_SEGMENT|932,938|false|false|false|||unable
Finding|Finding|SIMPLE_SEGMENT|932,938|false|false|false|C1299582|Unable|unable
Event|Event|SIMPLE_SEGMENT|943,947|false|false|false|||keep
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|953,957|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|953,957|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|953,957|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|953,957|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Food|SIMPLE_SEGMENT|958,963|false|false|false|C0016452|Food|foods
Event|Event|SIMPLE_SEGMENT|958,963|false|false|false|||foods
Event|Event|SIMPLE_SEGMENT|968,977|false|false|false|||presented
Finding|Idea or Concept|SIMPLE_SEGMENT|968,977|false|false|false|C0449450|Presentation|presented
Drug|Food|SIMPLE_SEGMENT|997,1002|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|Vital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|997,1008|false|false|false|C0488614;C0518766|Vital signs|Vital signs
Procedure|Health Care Activity|SIMPLE_SEGMENT|997,1008|false|false|false|C0150404|Taking vital signs|Vital signs
Event|Event|SIMPLE_SEGMENT|1003,1008|false|false|false|||signs
Finding|Finding|SIMPLE_SEGMENT|1003,1008|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|1003,1008|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Event|Activity|SIMPLE_SEGMENT|1012,1019|false|false|false|C1706079||arrival
Event|Event|SIMPLE_SEGMENT|1012,1019|false|false|false|||arrival
Finding|Functional Concept|SIMPLE_SEGMENT|1012,1019|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Event|Event|SIMPLE_SEGMENT|1039,1040|false|false|false|||P
Event|Event|SIMPLE_SEGMENT|1073,1083|false|false|false|||evaluation
Finding|Idea or Concept|SIMPLE_SEGMENT|1073,1083|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|SIMPLE_SEGMENT|1073,1083|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Event|Event|SIMPLE_SEGMENT|1098,1105|false|false|false|||notable
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|1110,1116|false|false|false|C0018302|guaiac|guaiac
Drug|Organic Chemical|SIMPLE_SEGMENT|1110,1116|false|false|false|C0018302|guaiac|guaiac
Event|Event|SIMPLE_SEGMENT|1110,1116|false|false|false|||guaiac
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|1118,1126|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Event|Event|SIMPLE_SEGMENT|1118,1126|false|false|false|||positive
Finding|Classification|SIMPLE_SEGMENT|1118,1126|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|SIMPLE_SEGMENT|1118,1126|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Event|Event|SIMPLE_SEGMENT|1127,1132|false|false|false|||stool
Finding|Body Substance|SIMPLE_SEGMENT|1127,1132|false|false|false|C0015733|Feces|stool
Anatomy|Cell|SIMPLE_SEGMENT|1136,1139|false|false|false|C0023516|Leukocytes|WBC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1136,1145|false|false|false|C0023508|White Blood Cell Count procedure|WBC count
Event|Event|SIMPLE_SEGMENT|1140,1145|false|false|false|||count
Finding|Finding|SIMPLE_SEGMENT|1161,1173|false|false|false|C0151539|Blood urea increased|elevated BUN
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1170,1173|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Drug|Inorganic Chemical|SIMPLE_SEGMENT|1170,1173|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Event|Event|SIMPLE_SEGMENT|1170,1173|false|false|false|||BUN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1170,1173|false|false|false|C0005845|Blood urea nitrogen measurement|BUN
Drug|Inorganic Chemical|SIMPLE_SEGMENT|1223,1229|false|false|false|C0036082|Saline Solution|saline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1223,1229|false|false|false|C0036082|Saline Solution|saline
Event|Event|SIMPLE_SEGMENT|1223,1229|false|false|false|||saline
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1223,1229|false|false|false|C0450082|Saline method|saline
Event|Event|SIMPLE_SEGMENT|1232,1238|false|false|false|||Review
Finding|Idea or Concept|SIMPLE_SEGMENT|1232,1238|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|Review
Finding|Intellectual Product|SIMPLE_SEGMENT|1232,1238|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|Review
Finding|Functional Concept|SIMPLE_SEGMENT|1232,1241|false|false|false|C0699752|Review of|Review of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1232,1249|false|false|false|C0488564;C0488565||Review of Systems
Procedure|Health Care Activity|SIMPLE_SEGMENT|1232,1249|false|false|false|C0489633|Review of systems (procedure)|Review of Systems
Event|Event|SIMPLE_SEGMENT|1242,1249|false|false|false|||Systems
Finding|Functional Concept|SIMPLE_SEGMENT|1242,1249|false|false|false|C0449913|System|Systems
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1251,1255|false|false|false|C2598155||Pain
Finding|Functional Concept|SIMPLE_SEGMENT|1251,1255|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1251,1255|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1251,1266|false|false|false|C0030198|Pain Measurement|Pain assessment
Event|Activity|SIMPLE_SEGMENT|1256,1266|false|false|false|C1516048|Assessed|assessment
Event|Event|SIMPLE_SEGMENT|1256,1266|false|false|false|||assessment
Finding|Intellectual Product|SIMPLE_SEGMENT|1256,1266|false|false|false|C0679207|Knowledge acquisition using a method of assessment|assessment
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1256,1266|false|false|false|C0028708;C0031809;C0220825;C0542573;C0549068;C0549070;C0549071;C0549072;C0549073;C0549074;C0549075;C0549076;C0549078;C0549079;C0549080;C1161151;C1261322;C2237115|Evaluation;Evaluation procedure;Nutrition Assessment;Personal care assessment;Physical Examination;assessment of cognitive functions|assessment
Procedure|Health Care Activity|SIMPLE_SEGMENT|1256,1266|false|false|false|C0028708;C0031809;C0220825;C0542573;C0549068;C0549070;C0549071;C0549072;C0549073;C0549074;C0549075;C0549076;C0549078;C0549079;C0549080;C1161151;C1261322;C2237115|Evaluation;Evaluation procedure;Nutrition Assessment;Personal care assessment;Physical Examination;assessment of cognitive functions|assessment
Event|Activity|SIMPLE_SEGMENT|1270,1277|false|false|false|C1706079||arrival
Event|Event|SIMPLE_SEGMENT|1270,1277|false|false|false|||arrival
Finding|Functional Concept|SIMPLE_SEGMENT|1270,1277|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|1285,1290|false|false|false|C3714591|Floor (anatomic)|floor
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1301,1305|true|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|1301,1305|true|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1301,1305|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1301,1305|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|1318,1327|true|false|false|||illnesses
Finding|Sign or Symptom|SIMPLE_SEGMENT|1318,1327|true|false|false|C0221423|Illness (finding)|illnesses
Event|Event|SIMPLE_SEGMENT|1332,1338|true|false|false|||fevers
Finding|Sign or Symptom|SIMPLE_SEGMENT|1332,1338|true|false|false|C0015967|Fever|fevers
Event|Event|SIMPLE_SEGMENT|1340,1346|true|false|false|||chills
Finding|Sign or Symptom|SIMPLE_SEGMENT|1340,1346|true|false|false|C0085593|Chills|chills
Event|Event|SIMPLE_SEGMENT|1358,1364|false|false|false|||sweats
Finding|Body Substance|SIMPLE_SEGMENT|1358,1364|false|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Finding|Finding|SIMPLE_SEGMENT|1358,1364|false|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Event|Event|SIMPLE_SEGMENT|1369,1372|true|false|false|||SOB
Finding|Sign or Symptom|SIMPLE_SEGMENT|1369,1372|true|false|false|C0013404|Dyspnea|SOB
Drug|Organic Chemical|SIMPLE_SEGMENT|1374,1379|true|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1374,1379|true|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|SIMPLE_SEGMENT|1374,1379|true|false|false|||cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|1374,1379|true|false|false|C0010200|Coughing|cough
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1384,1389|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|1384,1389|true|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1384,1394|true|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1384,1394|true|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1390,1394|true|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|1390,1394|true|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1390,1394|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1390,1394|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1399,1406|true|false|false|C0042027|Urinary tract|urinary
Finding|Sign or Symptom|SIMPLE_SEGMENT|1399,1415|true|false|false|C0426359|Urinary symptoms|urinary symptoms
Event|Event|SIMPLE_SEGMENT|1407,1415|true|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|1407,1415|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|1407,1415|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|1424,1431|false|false|false|C0449913|System|systems
Event|Event|SIMPLE_SEGMENT|1432,1440|false|false|false|||reviewed
Finding|Functional Concept|SIMPLE_SEGMENT|1444,1450|false|false|false|C1561567|detail - Response Level|detail
Event|Event|SIMPLE_SEGMENT|1469,1477|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|1469,1477|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|1469,1477|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1469,1477|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|SIMPLE_SEGMENT|1481,1501|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|1486,1493|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|1486,1493|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|1486,1493|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|1486,1493|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1486,1493|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|1486,1501|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1494,1501|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1494,1501|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1494,1501|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1503,1515|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|SIMPLE_SEGMENT|1503,1515|false|false|false|||Hypertension
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1516,1524|false|false|false|C0011265;C0497327|Dementia;Presenile dementia|Dementia
Event|Event|SIMPLE_SEGMENT|1516,1524|false|false|false|||Dementia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1525,1537|false|false|false|C0029456|Osteoporosis|Osteoporosis
Event|Event|SIMPLE_SEGMENT|1525,1537|false|false|false|||Osteoporosis
Finding|Finding|SIMPLE_SEGMENT|1525,1537|false|false|false|C2911643|Encounter due to family history of osteoporosis|Osteoporosis
Finding|Finding|SIMPLE_SEGMENT|1538,1547|false|false|false|C0022107;C2700617|Irritability - emotion;Irritable Mood|Irritable
Finding|Mental Process|SIMPLE_SEGMENT|1538,1547|false|false|false|C0022107;C2700617|Irritability - emotion;Irritable Mood|Irritable
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1538,1553|false|false|false|C0022104|Irritable Bowel Syndrome|Irritable bowel
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1538,1562|false|false|false|C0022104|Irritable Bowel Syndrome|Irritable bowel syndrome
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1548,1553|false|false|false|C0021853|Intestines|bowel
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1554,1562|false|false|false|C0039082|Syndrome|syndrome
Event|Event|SIMPLE_SEGMENT|1554,1562|false|false|false|||syndrome
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|1563,1575|false|false|false|C0085662;C2004480|Macrocytosis;Macrocytosis (morphologic abnormality)|Macrocytosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1563,1575|false|false|false|C0085662;C2004480|Macrocytosis;Macrocytosis (morphologic abnormality)|Macrocytosis
Event|Event|SIMPLE_SEGMENT|1563,1575|false|false|false|||Macrocytosis
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1563,1575|false|false|false|C0684332|Macrocytosis (finding)|Macrocytosis
Event|Event|SIMPLE_SEGMENT|1587,1595|false|false|false|||etiology
Finding|Conceptual Entity|SIMPLE_SEGMENT|1587,1595|false|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|etiology
Finding|Functional Concept|SIMPLE_SEGMENT|1587,1595|false|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|etiology
Finding|Functional Concept|SIMPLE_SEGMENT|1596,1600|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1596,1604|false|false|false|C0229299|Left ear structure|Left ear
Finding|Sign or Symptom|SIMPLE_SEGMENT|1596,1604|false|false|false|C2127178|left ear symptoms (symptom)|Left ear
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1601,1604|false|false|false|C0013443;C0521421|Ear structure|ear
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1601,1604|false|false|false|C0851354|Ear and labyrinth disorders|ear
Finding|Body Substance|SIMPLE_SEGMENT|1601,1604|false|false|false|C1546608;C1550629|SpecimenType - Ear|ear
Finding|Intellectual Product|SIMPLE_SEGMENT|1601,1604|false|false|false|C1546608;C1550629|SpecimenType - Ear|ear
Finding|Finding|SIMPLE_SEGMENT|1605,1612|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|hearing
Finding|Physiologic Function|SIMPLE_SEGMENT|1605,1612|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|hearing
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1605,1617|false|false|false|C1384666|hearing impairment|hearing loss
Finding|Finding|SIMPLE_SEGMENT|1605,1617|false|false|false|C0011053;C0018772;C2029884;C3887873|Deafness;Hearing Loss;Partial Hearing Loss;hearing loss by exam|hearing loss
Event|Event|SIMPLE_SEGMENT|1613,1617|false|false|false|||loss
Finding|Finding|SIMPLE_SEGMENT|1613,1617|false|false|false|C5890125|Loss (adaptation)|loss
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1618,1624|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|1618,1624|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|1618,1624|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|1630,1642|false|false|false|||hysterectomy
Finding|Finding|SIMPLE_SEGMENT|1630,1642|false|false|false|C1548863|Consent Type - Hysterectomy|hysterectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1630,1642|false|false|false|C0020699|Hysterectomy|hysterectomy
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1643,1649|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|1643,1649|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|1643,1649|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|1655,1667|false|false|false|||appendectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1655,1667|false|false|false|C0003611;C0003612|Appendectomy;Appendectomy; for ruptured appendix with abscess or generalized peritonitis|appendectomy
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1668,1674|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|1668,1674|false|false|false|C1546481|What subject filter - Status|Status
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1680,1687|false|false|false|C0205065|Ovarian|ovarian
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1680,1692|false|false|false|C0029927|Ovarian Cysts|ovarian cyst
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1680,1700|false|false|false|C0195488|Removal of ovarian cyst|ovarian cyst removal
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|1688,1692|false|false|false|C0010709|Cyst|cyst
Event|Event|SIMPLE_SEGMENT|1688,1692|false|false|false|||cyst
Finding|Body Substance|SIMPLE_SEGMENT|1688,1692|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Finding|Intellectual Product|SIMPLE_SEGMENT|1688,1692|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1688,1700|false|false|false|C0742962|Cyst removal|cyst removal
Event|Activity|SIMPLE_SEGMENT|1693,1700|false|false|false|C1883720|Removing (action)|removal
Event|Event|SIMPLE_SEGMENT|1693,1700|false|false|false|||removal
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1693,1700|false|false|false|C0015252;C0185115;C0728940|Excision;Extraction;removal technique|removal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1701,1709|false|false|false|C0086543|Cataract|Cataract
Finding|Finding|SIMPLE_SEGMENT|1701,1709|false|false|false|C1690964|cataract on exam (physical finding)|Cataract
Finding|Finding|SIMPLE_SEGMENT|1701,1717|false|false|false|C1548833;C2186377|Consent Type - Cataract Surgery;reported history of cataract surgery|Cataract surgery
Finding|Intellectual Product|SIMPLE_SEGMENT|1701,1717|false|false|false|C1548833;C2186377|Consent Type - Cataract Surgery;reported history of cataract surgery|Cataract surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1701,1717|false|false|false|C0007389;C2939459|Cataract Extraction;Cataract surgery|Cataract surgery
Event|Event|SIMPLE_SEGMENT|1710,1717|false|false|false|||surgery
Finding|Finding|SIMPLE_SEGMENT|1710,1717|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|1710,1717|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|1710,1717|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1710,1717|false|false|false|C0543467|Operative Surgical Procedures|surgery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1718,1726|false|false|false|C0017601|Glaucoma|Glaucoma
Event|Event|SIMPLE_SEGMENT|1718,1726|false|false|false|||Glaucoma
Finding|Functional Concept|SIMPLE_SEGMENT|1729,1735|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|1729,1743|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|1736,1743|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1736,1743|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1736,1743|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1736,1743|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|1749,1755|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|1749,1755|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|1749,1755|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|1749,1755|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|1749,1763|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|1756,1763|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1756,1763|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1756,1763|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1756,1763|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Event|Event|SIMPLE_SEGMENT|1769,1777|true|false|false|||relevant
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|1785,1792|true|false|false|C1705970|Electrical Current|current
Event|Event|SIMPLE_SEGMENT|1793,1802|true|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|1793,1802|true|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|1806,1814|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|1806,1814|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|1806,1814|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1806,1814|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|1806,1819|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1806,1819|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|1815,1819|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|1815,1819|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1815,1819|false|false|false|C0582103|Medical Examination|Exam
Drug|Food|SIMPLE_SEGMENT|1821,1826|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|Vital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1821,1832|false|false|false|C0488614;C0518766|Vital signs|Vital Signs
Procedure|Health Care Activity|SIMPLE_SEGMENT|1821,1832|false|false|false|C0150404|Taking vital signs|Vital Signs
Event|Event|SIMPLE_SEGMENT|1827,1832|false|false|false|||Signs
Finding|Finding|SIMPLE_SEGMENT|1827,1832|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|Signs
Finding|Functional Concept|SIMPLE_SEGMENT|1827,1832|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|Signs
Event|Event|SIMPLE_SEGMENT|1842,1843|false|false|false|||P
Finding|Finding|SIMPLE_SEGMENT|1871,1879|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|1871,1879|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1871,1879|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|1871,1891|false|false|false|C1509143|physical examination (physical finding)|Physical examination
Procedure|Health Care Activity|SIMPLE_SEGMENT|1871,1891|false|false|false|C0031809|Physical Examination|Physical examination
Event|Activity|SIMPLE_SEGMENT|1880,1891|false|false|false|C4321457|Examination|examination
Event|Event|SIMPLE_SEGMENT|1880,1891|false|false|false|||examination
Procedure|Health Care Activity|SIMPLE_SEGMENT|1880,1891|false|false|false|C0031809;C0582103|Medical Examination;Physical Examination|examination
Finding|Classification|SIMPLE_SEGMENT|1895,1898|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Finding|Gene or Genome|SIMPLE_SEGMENT|1895,1898|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Event|Event|SIMPLE_SEGMENT|1915,1922|false|false|false|||sitting
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1929,1932|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Event|Event|SIMPLE_SEGMENT|1929,1932|false|false|false|||bed
Finding|Intellectual Product|SIMPLE_SEGMENT|1929,1932|false|false|false|C2346952|Bachelor of Education|bed
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1936,1939|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1936,1939|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1936,1939|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|1936,1939|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1936,1939|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|1936,1939|false|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|1936,1939|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1943,1948|false|false|false|C1512338|HEENT|HEENT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1950,1965|false|false|false|C1384666|hearing impairment|Hard of hearing
Finding|Finding|SIMPLE_SEGMENT|1950,1965|false|false|false|C0018772|Partial Hearing Loss|Hard of hearing
Event|Event|SIMPLE_SEGMENT|1958,1965|false|false|false|||hearing
Finding|Finding|SIMPLE_SEGMENT|1958,1965|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|hearing
Finding|Physiologic Function|SIMPLE_SEGMENT|1958,1965|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|hearing
Finding|Functional Concept|SIMPLE_SEGMENT|1967,1972|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1967,1976|false|false|false|C0229298|Right ear structure|Right ear
Finding|Sign or Symptom|SIMPLE_SEGMENT|1967,1976|false|false|false|C2127177|right ear symptoms (symptom)|Right ear
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1973,1976|false|false|false|C0013443;C0521421|Ear structure|ear
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1973,1976|false|false|false|C0851354|Ear and labyrinth disorders|ear
Event|Event|SIMPLE_SEGMENT|1973,1976|false|false|false|||ear
Finding|Body Substance|SIMPLE_SEGMENT|1973,1976|false|false|false|C1546608;C1550629|SpecimenType - Ear|ear
Finding|Intellectual Product|SIMPLE_SEGMENT|1973,1976|false|false|false|C1546608;C1550629|SpecimenType - Ear|ear
Event|Event|SIMPLE_SEGMENT|1977,1983|false|false|false|||better
Finding|Idea or Concept|SIMPLE_SEGMENT|1977,1983|false|false|false|C1550462|Observation Interpretation - better|better
Event|Event|SIMPLE_SEGMENT|1989,1993|false|false|false|||left
Finding|Functional Concept|SIMPLE_SEGMENT|1989,1993|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1997,2002|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|SIMPLE_SEGMENT|1997,2002|false|false|false|C0741025|Chest problem|Chest
Event|Event|SIMPLE_SEGMENT|2011,2023|false|false|false|||respirations
Finding|Physiologic Function|SIMPLE_SEGMENT|2011,2023|false|false|false|C0035203|Respiration|respirations
Event|Event|SIMPLE_SEGMENT|2028,2037|false|false|false|||breathing
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2064,2069|false|false|false|C0024109|Lung|Lungs
Event|Event|SIMPLE_SEGMENT|2070,2075|false|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|2070,2075|false|false|false|C1550016|Remote control command - Clear|clear
Event|Event|SIMPLE_SEGMENT|2079,2091|false|false|false|||auscultation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2079,2091|false|false|false|C0004339|Auscultation|auscultation
Event|Event|SIMPLE_SEGMENT|2119,2125|false|false|false|||rhythm
Finding|Finding|SIMPLE_SEGMENT|2119,2125|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|SIMPLE_SEGMENT|2119,2125|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Event|Event|SIMPLE_SEGMENT|2145,2152|true|false|false|||murmurs
Finding|Finding|SIMPLE_SEGMENT|2145,2152|true|false|false|C0018808|Heart murmur|murmurs
Event|Event|SIMPLE_SEGMENT|2156,2163|true|false|false|||gallops
Event|Event|SIMPLE_SEGMENT|2165,2168|false|false|false|||JVP
Finding|Finding|SIMPLE_SEGMENT|2165,2168|false|false|false|C0428897|Jugular venous pressure|JVP
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2180,2187|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2180,2187|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Finding|Finding|SIMPLE_SEGMENT|2180,2187|false|false|false|C0941288|Abdomen problem|Abdomen
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2196,2201|false|false|false|C0021853|Intestines|bowel
Finding|Finding|SIMPLE_SEGMENT|2196,2208|false|false|false|C0232693|Bowel sounds|bowel sounds
Event|Event|SIMPLE_SEGMENT|2202,2208|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2202,2208|false|false|false|C0037709||sounds
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2210,2214|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|SIMPLE_SEGMENT|2210,2214|false|false|false|||Soft
Event|Event|SIMPLE_SEGMENT|2216,2225|false|false|false|||nontender
Event|Event|SIMPLE_SEGMENT|2227,2239|false|false|false|||nondistended
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2244,2255|false|false|false|C0015385;C0278454|All extremities;Limb structure|Extremities
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2260,2265|true|false|false|C0003086;C0003087;C4284979|Ankle;Ankle joint structure;Lower extremity>Ankle|ankle
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|2260,2265|true|false|false|C0003086;C0003087;C4284979|Ankle;Ankle joint structure;Lower extremity>Ankle|ankle
Finding|Pathologic Function|SIMPLE_SEGMENT|2260,2271|true|false|false|C0235439|Ankle edema (finding)|ankle edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2266,2271|true|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|2266,2271|true|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|2266,2271|true|false|false|C0013604|Edema|edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2282,2287|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|2282,2287|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2282,2287|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|2282,2287|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|2282,2287|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|2282,2287|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|2282,2287|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|2289,2297|false|false|false|||oriented
Event|Event|SIMPLE_SEGMENT|2313,2320|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|2313,2320|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2313,2320|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|2313,2320|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Idea or Concept|SIMPLE_SEGMENT|2355,2359|true|true|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|2355,2359|true|true|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|2355,2359|true|true|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2360,2371|true|true|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2360,2371|true|true|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|2360,2371|true|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|2360,2371|true|true|false|C4284232|Medications|medications
Event|Event|SIMPLE_SEGMENT|2375,2384|true|false|false|||specifics
Event|Event|SIMPLE_SEGMENT|2385,2391|true|false|false|||timing
Finding|Intellectual Product|SIMPLE_SEGMENT|2385,2391|true|false|false|C1704250|Timing, LOINC Axis 3|timing
Finding|Finding|SIMPLE_SEGMENT|2396,2409|false|false|false|C2133635|recent events relating to health|recent events
Event|Event|SIMPLE_SEGMENT|2403,2409|false|false|false|||events
Event|Event|SIMPLE_SEGMENT|2403,2409|false|false|false|C0441471|Event|events
Finding|Mental Process|SIMPLE_SEGMENT|2415,2432|false|false|false|C0025265|Memory, Short-Term|short-term memory
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2415,2443|false|false|false|C0701811|Poor short-term memory|short-term memory impairment
Finding|Idea or Concept|SIMPLE_SEGMENT|2421,2425|false|false|false|C0233324;C1705313|Term (lexical);Term Birth|term
Finding|Organism Function|SIMPLE_SEGMENT|2421,2425|false|false|false|C0233324;C1705313|Term (lexical);Term Birth|term
Finding|Finding|SIMPLE_SEGMENT|2426,2432|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Intellectual Product|SIMPLE_SEGMENT|2426,2432|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Mental Process|SIMPLE_SEGMENT|2426,2432|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2426,2443|false|false|false|C0233794|Memory impairment|memory impairment
Finding|Sign or Symptom|SIMPLE_SEGMENT|2426,2443|false|false|false|C0542476|Forgetful|memory impairment
Event|Event|SIMPLE_SEGMENT|2433,2443|false|false|false|||impairment
Finding|Finding|SIMPLE_SEGMENT|2433,2443|false|false|false|C0221099;C0684336|Impaired;Impaired health|impairment
Finding|Functional Concept|SIMPLE_SEGMENT|2433,2443|false|false|false|C0221099;C0684336|Impaired;Impaired health|impairment
Event|Event|SIMPLE_SEGMENT|2445,2451|false|false|false|||Speech
Finding|Organism Function|SIMPLE_SEGMENT|2445,2451|false|false|false|C0037817|Speech|Speech
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2445,2451|false|false|false|C0846595|Speech assessment|Speech
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2457,2465|false|false|false|C2706915||language
Event|Event|SIMPLE_SEGMENT|2457,2465|false|false|false|||language
Finding|Intellectual Product|SIMPLE_SEGMENT|2457,2465|false|false|false|C0033348|Programming Languages|language
Event|Event|SIMPLE_SEGMENT|2470,2476|false|false|false|||normal
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2481,2486|false|false|false|C0004936;C1306597|Mental disorders;Psychiatric problem|Psych
Event|Event|SIMPLE_SEGMENT|2481,2486|false|false|false|||Psych
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2488,2498|false|false|false|C0550215||Appearance
Event|Event|SIMPLE_SEGMENT|2488,2498|false|false|false|||Appearance
Procedure|Health Care Activity|SIMPLE_SEGMENT|2488,2498|false|false|false|C2051406|patient appearance regarding mental status exam|Appearance
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2500,2508|false|false|false|C2707008||behavior
Event|Event|SIMPLE_SEGMENT|2500,2508|false|false|false|||behavior
Finding|Behavior|SIMPLE_SEGMENT|2500,2508|false|false|false|C0004927|Behavior|behavior
Event|Event|SIMPLE_SEGMENT|2514,2520|false|false|false|||affect
Event|Event|SIMPLE_SEGMENT|2525,2531|false|false|false|||normal
Procedure|Health Care Activity|SIMPLE_SEGMENT|2555,2564|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Event|Event|SIMPLE_SEGMENT|2565,2569|false|false|false|||Labs
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2565,2569|false|false|false|C0587081|Laboratory test finding|Labs
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2583,2588|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|2583,2588|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2583,2588|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|2589,2592|false|false|false|C0023516|Leukocytes|WBC
Event|Event|SIMPLE_SEGMENT|2615,2621|false|false|false|||Lymphs
Finding|Body Substance|SIMPLE_SEGMENT|2615,2621|false|false|false|C0024202|Lymph|Lymphs
Drug|Antibiotic|SIMPLE_SEGMENT|2626,2631|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2626,2631|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|SIMPLE_SEGMENT|2626,2631|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2636,2639|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Finding|Gene or Genome|SIMPLE_SEGMENT|2636,2639|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Anatomy|Cell|SIMPLE_SEGMENT|2663,2666|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2663,2666|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2663,2666|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2673,2676|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2673,2676|false|false|false|C0019046|Hemoglobin|Hgb
Event|Event|SIMPLE_SEGMENT|2673,2676|false|false|false|||Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|2673,2676|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2673,2676|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2682,2685|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2682,2685|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|2691,2694|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|2691,2694|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2691,2694|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2691,2694|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2691,2694|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|2699,2702|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2699,2702|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|2699,2702|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|2699,2702|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|2699,2702|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2699,2702|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2709,2713|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Event|Event|SIMPLE_SEGMENT|2728,2731|false|false|false|||Plt
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2728,2731|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2749,2754|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|2749,2754|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|2749,2754|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|2749,2762|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2749,2762|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2749,2762|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2755,2762|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|2755,2762|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2755,2762|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|2755,2762|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2755,2762|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2755,2762|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|2809,2813|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2809,2813|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2809,2813|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2827,2830|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2827,2830|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|2827,2830|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|2827,2830|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|2827,2830|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|2827,2830|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|2827,2830|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2827,2830|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|2834,2837|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2834,2837|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2834,2837|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2834,2837|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|2834,2837|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|2834,2837|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|2834,2837|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2841,2848|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|SIMPLE_SEGMENT|2841,2848|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2865,2871|false|false|false|C0023764|lipase|Lipase
Drug|Enzyme|SIMPLE_SEGMENT|2865,2871|false|false|false|C0023764|lipase|Lipase
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2865,2871|false|false|false|C0023764|lipase|Lipase
Event|Event|SIMPLE_SEGMENT|2865,2871|false|false|false|||Lipase
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2865,2871|false|false|false|C0373670|Lipase measurement|Lipase
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2875,2882|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2875,2882|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2875,2882|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Event|Event|SIMPLE_SEGMENT|2875,2882|false|false|false|||Albumin
Finding|Gene or Genome|SIMPLE_SEGMENT|2875,2882|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Finding|Physiologic Function|SIMPLE_SEGMENT|2875,2882|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2875,2882|false|false|false|C0201838|Albumin measurement|Albumin
Finding|Body Substance|SIMPLE_SEGMENT|2902,2907|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|2902,2907|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|2902,2907|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Finding|SIMPLE_SEGMENT|2902,2913|false|false|false|C0278030|Color of urine|URINE Color
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2908,2913|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|Color
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|2908,2913|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|Color
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2941,2946|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Event|Event|SIMPLE_SEGMENT|2941,2946|false|false|false|||Blood
Finding|Body Substance|SIMPLE_SEGMENT|2941,2946|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Event|Event|SIMPLE_SEGMENT|2947,2950|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|2947,2950|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2951,2958|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Drug|Inorganic Chemical|SIMPLE_SEGMENT|2951,2958|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2951,2958|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Event|Event|SIMPLE_SEGMENT|2959,2962|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|2959,2962|false|false|false|C5848551|Neg - answer|NEG
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2963,2970|false|false|false|C0033684|Proteins|Protein
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2963,2970|false|false|false|C0033684|Proteins|Protein
Event|Event|SIMPLE_SEGMENT|2963,2970|false|false|false|||Protein
Finding|Conceptual Entity|SIMPLE_SEGMENT|2963,2970|false|false|false|C1521746|Protein Info|Protein
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2963,2970|false|false|false|C0202202|Protein measurement|Protein
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2974,2981|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|2974,2981|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2974,2981|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|2974,2981|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2974,2981|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2974,2981|false|false|false|C0337438|Glucose measurement|Glucose
Event|Event|SIMPLE_SEGMENT|2982,2985|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|2982,2985|false|false|false|C5848551|Neg - answer|NEG
Drug|Organic Chemical|SIMPLE_SEGMENT|2986,2992|false|false|false|C0022634|Ketones|Ketone
Event|Event|SIMPLE_SEGMENT|2993,2996|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|2993,2996|false|false|false|C5848551|Neg - answer|NEG
Event|Event|SIMPLE_SEGMENT|3006,3009|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|3006,3009|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|SIMPLE_SEGMENT|3018,3021|false|false|false|C5848551|Neg - answer|NEG
Event|Event|SIMPLE_SEGMENT|3035,3038|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|3035,3038|false|false|false|C5848551|Neg - answer|NEG
Anatomy|Cell|SIMPLE_SEGMENT|3039,3042|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3039,3042|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3039,3042|false|false|false|C0014792|Erythrocytes|RBC
Anatomy|Cell|SIMPLE_SEGMENT|3045,3048|false|false|false|C0023516|Leukocytes|WBC
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3059,3062|true|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|MOD
Event|Event|SIMPLE_SEGMENT|3059,3062|true|false|false|||MOD
Drug|Food|SIMPLE_SEGMENT|3064,3069|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Immunologic Factor|SIMPLE_SEGMENT|3064,3069|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|3064,3069|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3064,3069|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3075,3078|true|false|false|C0267963|Exocrine pancreatic insufficiency|Epi
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3075,3078|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3075,3078|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Hormone|SIMPLE_SEGMENT|3075,3078|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Organic Chemical|SIMPLE_SEGMENT|3075,3078|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3075,3078|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Event|Event|SIMPLE_SEGMENT|3075,3078|true|false|false|||Epi
Finding|Gene or Genome|SIMPLE_SEGMENT|3075,3078|true|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|Epi
Finding|Intellectual Product|SIMPLE_SEGMENT|3075,3078|true|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|Epi
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3075,3078|true|false|false|C0162734;C3641909|Echo-Planar Imaging;Electronic Portal Imaging|Epi
Event|Event|SIMPLE_SEGMENT|3115,3127|false|false|false|||Microbiology
Finding|Functional Concept|SIMPLE_SEGMENT|3115,3127|false|false|false|C0025953;C1571921;C4049106|Microbiological;Microbiology - Laboratory Class;Microbiology Diagnostic Service Section ID|Microbiology
Finding|Intellectual Product|SIMPLE_SEGMENT|3115,3127|false|false|false|C0025953;C1571921;C4049106|Microbiological;Microbiology - Laboratory Class;Microbiology Diagnostic Service Section ID|Microbiology
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3115,3127|false|false|false|C0085672|Microbiology procedure|Microbiology
Finding|Body Substance|SIMPLE_SEGMENT|3133,3138|false|false|false|C0015733|Feces|Stool
Event|Event|SIMPLE_SEGMENT|3139,3147|false|false|false|||Cultures
Finding|Idea or Concept|SIMPLE_SEGMENT|3139,3147|false|true|false|C0010453|Culture (Anthropological)|Cultures
Finding|Body Substance|SIMPLE_SEGMENT|3161,3166|false|false|false|C0015733|Feces|STOOL
Finding|Finding|SIMPLE_SEGMENT|3161,3182|false|false|false|C0426740|Consistency of stool|STOOL     CONSISTENCY
Event|Event|SIMPLE_SEGMENT|3196,3202|false|false|false|||Source
Finding|Finding|SIMPLE_SEGMENT|3196,3202|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|Source
Finding|Functional Concept|SIMPLE_SEGMENT|3196,3202|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|Source
Finding|Intellectual Product|SIMPLE_SEGMENT|3196,3202|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|Source
Event|Event|SIMPLE_SEGMENT|3205,3210|false|false|false|||Stool
Finding|Body Substance|SIMPLE_SEGMENT|3205,3210|false|false|false|C0015733|Feces|Stool
Finding|Body Substance|SIMPLE_SEGMENT|3216,3221|false|false|false|C0015733|Feces|FECAL
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3216,3229|false|false|false|C0430414|Stool culture|FECAL CULTURE
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3222,3229|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|SIMPLE_SEGMENT|3222,3229|false|false|false|||CULTURE
Finding|Functional Concept|SIMPLE_SEGMENT|3222,3229|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|3222,3229|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3222,3229|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|SIMPLE_SEGMENT|3231,3238|false|false|false|||Pending
Finding|Idea or Concept|SIMPLE_SEGMENT|3231,3238|false|false|false|C1691786;C1704475|Pending - Allergy Clinical Status;Pending - referral status|Pending
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3245,3266|false|false|false|C1294214|Campylobacter culture|CAMPYLOBACTER CULTURE
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3259,3266|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|SIMPLE_SEGMENT|3259,3266|false|false|false|||CULTURE
Finding|Functional Concept|SIMPLE_SEGMENT|3259,3266|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|3259,3266|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3259,3266|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|SIMPLE_SEGMENT|3268,3275|false|false|false|||Pending
Finding|Idea or Concept|SIMPLE_SEGMENT|3268,3275|false|false|false|C1691786;C1704475|Pending - Allergy Clinical Status;Pending - referral status|Pending
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3282,3309|false|false|false|C0314765|Clostridium difficile toxin|CLOSTRIDIUM DIFFICILE TOXIN
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3282,3309|false|false|false|C0314765|Clostridium difficile toxin|CLOSTRIDIUM DIFFICILE TOXIN
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|3282,3309|false|false|false|C0314765|Clostridium difficile toxin|CLOSTRIDIUM DIFFICILE TOXIN
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3282,3311|false|false|false|C0055948|tcdA protein, Clostridium difficile|CLOSTRIDIUM DIFFICILE TOXIN A
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3282,3311|false|false|false|C0055948|tcdA protein, Clostridium difficile|CLOSTRIDIUM DIFFICILE TOXIN A
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|3282,3311|false|false|false|C0055948|tcdA protein, Clostridium difficile|CLOSTRIDIUM DIFFICILE TOXIN A
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3304,3309|false|false|false|C0040549|Toxin|TOXIN
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|3304,3309|false|false|false|C0040549|Toxin|TOXIN
Event|Event|SIMPLE_SEGMENT|3304,3309|false|false|false|||TOXIN
Event|Event|SIMPLE_SEGMENT|3310,3311|false|false|false|||A
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3316,3320|false|false|false|C4318744|Test - temporal region|TEST
Event|Event|SIMPLE_SEGMENT|3316,3320|false|false|false|||TEST
Finding|Functional Concept|SIMPLE_SEGMENT|3316,3320|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|TEST
Finding|Intellectual Product|SIMPLE_SEGMENT|3316,3320|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|TEST
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3316,3320|false|false|false|C0456984|Test Result|TEST
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3316,3320|false|false|false|C0022885|Laboratory Procedures|TEST
Event|Event|SIMPLE_SEGMENT|3322,3327|false|false|false|||Final
Finding|Idea or Concept|SIMPLE_SEGMENT|3322,3327|false|false|false|C1546485|Diagnosis Type - Final|Final
Finding|Body Substance|SIMPLE_SEGMENT|3340,3345|true|false|false|C0015733|Feces|Feces
Event|Event|SIMPLE_SEGMENT|3346,3354|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|3346,3354|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|3346,3354|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3346,3354|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|SIMPLE_SEGMENT|3346,3358|false|false|false|C0205160|Negative|negative for
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3371,3376|false|false|false|C0040549|Toxin|toxin
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|3371,3376|false|false|false|C0040549|Toxin|toxin
Event|Event|SIMPLE_SEGMENT|3377,3378|false|false|false|||A
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3386,3389|false|false|false|C0014661;C5400664|Endocrine Therapy-Induced Alopecia;Equine Infectious Anemia|EIA
Event|Event|SIMPLE_SEGMENT|3386,3389|false|false|false|||EIA
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3386,3389|false|false|false|C0086231|Enzyme Immunoassay|EIA
Finding|Conceptual Entity|SIMPLE_SEGMENT|3404,3413|false|false|false|C1514811;C1561577;C1706462;C3244318;C4266518|Bibliographic Reference;Reference - HL7UpdateMode;Reference - MdfHmdMetSourceType;Reference Object;Reference source|Reference
Finding|Idea or Concept|SIMPLE_SEGMENT|3404,3413|false|false|false|C1514811;C1561577;C1706462;C3244318;C4266518|Bibliographic Reference;Reference - HL7UpdateMode;Reference - MdfHmdMetSourceType;Reference Object;Reference source|Reference
Finding|Intellectual Product|SIMPLE_SEGMENT|3404,3413|false|false|false|C1514811;C1561577;C1706462;C3244318;C4266518|Bibliographic Reference;Reference - HL7UpdateMode;Reference - MdfHmdMetSourceType;Reference Object;Reference source|Reference
Finding|Intellectual Product|SIMPLE_SEGMENT|3414,3419|false|false|false|C3542016|Concept model range (foundation metadata concept)|Range
Event|Event|SIMPLE_SEGMENT|3420,3428|false|false|false|||Negative
Finding|Classification|SIMPLE_SEGMENT|3420,3428|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Finding|Finding|SIMPLE_SEGMENT|3420,3428|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3420,3428|false|false|false|C5237010|Expression Negative|Negative
Finding|Body Substance|SIMPLE_SEGMENT|3438,3443|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Functional Concept|SIMPLE_SEGMENT|3438,3443|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Intellectual Product|SIMPLE_SEGMENT|3438,3443|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Event|Event|SIMPLE_SEGMENT|3444,3452|false|false|false|||Cultures
Finding|Idea or Concept|SIMPLE_SEGMENT|3444,3452|false|true|false|C0010453|Culture (Anthropological)|Cultures
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3470,3475|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3470,3475|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3470,3475|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|3476,3479|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|3485,3488|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3485,3488|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3485,3488|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3495,3498|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3495,3498|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|3495,3498|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3495,3498|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3504,3507|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3504,3507|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|3514,3517|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|3514,3517|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3514,3517|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3514,3517|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3514,3517|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|3521,3524|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3521,3524|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|3521,3524|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|3521,3524|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|3521,3524|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3521,3524|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3531,3535|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3550,3553|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3570,3575|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3570,3575|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3570,3575|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|3570,3583|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3570,3583|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3570,3583|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3576,3583|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|3576,3583|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3576,3583|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|3576,3583|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3576,3583|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3576,3583|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3628,3632|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3628,3632|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3628,3632|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3657,3662|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3657,3662|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3657,3662|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3663,3666|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3663,3666|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|3663,3666|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|3663,3666|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|3663,3666|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|3663,3666|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|3663,3666|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3663,3666|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|3670,3673|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3670,3673|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3670,3673|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3670,3673|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|3670,3673|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|3670,3673|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|3670,3673|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3677,3684|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|SIMPLE_SEGMENT|3677,3684|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3712,3717|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3712,3717|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3712,3717|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3744,3749|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3744,3749|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3744,3749|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3744,3757|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3750,3757|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|3750,3757|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3750,3757|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3750,3757|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|3750,3757|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|3750,3757|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|3750,3757|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3750,3757|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|3801,3804|false|false|false|C0022104;C0432306|Ichthyosis Bullosa of Siemens;Irritable Bowel Syndrome|IBS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3801,3804|false|false|false|C0022104;C0432306|Ichthyosis Bullosa of Siemens;Irritable Bowel Syndrome|IBS
Event|Event|SIMPLE_SEGMENT|3801,3804|false|false|false|||IBS
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|3809,3817|false|false|false|C0011265;C0497327|Dementia;Presenile dementia|Dementia
Event|Event|SIMPLE_SEGMENT|3809,3817|false|false|false|||Dementia
Event|Event|SIMPLE_SEGMENT|3822,3831|false|false|false|||presented
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3850,3856|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|3850,3856|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|3850,3856|false|false|false|C0027497|Nausea|nausea
Event|Event|SIMPLE_SEGMENT|3858,3866|false|false|false|||vomiting
Finding|Sign or Symptom|SIMPLE_SEGMENT|3858,3866|false|false|false|C0042963|Vomiting|vomiting
Event|Event|SIMPLE_SEGMENT|3882,3890|false|false|false|||diarrhea
Finding|Finding|SIMPLE_SEGMENT|3882,3890|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|3882,3890|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3908,3918|false|false|false|C0011175|Dehydration|dehydrated
Event|Event|SIMPLE_SEGMENT|3908,3918|false|false|false|||dehydrated
Event|Event|SIMPLE_SEGMENT|3922,3931|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|3922,3931|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Intellectual Product|SIMPLE_SEGMENT|3937,3942|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3937,3956|false|false|false|C0022660|Kidney Failure, Acute|acute renal failure
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3943,3948|false|false|false|C0022646|Kidney|renal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3943,3948|false|false|false|C0042075|Urologic Diseases|renal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3943,3956|false|false|false|C0035078|Kidney Failure|renal failure
Event|Event|SIMPLE_SEGMENT|3949,3956|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|3949,3956|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|3949,3956|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|3949,3956|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|SIMPLE_SEGMENT|3961,3972|false|false|false|||symptomatic
Finding|Functional Concept|SIMPLE_SEGMENT|3961,3972|false|false|false|C0231220|Symptomatic|symptomatic
Event|Event|SIMPLE_SEGMENT|3974,3985|false|false|false|||orthostasis
Finding|Finding|SIMPLE_SEGMENT|3974,3985|false|false|false|C0149746;C1535893|Orthostasis;Orthostatic intolerance|orthostasis
Finding|Sign or Symptom|SIMPLE_SEGMENT|3974,3985|false|false|false|C0149746;C1535893|Orthostasis;Orthostatic intolerance|orthostasis
Event|Event|SIMPLE_SEGMENT|3995,4002|false|false|false|||treated
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4008,4011|false|false|false|C0016520|Structure of interventricular foramen|IVF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4008,4011|false|false|false|C2751898|Ventricular Fibrillation, Paroxysmal Familial, 1|IVF
Event|Event|SIMPLE_SEGMENT|4008,4011|false|false|false|||IVF
Finding|Gene or Genome|SIMPLE_SEGMENT|4008,4011|false|false|false|C1419864;C4321334|SCN5A gene;SCN5A wt Allele|IVF
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4008,4011|false|false|false|C0015915;C0872104|Assisted Reproductive Technologies;Fertilization in Vitro|IVF
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4016,4021|false|false|false|C0021853|Intestines|bowel
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4022,4026|false|false|false|C1742913|REST protein, human|rest
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4022,4026|false|false|false|C1742913|REST protein, human|rest
Event|Event|SIMPLE_SEGMENT|4022,4026|false|false|false|||rest
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|4022,4026|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Gene or Genome|SIMPLE_SEGMENT|4022,4026|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Molecular Function|SIMPLE_SEGMENT|4022,4026|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4030,4040|false|false|false|C0009450|Communicable Diseases|Infectious
Event|Event|SIMPLE_SEGMENT|4041,4045|false|false|false|||work
Event|Occupational Activity|SIMPLE_SEGMENT|4041,4045|false|false|false|C0043227|Work|work
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4041,4048|false|false|false|C0750430|Work-up|work up
Event|Event|SIMPLE_SEGMENT|4065,4073|false|false|false|||returned
Finding|Classification|SIMPLE_SEGMENT|4074,4082|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|4074,4082|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4074,4082|false|false|false|C5237010|Expression Negative|negative
Event|Event|SIMPLE_SEGMENT|4088,4100|false|false|false|||presentation
Finding|Idea or Concept|SIMPLE_SEGMENT|4088,4100|false|false|false|C0449450|Presentation|presentation
Event|Event|SIMPLE_SEGMENT|4110,4120|false|false|false|||consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|4110,4120|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|4110,4125|false|false|false|C0332290|Consistent with|consistent with
Event|Event|SIMPLE_SEGMENT|4126,4135|false|false|false|||norovirus
Event|Event|SIMPLE_SEGMENT|4153,4161|false|false|false|||advanced
Drug|Food|SIMPLE_SEGMENT|4164,4168|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|SIMPLE_SEGMENT|4164,4168|false|false|false|||diet
Finding|Functional Concept|SIMPLE_SEGMENT|4164,4168|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|SIMPLE_SEGMENT|4164,4168|false|false|false|C0012159|Diet therapy|diet
Event|Event|SIMPLE_SEGMENT|4173,4181|false|false|false|||diarrhea
Finding|Finding|SIMPLE_SEGMENT|4173,4181|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|4173,4181|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Event|Event|SIMPLE_SEGMENT|4182,4190|false|false|false|||improved
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4193,4198|false|false|false|C0022646|Kidney|Renal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4193,4198|false|false|false|C0042075|Urologic Diseases|Renal
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4193,4207|false|false|false|C0232804|Renal function|Renal function
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4193,4207|false|false|false|C0022662|Kidney Function Tests|Renal function
Event|Event|SIMPLE_SEGMENT|4199,4207|false|false|false|||function
Finding|Finding|SIMPLE_SEGMENT|4199,4207|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|4199,4207|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|4199,4207|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|SIMPLE_SEGMENT|4199,4207|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Event|Event|SIMPLE_SEGMENT|4208,4216|false|false|false|||returned
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4221,4229|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|SIMPLE_SEGMENT|4221,4229|false|false|false|||baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|4221,4229|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4235,4238|false|false|false|C0016520|Structure of interventricular foramen|IVF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4235,4238|false|false|false|C2751898|Ventricular Fibrillation, Paroxysmal Familial, 1|IVF
Event|Event|SIMPLE_SEGMENT|4235,4238|false|false|false|||IVF
Finding|Gene or Genome|SIMPLE_SEGMENT|4235,4238|false|false|false|C1419864;C4321334|SCN5A gene;SCN5A wt Allele|IVF
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4235,4238|false|false|false|C0015915;C0872104|Assisted Reproductive Technologies;Fertilization in Vitro|IVF
Event|Event|SIMPLE_SEGMENT|4250,4260|true|false|false|||tolerating
Finding|Finding|SIMPLE_SEGMENT|4263,4273|true|false|false|C0301572|Bland diet|bland diet
Drug|Food|SIMPLE_SEGMENT|4269,4273|true|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|SIMPLE_SEGMENT|4269,4273|true|false|false|||diet
Finding|Functional Concept|SIMPLE_SEGMENT|4269,4273|true|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|SIMPLE_SEGMENT|4269,4273|true|false|false|C0012159|Diet therapy|diet
Event|Event|SIMPLE_SEGMENT|4287,4295|true|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|4287,4295|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|4287,4298|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Event|Event|SIMPLE_SEGMENT|4299,4310|true|false|false|||orthostasis
Finding|Finding|SIMPLE_SEGMENT|4299,4310|true|false|false|C0149746;C1535893|Orthostasis;Orthostatic intolerance|orthostasis
Finding|Sign or Symptom|SIMPLE_SEGMENT|4299,4310|true|false|false|C0149746;C1535893|Orthostasis;Orthostatic intolerance|orthostasis
Finding|Idea or Concept|SIMPLE_SEGMENT|4318,4321|true|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|4318,4321|true|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|4325,4334|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|4325,4334|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|4325,4334|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|4325,4334|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|4325,4334|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|4345,4349|false|false|false|||seen
Event|Event|SIMPLE_SEGMENT|4361,4365|false|false|false|||felt
Event|Event|SIMPLE_SEGMENT|4379,4383|true|false|false|||safe
Finding|Intellectual Product|SIMPLE_SEGMENT|4379,4383|true|false|false|C4684764|SAFE-Biopharma Standard|safe
Event|Event|SIMPLE_SEGMENT|4388,4397|true|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|4388,4397|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|4388,4397|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|4388,4397|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|4388,4397|true|false|false|C0030685|Patient Discharge|discharge
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4388,4402|true|false|false|C0184713|Discharge to home|discharge home
Event|Event|SIMPLE_SEGMENT|4398,4402|true|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|4398,4402|true|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|4398,4402|true|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|4398,4402|true|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|4412,4420|true|false|false|||services
Event|Occupational Activity|SIMPLE_SEGMENT|4412,4420|true|false|false|C0557854|Services|services
Procedure|Health Care Activity|SIMPLE_SEGMENT|4412,4420|true|false|false|C1704289|Clinical Service|services
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4426,4440|false|false|false|C0009763|Conjunctivitis|Conjunctivitis
Event|Event|SIMPLE_SEGMENT|4426,4440|false|false|false|||Conjunctivitis
Finding|Functional Concept|SIMPLE_SEGMENT|4442,4446|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4442,4450|false|false|false|C0229090|Left eye structure|left eye
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4442,4450|false|false|false|C2141124|examination of left eye|left eye
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4447,4450|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4447,4450|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4447,4450|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4447,4450|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Finding|Body Substance|SIMPLE_SEGMENT|4447,4450|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Finding|SIMPLE_SEGMENT|4447,4450|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Intellectual Product|SIMPLE_SEGMENT|4447,4450|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Finding|SIMPLE_SEGMENT|4460,4464|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|4460,4464|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|4460,4464|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|SIMPLE_SEGMENT|4468,4477|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|4468,4477|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|4482,4490|false|false|false|||reported
Event|Event|SIMPLE_SEGMENT|4498,4505|false|false|false|||treated
Drug|Antibiotic|SIMPLE_SEGMENT|4511,4523|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|SIMPLE_SEGMENT|4511,4523|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|SIMPLE_SEGMENT|4511,4523|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4524,4529|false|false|false|C0991568|Drops - Drug Form|drops
Event|Event|SIMPLE_SEGMENT|4524,4529|false|false|false|||drops
Finding|Functional Concept|SIMPLE_SEGMENT|4534,4538|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4534,4542|false|false|false|C0229090|Left eye structure|left eye
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4534,4542|false|false|false|C2141124|examination of left eye|left eye
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4539,4542|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4539,4542|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4539,4542|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4539,4542|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Event|Event|SIMPLE_SEGMENT|4539,4542|false|false|false|||eye
Finding|Body Substance|SIMPLE_SEGMENT|4539,4542|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Finding|SIMPLE_SEGMENT|4539,4542|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Intellectual Product|SIMPLE_SEGMENT|4539,4542|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4544,4558|false|false|false|C0009763|Conjunctivitis|conjunctivitis
Event|Event|SIMPLE_SEGMENT|4544,4558|false|false|false|||conjunctivitis
Finding|Idea or Concept|SIMPLE_SEGMENT|4574,4581|false|false|false|C0549178|Continuous|ongoing
Event|Event|SIMPLE_SEGMENT|4582,4590|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|4582,4590|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|4582,4590|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|SIMPLE_SEGMENT|4599,4606|false|false|false|||started
Drug|Antibiotic|SIMPLE_SEGMENT|4611,4623|false|false|false|C0014806|erythromycin|erythromycin
Drug|Organic Chemical|SIMPLE_SEGMENT|4611,4623|false|false|false|C0014806|erythromycin|erythromycin
Event|Event|SIMPLE_SEGMENT|4611,4623|false|false|false|||erythromycin
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4634,4642|false|false|false|C0028912|Ointments|ointment
Event|Event|SIMPLE_SEGMENT|4634,4642|false|false|false|||ointment
Event|Event|SIMPLE_SEGMENT|4653,4664|false|false|false|||improvement
Finding|Conceptual Entity|SIMPLE_SEGMENT|4653,4664|false|false|false|C2986411|Improvement|improvement
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4669,4681|false|false|false|C0009758|conjunctiva|conjunctival
Finding|Functional Concept|SIMPLE_SEGMENT|4669,4681|false|false|false|C1522483|Conjunctival Route of Administration|conjunctival
Finding|Finding|SIMPLE_SEGMENT|4669,4691|false|false|false|C1761613|Conjunctival hyperemia|conjunctival injection
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4682,4691|false|false|false|C1272883|Injection|injection
Event|Event|SIMPLE_SEGMENT|4682,4691|false|false|false|||injection
Finding|Functional Concept|SIMPLE_SEGMENT|4682,4691|false|false|false|C1828121|Injection Route of Administration|injection
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4682,4691|false|false|false|C0021485;C1533685|Injection of therapeutic agent;Injection procedure|injection
Event|Event|SIMPLE_SEGMENT|4702,4712|true|false|false|||instructed
Event|Event|SIMPLE_SEGMENT|4716,4723|true|false|false|||monitor
Event|Event|SIMPLE_SEGMENT|4733,4742|true|false|false|||worsening
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4746,4749|true|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4746,4749|true|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4746,4749|true|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4746,4749|true|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Finding|Body Substance|SIMPLE_SEGMENT|4746,4749|true|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Finding|SIMPLE_SEGMENT|4746,4749|true|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Intellectual Product|SIMPLE_SEGMENT|4746,4749|true|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Finding|SIMPLE_SEGMENT|4746,4758|true|false|false|C0586406|Eye symptom|eye symptoms
Event|Event|SIMPLE_SEGMENT|4750,4758|true|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|4750,4758|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|4750,4758|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|SIMPLE_SEGMENT|4767,4776|false|false|false|||scheduled
Finding|Functional Concept|SIMPLE_SEGMENT|4781,4787|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|4781,4787|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|SIMPLE_SEGMENT|4781,4790|false|false|false|C0589120|Follow-up status|follow up
Procedure|Health Care Activity|SIMPLE_SEGMENT|4781,4790|false|false|false|C1522577|follow-up|follow up
Event|Event|SIMPLE_SEGMENT|4788,4790|false|false|false|||up
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4801,4804|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|4801,4804|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4801,4804|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4801,4804|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|4801,4804|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|4801,4804|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|4801,4804|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4801,4804|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|4801,4804|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|4801,4804|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|4801,4804|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|SIMPLE_SEGMENT|4833,4840|true|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|4833,4840|true|false|false|C0392747|Changing|changes
Finding|Intellectual Product|SIMPLE_SEGMENT|4853,4860|true|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|4853,4860|true|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4861,4871|true|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|4861,4871|true|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|4861,4871|true|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|4873,4880|false|false|false|||regimen
Finding|Intellectual Product|SIMPLE_SEGMENT|4873,4880|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4873,4880|false|false|false|C0040808|Treatment Protocols|regimen
Event|Occupational Activity|SIMPLE_SEGMENT|4884,4888|false|false|false|C0009219|Coding|Code
Finding|Intellectual Product|SIMPLE_SEGMENT|4884,4888|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|Code
Procedure|Health Care Activity|SIMPLE_SEGMENT|4884,4895|false|false|false|C0742531|CODE STATUS|Code Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4889,4895|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|4889,4895|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|4889,4895|false|false|false|C1546481|What subject filter - Status|Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4897,4900|false|false|false|C4285234||DNR
Drug|Antibiotic|SIMPLE_SEGMENT|4897,4900|false|false|false|C0011015|daunorubicin|DNR
Drug|Organic Chemical|SIMPLE_SEGMENT|4897,4900|false|false|false|C0011015|daunorubicin|DNR
Event|Event|SIMPLE_SEGMENT|4897,4900|false|false|false|||DNR
Finding|Finding|SIMPLE_SEGMENT|4897,4900|false|false|false|C0079252;C0582114|Do not resuscitate status;Do-Not-Resuscitate Orders|DNR
Finding|Intellectual Product|SIMPLE_SEGMENT|4897,4900|false|false|false|C0079252;C0582114|Do not resuscitate status;Do-Not-Resuscitate Orders|DNR
Event|Event|SIMPLE_SEGMENT|4905,4914|false|false|false|||confirmed
Event|Event|SIMPLE_SEGMENT|4918,4927|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|4918,4927|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Body Substance|SIMPLE_SEGMENT|4933,4940|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|4933,4940|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|4933,4940|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4950,4953|false|false|false|C0162531|Hereditary Coproporphyria|HCP
Event|Event|SIMPLE_SEGMENT|4950,4953|false|false|false|||HCP
Finding|Gene or Genome|SIMPLE_SEGMENT|4950,4953|false|false|false|C1335283;C1412376;C1413681;C1705637;C5780748|AMBP gene;AMBP wt Allele;CPOX gene;PTPN6 gene;PTPN6 wt Allele|HCP
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4958,4969|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4958,4969|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|4958,4969|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|4958,4969|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|4958,4982|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|SIMPLE_SEGMENT|4973,4982|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|4973,4982|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Event|Event|SIMPLE_SEGMENT|4985,4989|false|false|false|||list
Finding|Intellectual Product|SIMPLE_SEGMENT|4985,4989|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|SIMPLE_SEGMENT|4990,4999|false|false|false|||confirmed
Event|Event|SIMPLE_SEGMENT|5013,5022|false|false|false|||caregiver
Event|Event|SIMPLE_SEGMENT|5026,5035|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|5026,5035|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Drug|Organic Chemical|SIMPLE_SEGMENT|5054,5061|false|false|false|C1330412|Namenda|Namenda
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5054,5061|false|false|false|C1330412|Namenda|Namenda
Drug|Organic Chemical|SIMPLE_SEGMENT|5074,5081|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5074,5081|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|5101,5111|false|false|false|C0244404|raloxifene|Raloxifene
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5101,5111|false|false|false|C0244404|raloxifene|Raloxifene
Event|Event|SIMPLE_SEGMENT|5101,5111|false|false|false|||Raloxifene
Drug|Organic Chemical|SIMPLE_SEGMENT|5113,5119|false|false|false|C0720318|Evista|Evista
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5113,5119|false|false|false|C0720318|Evista|Evista
Drug|Organic Chemical|SIMPLE_SEGMENT|5136,5148|false|false|false|C0301532|Multivitamin preparation|Multivitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5136,5148|false|false|false|C0301532|Multivitamin preparation|Multivitamin
Drug|Vitamin|SIMPLE_SEGMENT|5136,5148|false|false|false|C0301532|Multivitamin preparation|Multivitamin
Drug|Organic Chemical|SIMPLE_SEGMENT|5155,5166|false|false|false|C0017718|glucosamine|Glucosamine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5155,5166|false|false|false|C0017718|glucosamine|Glucosamine
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5171,5178|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|5171,5178|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5171,5178|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5171,5178|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|5171,5178|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|5171,5178|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|5171,5178|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5171,5178|false|false|false|C0201925|Calcium measurement|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5171,5189|false|false|false|C3540037|CALCIUM SUPPLEMENTS|Calcium supplement
Drug|Vitamin|SIMPLE_SEGMENT|5171,5189|false|false|false|C3540037|CALCIUM SUPPLEMENTS|Calcium supplement
Drug|Food|SIMPLE_SEGMENT|5179,5189|false|false|false|C0242295|Dietary Supplements|supplement
Event|Event|SIMPLE_SEGMENT|5179,5189|false|false|false|||supplement
Finding|Functional Concept|SIMPLE_SEGMENT|5179,5189|false|false|false|C1549514;C1947943;C2348609|Supplement;Supplement (document);Supplement - Diet Code Specification Type|supplement
Finding|Idea or Concept|SIMPLE_SEGMENT|5179,5189|false|false|false|C1549514;C1947943;C2348609|Supplement;Supplement (document);Supplement - Diet Code Specification Type|supplement
Finding|Intellectual Product|SIMPLE_SEGMENT|5179,5189|false|false|false|C1549514;C1947943;C2348609|Supplement;Supplement (document);Supplement - Diet Code Specification Type|supplement
Drug|Organic Chemical|SIMPLE_SEGMENT|5190,5205|false|false|false|C0008318|cholecalciferol|Cholecalciferol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5190,5205|false|false|false|C0008318|cholecalciferol|Cholecalciferol
Drug|Vitamin|SIMPLE_SEGMENT|5190,5205|false|false|false|C0008318|cholecalciferol|Cholecalciferol
Event|Event|SIMPLE_SEGMENT|5190,5205|false|false|false|||Cholecalciferol
Drug|Organic Chemical|SIMPLE_SEGMENT|5190,5218|false|false|false|C0008318|cholecalciferol|Cholecalciferol (Vitamin D3)
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5190,5218|false|false|false|C0008318|cholecalciferol|Cholecalciferol (Vitamin D3)
Drug|Vitamin|SIMPLE_SEGMENT|5190,5218|false|false|false|C0008318|cholecalciferol|Cholecalciferol (Vitamin D3)
Drug|Organic Chemical|SIMPLE_SEGMENT|5207,5214|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5207,5214|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|SIMPLE_SEGMENT|5207,5214|false|false|false|C0042890|Vitamins|Vitamin
Drug|Organic Chemical|SIMPLE_SEGMENT|5207,5217|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|Vitamin D3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5207,5217|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|Vitamin D3
Drug|Vitamin|SIMPLE_SEGMENT|5207,5217|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|Vitamin D3
Drug|Organic Chemical|SIMPLE_SEGMENT|5240,5253|false|false|false|C0003968|ascorbic acid|Ascorbic Acid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5240,5253|false|false|false|C0003968|ascorbic acid|Ascorbic Acid
Drug|Vitamin|SIMPLE_SEGMENT|5240,5253|false|false|false|C0003968|ascorbic acid|Ascorbic Acid
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5240,5253|false|false|false|C0201898|Ascorbic acid measurement|Ascorbic Acid
Event|Event|SIMPLE_SEGMENT|5249,5253|false|false|false|||Acid
Event|Event|SIMPLE_SEGMENT|5272,5281|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|5272,5281|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|5272,5281|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|5272,5281|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|5272,5281|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|5272,5293|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5282,5293|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5282,5293|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|5282,5293|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|5282,5293|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|5298,5307|false|false|false|C0527316|donepezil|donepezil
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5298,5307|false|false|false|C0527316|donepezil|donepezil
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5313,5319|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5333,5339|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|5333,5339|false|false|false|||Tablet
Drug|Organic Chemical|SIMPLE_SEGMENT|5366,5373|false|false|false|C1330412|Namenda|Namenda
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5366,5373|false|false|false|C1330412|Namenda|Namenda
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5380,5386|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5400,5406|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|5400,5406|false|false|false|||Tablet
Drug|Organic Chemical|SIMPLE_SEGMENT|5423,5430|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5423,5430|false|false|false|C0004057|aspirin|aspirin
Event|Event|SIMPLE_SEGMENT|5423,5430|false|false|false|||aspirin
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5438,5444|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|5438,5444|false|false|false|||Tablet
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5446,5453|false|false|false|C1545665|Views delayed|Delayed
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5446,5461|false|false|false|C1707664|Delayed Release Dosage Form|Delayed Release
Event|Event|SIMPLE_SEGMENT|5454,5461|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|5454,5461|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|5454,5461|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5454,5461|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Event|Event|SIMPLE_SEGMENT|5469,5472|false|false|false|||Sig
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5483,5489|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|5483,5489|false|false|false|||Tablet
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5491,5498|false|false|false|C1545665|Views delayed|Delayed
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5491,5506|false|false|false|C1707664|Delayed Release Dosage Form|Delayed Release
Event|Event|SIMPLE_SEGMENT|5499,5506|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|5499,5506|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|5499,5506|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5499,5506|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Finding|Intellectual Product|SIMPLE_SEGMENT|5517,5521|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5517,5527|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|SIMPLE_SEGMENT|5524,5527|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|5524,5527|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|SIMPLE_SEGMENT|5534,5544|false|false|false|C0244404|raloxifene|raloxifene
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5534,5544|false|false|false|C0244404|raloxifene|raloxifene
Event|Event|SIMPLE_SEGMENT|5534,5544|false|false|false|||raloxifene
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5551,5557|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|5558,5561|false|false|false|||Sig
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5571,5577|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Intellectual Product|SIMPLE_SEGMENT|5581,5585|false|false|false|C1720092|Once - dosing instruction fragment|once
Finding|Intellectual Product|SIMPLE_SEGMENT|5588,5592|false|false|false|C1561540|Transaction counts and value totals - week|week
Drug|Organic Chemical|SIMPLE_SEGMENT|5599,5611|false|false|false|C0301532|Multivitamin preparation|multivitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5599,5611|false|false|false|C0301532|Multivitamin preparation|multivitamin
Drug|Vitamin|SIMPLE_SEGMENT|5599,5611|false|false|false|C0301532|Multivitamin preparation|multivitamin
Event|Event|SIMPLE_SEGMENT|5599,5611|false|false|false|||multivitamin
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5613,5617|false|false|false|C0226896|Oral cavity|Oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5613,5617|false|false|false|C1272919|Oral Dosage Form|Oral
Event|Event|SIMPLE_SEGMENT|5613,5617|false|false|false|||Oral
Finding|Finding|SIMPLE_SEGMENT|5613,5617|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Finding|Functional Concept|SIMPLE_SEGMENT|5613,5617|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Drug|Organic Chemical|SIMPLE_SEGMENT|5621,5632|false|false|false|C0017718|glucosamine|Glucosamine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5621,5632|false|false|false|C0017718|glucosamine|Glucosamine
Event|Event|SIMPLE_SEGMENT|5621,5632|false|false|false|||Glucosamine
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5634,5638|false|false|false|C0226896|Oral cavity|Oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5634,5638|false|false|false|C1272919|Oral Dosage Form|Oral
Event|Event|SIMPLE_SEGMENT|5634,5638|false|false|false|||Oral
Finding|Finding|SIMPLE_SEGMENT|5634,5638|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Finding|Functional Concept|SIMPLE_SEGMENT|5634,5638|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Drug|Organic Chemical|SIMPLE_SEGMENT|5642,5649|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5642,5649|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|SIMPLE_SEGMENT|5642,5649|false|false|false|C0042890|Vitamins|Vitamin
Event|Event|SIMPLE_SEGMENT|5642,5649|false|false|false|||Vitamin
Drug|Hormone|SIMPLE_SEGMENT|5642,5651|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|SIMPLE_SEGMENT|5642,5651|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5642,5651|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|SIMPLE_SEGMENT|5642,5651|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5642,5651|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5653,5657|false|false|false|C0226896|Oral cavity|Oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5653,5657|false|false|false|C1272919|Oral Dosage Form|Oral
Finding|Finding|SIMPLE_SEGMENT|5653,5657|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Finding|Functional Concept|SIMPLE_SEGMENT|5653,5657|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Drug|Organic Chemical|SIMPLE_SEGMENT|5661,5674|false|false|false|C0003968|ascorbic acid|ascorbic acid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5661,5674|false|false|false|C0003968|ascorbic acid|ascorbic acid
Drug|Vitamin|SIMPLE_SEGMENT|5661,5674|false|false|false|C0003968|ascorbic acid|ascorbic acid
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5661,5674|false|false|false|C0201898|Ascorbic acid measurement|ascorbic acid
Event|Event|SIMPLE_SEGMENT|5670,5674|false|false|false|||acid
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5676,5680|false|false|false|C0226896|Oral cavity|Oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5676,5680|false|false|false|C1272919|Oral Dosage Form|Oral
Finding|Finding|SIMPLE_SEGMENT|5676,5680|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Finding|Functional Concept|SIMPLE_SEGMENT|5676,5680|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5684,5691|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|5684,5691|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5684,5691|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5684,5691|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|5684,5691|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|5684,5691|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|5684,5691|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5684,5691|false|false|false|C0201925|Calcium measurement|Calcium
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5697,5701|false|false|false|C0226896|Oral cavity|Oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5697,5701|false|false|false|C1272919|Oral Dosage Form|Oral
Finding|Finding|SIMPLE_SEGMENT|5697,5701|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Finding|Functional Concept|SIMPLE_SEGMENT|5697,5701|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Drug|Antibiotic|SIMPLE_SEGMENT|5706,5718|false|false|false|C0014806|erythromycin|erythromycin
Drug|Organic Chemical|SIMPLE_SEGMENT|5706,5718|false|false|false|C0014806|erythromycin|erythromycin
Event|Event|SIMPLE_SEGMENT|5706,5718|false|false|false|||erythromycin
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5737,5745|false|false|false|C0028912|Ointments|Ointment
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5761,5771|false|false|false|C0015392|Eye|Ophthalmic
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5761,5771|false|false|false|C2347396|Ophthalmic Dosage Form|Ophthalmic
Finding|Functional Concept|SIMPLE_SEGMENT|5761,5771|false|false|false|C1522230|Ophthalmic Route of Administration|Ophthalmic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5777,5782|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|SIMPLE_SEGMENT|5785,5788|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|5785,5788|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|5801,5806|false|false|false|||apply
Finding|Functional Concept|SIMPLE_SEGMENT|5810,5814|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5810,5818|false|false|false|C0229090|Left eye structure|left eye
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5810,5818|false|false|false|C2141124|examination of left eye|left eye
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5815,5818|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5815,5818|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5815,5818|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5815,5818|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Event|Event|SIMPLE_SEGMENT|5815,5818|false|false|false|||eye
Finding|Body Substance|SIMPLE_SEGMENT|5815,5818|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Finding|SIMPLE_SEGMENT|5815,5818|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Intellectual Product|SIMPLE_SEGMENT|5815,5818|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Functional Concept|SIMPLE_SEGMENT|5851,5855|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Finding|Gene or Genome|SIMPLE_SEGMENT|5851,5855|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Finding|Idea or Concept|SIMPLE_SEGMENT|5857,5864|false|false|false|C0807726|refill|Refills
Event|Event|SIMPLE_SEGMENT|5872,5881|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|5872,5881|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|5872,5881|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|5872,5881|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|5872,5881|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5872,5893|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|5872,5893|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5882,5893|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|5882,5893|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|5882,5893|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|SIMPLE_SEGMENT|5895,5899|false|false|false|||Home
Finding|Idea or Concept|SIMPLE_SEGMENT|5895,5899|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|5895,5899|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|5895,5899|false|false|false|C1553498|home health encounter|Home
Event|Event|SIMPLE_SEGMENT|5902,5911|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|5902,5911|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|5902,5911|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|5902,5911|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|5902,5911|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|5902,5921|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5912,5921|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|5912,5921|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|5912,5921|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|5912,5921|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5912,5921|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Intellectual Product|SIMPLE_SEGMENT|5933,5949|false|false|false|C1314977|Gastrointestinal attachment|Gastrointestinal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5950,5955|false|false|false|C0042769;C0042776;C0319157|AS virus;Virus;Virus Diseases|Virus
Disorder|Virus|SIMPLE_SEGMENT|5950,5955|false|false|false|C0042769;C0042776;C0319157|AS virus;Virus;Virus Diseases|Virus
Event|Event|SIMPLE_SEGMENT|5950,5955|false|false|false|||Virus
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5956,5967|false|false|false|C0011175;C2062903|Dehydration;dehydration (Na, H2O)|Dehydration
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|5956,5967|false|false|false|C0011175;C2062903|Dehydration;dehydration (Na, H2O)|Dehydration
Event|Event|SIMPLE_SEGMENT|5956,5967|false|false|false|||Dehydration
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5956,5967|false|false|false|C4284399|Dehydration procedure|Dehydration
Finding|Functional Concept|SIMPLE_SEGMENT|5969,5980|false|false|false|C0231220|Symptomatic|Symptomatic
Event|Event|SIMPLE_SEGMENT|5981,5992|false|false|false|||orthostasis
Finding|Finding|SIMPLE_SEGMENT|5981,5992|false|false|false|C0149746;C1535893|Orthostasis;Orthostatic intolerance|orthostasis
Finding|Sign or Symptom|SIMPLE_SEGMENT|5981,5992|false|false|false|C0149746;C1535893|Orthostasis;Orthostatic intolerance|orthostasis
Event|Event|SIMPLE_SEGMENT|5996,6005|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|5996,6005|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|5996,6005|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|5996,6005|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|5996,6005|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6006,6015|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6006,6015|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|6006,6015|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|6006,6015|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|6017,6023|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6017,6030|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|6017,6030|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6024,6030|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|6024,6030|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|6032,6037|false|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|6032,6037|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|6042,6050|false|false|false|||coherent
Finding|Finding|SIMPLE_SEGMENT|6042,6050|false|false|false|C4068804|Coherent|coherent
Event|Event|SIMPLE_SEGMENT|6052,6057|false|false|false|||Level
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6052,6074|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|6052,6074|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|SIMPLE_SEGMENT|6061,6074|false|false|false|||Consciousness
Finding|Finding|SIMPLE_SEGMENT|6061,6074|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|6061,6074|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6076,6081|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|6076,6081|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6076,6081|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|6076,6081|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|6076,6081|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|6076,6081|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|6076,6081|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|6086,6097|false|false|false|||interactive
Finding|Functional Concept|SIMPLE_SEGMENT|6086,6097|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|6099,6107|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|6099,6107|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|6099,6107|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6108,6114|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|6108,6114|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|6108,6114|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|6116,6126|false|false|false|||Ambulatory
Finding|Functional Concept|SIMPLE_SEGMENT|6116,6126|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|6116,6126|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|6116,6126|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|6116,6126|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|SIMPLE_SEGMENT|6129,6140|false|false|false|||Independent
Finding|Finding|SIMPLE_SEGMENT|6129,6140|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|SIMPLE_SEGMENT|6129,6140|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Event|Event|SIMPLE_SEGMENT|6145,6154|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|6145,6154|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6145,6154|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6145,6154|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6145,6154|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6145,6167|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|6145,6167|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|6145,6167|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6155,6167|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|6155,6167|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|6155,6167|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Event|Event|SIMPLE_SEGMENT|6178,6186|false|false|false|||admitted
Finding|Intellectual Product|SIMPLE_SEGMENT|6195,6200|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Sign or Symptom|SIMPLE_SEGMENT|6211,6218|false|false|false|C0221423|Illness (finding)|illness
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6224,6235|false|false|false|C0011175;C2062903|Dehydration;dehydration (Na, H2O)|dehydration
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|6224,6235|false|false|false|C0011175;C2062903|Dehydration;dehydration (Na, H2O)|dehydration
Event|Event|SIMPLE_SEGMENT|6224,6235|false|false|false|||dehydration
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6224,6235|false|false|false|C4284399|Dehydration procedure|dehydration
Finding|Finding|SIMPLE_SEGMENT|6247,6253|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|6247,6253|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6263,6268|false|false|false|C0042769;C0042776;C0319157|AS virus;Virus;Virus Diseases|virus
Disorder|Virus|SIMPLE_SEGMENT|6263,6268|false|false|false|C0042769;C0042776;C0319157|AS virus;Virus;Virus Diseases|virus
Event|Event|SIMPLE_SEGMENT|6263,6268|false|false|false|||virus
Event|Event|SIMPLE_SEGMENT|6288,6298|false|false|false|||contagious
Event|Event|SIMPLE_SEGMENT|6315,6322|false|false|false|||treated
Drug|Substance|SIMPLE_SEGMENT|6331,6337|false|false|false|C0302908|Liquid substance|fluids
Event|Event|SIMPLE_SEGMENT|6331,6337|false|false|false|||fluids
Finding|Body Substance|SIMPLE_SEGMENT|6331,6337|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6331,6337|false|false|false|C0016286|Fluid Therapy|fluids
Event|Event|SIMPLE_SEGMENT|6342,6352|false|false|false|||supportive
Finding|Conceptual Entity|SIMPLE_SEGMENT|6342,6352|false|false|false|C1521721|Supportive assistance|supportive
Event|Activity|SIMPLE_SEGMENT|6354,6358|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|6354,6358|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|6354,6358|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|6354,6358|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Event|Event|SIMPLE_SEGMENT|6364,6375|false|false|false|||improvement
Finding|Conceptual Entity|SIMPLE_SEGMENT|6364,6375|false|false|false|C2986411|Improvement|improvement
Event|Event|SIMPLE_SEGMENT|6384,6392|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|6384,6392|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|6384,6392|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|SIMPLE_SEGMENT|6409,6413|false|false|false|||seen
Finding|Finding|SIMPLE_SEGMENT|6418,6426|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Finding|Functional Concept|SIMPLE_SEGMENT|6418,6426|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|6418,6426|false|false|false|C0031809|Physical Examination|physical
Finding|Intellectual Product|SIMPLE_SEGMENT|6418,6434|false|false|false|C1547999|Diagnostic Service Section ID - Physical Therapy|physical therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6418,6434|false|false|false|C0949766|Physical therapy|physical therapy
Event|Event|SIMPLE_SEGMENT|6427,6434|false|false|false|||therapy
Finding|Finding|SIMPLE_SEGMENT|6427,6434|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|SIMPLE_SEGMENT|6427,6434|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6427,6434|false|false|false|C0087111|Therapeutic procedure|therapy
Event|Event|SIMPLE_SEGMENT|6439,6444|false|false|false|||agree
Event|Event|SIMPLE_SEGMENT|6458,6462|false|false|false|||safe
Finding|Intellectual Product|SIMPLE_SEGMENT|6458,6462|false|false|false|C4684764|SAFE-Biopharma Standard|safe
Event|Event|SIMPLE_SEGMENT|6466,6472|false|false|false|||return
Event|Event|SIMPLE_SEGMENT|6473,6477|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|6473,6477|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|6473,6477|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|6473,6477|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|6490,6499|false|false|false|||encourage
Event|Event|SIMPLE_SEGMENT|6504,6508|false|false|false|||take
Finding|Finding|SIMPLE_SEGMENT|6512,6516|false|false|false|C4281574|Much|much
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6517,6521|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6517,6521|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|6517,6521|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|6517,6521|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|SIMPLE_SEGMENT|6522,6531|false|false|false|||hydration
Finding|Finding|SIMPLE_SEGMENT|6522,6531|false|false|false|C1321013;C4520800|Hydration;Hydration status|hydration
Finding|Physiologic Function|SIMPLE_SEGMENT|6522,6531|false|false|false|C1321013;C4520800|Hydration;Hydration status|hydration
Finding|Finding|SIMPLE_SEGMENT|6535,6543|false|false|false|C0332149|Possible|possible
Event|Event|SIMPLE_SEGMENT|6549,6557|false|false|false|||continue
Event|Event|SIMPLE_SEGMENT|6558,6567|false|false|false|||advancing
Drug|Food|SIMPLE_SEGMENT|6573,6577|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|SIMPLE_SEGMENT|6573,6577|false|false|false|||diet
Finding|Functional Concept|SIMPLE_SEGMENT|6573,6577|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|SIMPLE_SEGMENT|6573,6577|false|false|false|C0012159|Diet therapy|diet
Event|Event|SIMPLE_SEGMENT|6581,6590|false|false|false|||tolerated
Event|Event|SIMPLE_SEGMENT|6600,6604|false|false|false|||keep
Event|Activity|SIMPLE_SEGMENT|6611,6622|false|false|false|C0003629|Appointments|appointment
Event|Event|SIMPLE_SEGMENT|6611,6622|false|false|false|||appointment
Finding|Finding|SIMPLE_SEGMENT|6666,6669|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|6666,6669|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6670,6682|false|false|false|C5886759|Prescription (attribute)|prescription
Event|Event|SIMPLE_SEGMENT|6670,6682|false|false|false|||prescription
Finding|Intellectual Product|SIMPLE_SEGMENT|6670,6682|false|false|false|C1521941|prescription document|prescription
Procedure|Health Care Activity|SIMPLE_SEGMENT|6670,6682|false|false|false|C0033080|Prescription (procedure)|prescription
Event|Event|SIMPLE_SEGMENT|6686,6690|false|false|false|||help
Event|Event|SIMPLE_SEGMENT|6691,6696|false|false|false|||treat
Finding|Functional Concept|SIMPLE_SEGMENT|6701,6705|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6701,6709|false|false|false|C0229090|Left eye structure|left eye
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6701,6709|false|false|false|C2141124|examination of left eye|left eye
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6706,6709|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6706,6709|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6706,6709|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6706,6709|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Event|Event|SIMPLE_SEGMENT|6706,6709|false|false|false|||eye
Finding|Body Substance|SIMPLE_SEGMENT|6706,6709|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Finding|SIMPLE_SEGMENT|6706,6709|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Intellectual Product|SIMPLE_SEGMENT|6706,6709|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6711,6725|false|false|false|C0009763|Conjunctivitis|conjunctivitis
Event|Event|SIMPLE_SEGMENT|6711,6725|false|false|false|||conjunctivitis
Event|Event|SIMPLE_SEGMENT|6734,6742|false|false|false|||continue
Event|Event|SIMPLE_SEGMENT|6743,6748|false|false|false|||using
Drug|Antibiotic|SIMPLE_SEGMENT|6753,6765|false|false|false|C0014806|erythromycin|erythromycin
Drug|Organic Chemical|SIMPLE_SEGMENT|6753,6765|false|false|false|C0014806|erythromycin|erythromycin
Drug|Clinical Drug|SIMPLE_SEGMENT|6753,6774|false|false|false|C1248462||erythromycin ointment
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6766,6774|false|false|false|C0028912|Ointments|ointment
Event|Event|SIMPLE_SEGMENT|6766,6774|false|false|false|||ointment
Event|Event|SIMPLE_SEGMENT|6804,6811|true|false|false|||develop
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6816,6820|true|false|false|C5779629|Eruption of skin (disorder)|rash
Event|Event|SIMPLE_SEGMENT|6816,6820|true|false|false|||rash
Finding|Pathologic Function|SIMPLE_SEGMENT|6816,6820|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|SIMPLE_SEGMENT|6816,6820|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6829,6833|true|false|false|C0015450;C4266571|Face;Head>Face|face
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6829,6833|true|false|false|C3160739|FANCONI ANEMIA, COMPLEMENTATION GROUP E|face
Event|Event|SIMPLE_SEGMENT|6829,6833|true|false|false|||face
Finding|Gene or Genome|SIMPLE_SEGMENT|6829,6833|true|false|false|C1414531;C1423759;C2828055|ELOVL6 gene;FANCE gene;FANCE wt Allele|face
Event|Event|SIMPLE_SEGMENT|6836,6842|true|false|false|||fevers
Finding|Sign or Symptom|SIMPLE_SEGMENT|6836,6842|true|false|false|C0015967|Fever|fevers
Finding|Functional Concept|SIMPLE_SEGMENT|6844,6850|false|false|false|C0234621|Visual|visual
Finding|Finding|SIMPLE_SEGMENT|6844,6858|false|false|false|C0750280|Visual changes|visual changes
Event|Event|SIMPLE_SEGMENT|6851,6858|false|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|6851,6858|false|false|false|C0392747|Changing|changes
Event|Event|SIMPLE_SEGMENT|6862,6871|false|false|false|||worsening
Finding|Idea or Concept|SIMPLE_SEGMENT|6862,6871|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6875,6878|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6875,6878|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6875,6878|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6875,6878|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Finding|Body Substance|SIMPLE_SEGMENT|6875,6878|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Finding|SIMPLE_SEGMENT|6875,6878|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Intellectual Product|SIMPLE_SEGMENT|6875,6878|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Finding|SIMPLE_SEGMENT|6875,6887|false|false|false|C0586406|Eye symptom|eye symptoms
Event|Event|SIMPLE_SEGMENT|6879,6887|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|6879,6887|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|6879,6887|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|SIMPLE_SEGMENT|6896,6900|false|false|false|||call
Finding|Functional Concept|SIMPLE_SEGMENT|6896,6900|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Gene or Genome|SIMPLE_SEGMENT|6896,6900|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Intellectual Product|SIMPLE_SEGMENT|6896,6900|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Mental Process|SIMPLE_SEGMENT|6896,6900|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6907,6910|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|6907,6910|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6907,6910|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6907,6910|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|6907,6910|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|6907,6910|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|6907,6910|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6907,6910|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|6907,6910|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|6907,6910|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|6907,6910|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|SIMPLE_SEGMENT|6914,6920|false|false|false|||return
Finding|Intellectual Product|SIMPLE_SEGMENT|6925,6931|false|false|false|C1546403;C1546845;C1547230;C1561556|Admission Type - Urgent;Certification patient type - Urgent;Triage Code - Urgent;Visit Priority Code - Urgent|urgent
Event|Event|SIMPLE_SEGMENT|6932,6942|false|false|false|||evaluation
Finding|Idea or Concept|SIMPLE_SEGMENT|6932,6942|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|SIMPLE_SEGMENT|6932,6942|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Event|Event|SIMPLE_SEGMENT|6969,6973|true|false|false|||made
Event|Event|SIMPLE_SEGMENT|6978,6985|true|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|6978,6985|true|false|false|C0392747|Changing|changes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6994,7005|true|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6994,7005|true|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|6994,7005|true|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|6994,7005|true|false|false|C4284232|Medications|medications
Procedure|Health Care Activity|SIMPLE_SEGMENT|7008,7016|true|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7017,7029|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|7017,7029|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|7017,7029|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

