 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|46,55|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|46,55|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|46,60|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|80,89|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|80,89|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|80,94|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|136,139|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|147,154|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|147,154|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|156,164|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|167,176|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|167,176|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|167,176|false|false|false|C0020517|Hypersensitivity|Allergies
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|179,189|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|179,189|false|false|false|C0065374|lisinopril|lisinopril
Event|Event|SIMPLE_SEGMENT|179,189|false|false|false|||lisinopril
Event|Event|SIMPLE_SEGMENT|192,201|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|192,201|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|210,225|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|216,225|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|216,225|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|216,225|false|false|false|C5441521|Complaint (finding)|Complaint
Anatomy|Body Location or Region|SIMPLE_SEGMENT|227,232|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|SIMPLE_SEGMENT|227,232|false|false|false|C0741025|Chest problem|Chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|227,237|false|false|false|C2926613||Chest Pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|227,237|false|false|false|C0008031|Chest Pain|Chest Pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|233,237|false|true|false|C2598155||Pain
Finding|Functional Concept|SIMPLE_SEGMENT|233,237|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|233,237|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Classification|SIMPLE_SEGMENT|240,245|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|246,254|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|246,254|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|258,276|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|267,276|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|267,276|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|267,276|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|267,276|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|267,276|false|false|false|C0184661|Interventional procedure|Procedure
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|278,286|false|false|false|C0015259|Exercise|Exercise
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|278,286|false|false|false|C1522704|Exercise Pain Management|Exercise
Event|Event|SIMPLE_SEGMENT|287,303|false|false|false|||Echocardiography
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|287,303|false|false|false|C0013516;C2729489|Echocardiography;echocardiography service|Echocardiography
Procedure|Health Care Activity|SIMPLE_SEGMENT|287,303|false|false|false|C0013516;C2729489|Echocardiography;echocardiography service|Echocardiography
Event|Event|SIMPLE_SEGMENT|307,314|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|307,314|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|307,314|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|307,314|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|307,317|false|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|307,333|false|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|307,333|false|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|318,325|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|318,325|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|318,333|false|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|326,333|false|false|false|C0221423|Illness (finding)|Illness
Finding|Finding|SIMPLE_SEGMENT|339,342|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|pmh
Finding|Finding|SIMPLE_SEGMENT|343,349|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|343,349|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|356,359|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|356,359|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|356,359|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|356,359|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|356,359|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|356,359|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|356,359|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|356,359|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|SIMPLE_SEGMENT|364,368|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|364,368|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Event|Event|SIMPLE_SEGMENT|394,401|false|false|false|||chronic
Finding|Intellectual Product|SIMPLE_SEGMENT|394,401|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|394,401|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Event|Occupational Activity|SIMPLE_SEGMENT|411,418|false|false|false|C1273870|Management procedure|managed
Attribute|Clinical Attribute|SIMPLE_SEGMENT|419,425|false|false|false|C2926611||angina
Event|Event|SIMPLE_SEGMENT|419,425|false|false|false|||angina
Finding|Finding|SIMPLE_SEGMENT|419,425|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Finding|Sign or Symptom|SIMPLE_SEGMENT|419,425|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|432,435|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|432,435|false|false|false|||HTN
Event|Event|SIMPLE_SEGMENT|444,452|false|false|false|||presents
Event|Event|SIMPLE_SEGMENT|459,467|false|false|false|||atypical
Finding|Finding|SIMPLE_SEGMENT|459,467|false|false|false|C0741302|atypia morphology|atypical
Finding|Sign or Symptom|SIMPLE_SEGMENT|459,478|false|false|false|C0262384|Atypical chest pain|atypical chest pain
Anatomy|Body Location or Region|SIMPLE_SEGMENT|468,473|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|468,473|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|468,478|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|468,478|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|474,478|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|474,478|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|474,478|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|474,478|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Body Substance|SIMPLE_SEGMENT|486,493|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|486,493|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|486,493|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Functional Concept|SIMPLE_SEGMENT|486,497|false|false|false|C0332310|Has patient|Patient has
Event|Event|SIMPLE_SEGMENT|498,505|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|498,505|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|498,505|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|498,505|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|498,508|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|509,512|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|509,512|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|509,512|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|509,512|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|509,512|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|509,512|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|509,512|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|509,512|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Anatomy|Body Location or Region|SIMPLE_SEGMENT|526,532|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|526,532|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Event|Event|SIMPLE_SEGMENT|533,537|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|533,537|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|544,547|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|544,547|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|SIMPLE_SEGMENT|544,547|false|false|false|||LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|544,547|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Event|SIMPLE_SEGMENT|599,607|false|false|false|||admitted
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|619,625|false|false|false|C4255010||NSTEMI
Event|Event|SIMPLE_SEGMENT|619,625|false|false|false|||NSTEMI
Finding|Finding|SIMPLE_SEGMENT|619,625|false|false|false|C3537184||NSTEMI
Event|Event|SIMPLE_SEGMENT|634,638|false|false|false|||cath
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|634,638|false|false|false|C0007430|Catheterization|cath
Event|Event|SIMPLE_SEGMENT|645,651|false|false|false|||showed
Finding|Finding|SIMPLE_SEGMENT|653,661|false|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Finding|Functional Concept|SIMPLE_SEGMENT|653,661|false|false|false|C0028778;C1947917|Obstruction;Occluded|occluded
Anatomy|Tissue|SIMPLE_SEGMENT|662,667|false|false|false|C0332835|Transplanted tissue|graft
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|662,667|false|false|false|C0181074;C1705210|Graft Dosage Form;Graft material|graft
Event|Event|SIMPLE_SEGMENT|662,667|false|false|false|||graft
Finding|Intellectual Product|SIMPLE_SEGMENT|662,667|false|false|false|C1546653|Graft - Specimen Source Codes|graft
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|662,667|false|false|false|C1961139;C3683798|Graft Procedures on the Head;Grafting procedure|graft
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|688,694|false|false|false|C1881507|Macromolecular Branch|branch
Event|Event|SIMPLE_SEGMENT|688,694|false|false|false|||branch
Finding|Finding|SIMPLE_SEGMENT|699,703|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|714,722|false|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|714,722|false|false|false|C1261287|Stenosis|stenosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|730,733|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|730,733|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|730,733|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Event|SIMPLE_SEGMENT|734,739|false|false|false|||stent
Event|Event|SIMPLE_SEGMENT|753,761|false|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|753,761|false|false|false|C1261287|Stenosis|stenosis
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|769,772|false|false|false|C2987138|Methylcytosine Dioxygenase TET1|LCx
Drug|Enzyme|SIMPLE_SEGMENT|769,772|false|false|false|C2987138|Methylcytosine Dioxygenase TET1|LCx
Event|Event|SIMPLE_SEGMENT|769,772|false|false|false|||LCx
Finding|Gene or Genome|SIMPLE_SEGMENT|769,772|false|false|false|C1428863;C2987137|TET1 gene;TET1 wt Allele|LCx
Event|Event|SIMPLE_SEGMENT|774,780|false|false|false|||origin
Finding|Classification|SIMPLE_SEGMENT|774,780|false|false|false|C0079946;C1550512|National origin;Participation Type - origin|origin
Finding|Intellectual Product|SIMPLE_SEGMENT|774,780|false|false|false|C0079946;C1550512|National origin;Participation Type - origin|origin
Event|Event|SIMPLE_SEGMENT|800,807|false|false|false|||managed
Event|Event|SIMPLE_SEGMENT|813,824|false|false|false|||uptitration
Drug|Organic Chemical|SIMPLE_SEGMENT|840,845|false|false|false|C0590690|Imdur|Imdur
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|840,845|false|false|false|C0590690|Imdur|Imdur
Event|Event|SIMPLE_SEGMENT|850,860|false|false|false|||initiation
Finding|Functional Concept|SIMPLE_SEGMENT|850,860|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Finding|Genetic Function|SIMPLE_SEGMENT|850,860|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Finding|Mental Process|SIMPLE_SEGMENT|850,860|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Drug|Organic Chemical|SIMPLE_SEGMENT|864,872|false|false|false|C0126174|losartan|losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|864,872|false|false|false|C0126174|losartan|losartan
Event|Event|SIMPLE_SEGMENT|864,872|false|false|false|||losartan
Finding|Idea or Concept|SIMPLE_SEGMENT|877,883|false|false|false|C1550462|Observation Interpretation - better|better
Drug|Organic Chemical|SIMPLE_SEGMENT|887,894|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|887,894|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|SIMPLE_SEGMENT|887,894|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Event|Event|SIMPLE_SEGMENT|887,894|false|false|false|||control
Finding|Conceptual Entity|SIMPLE_SEGMENT|887,894|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|SIMPLE_SEGMENT|887,894|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|SIMPLE_SEGMENT|887,894|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Intellectual Product|SIMPLE_SEGMENT|901,906|false|false|false|C4050225|Often - answer to question|often
Attribute|Clinical Attribute|SIMPLE_SEGMENT|911,917|false|false|false|C2926611||angina
Event|Event|SIMPLE_SEGMENT|911,917|false|false|false|||angina
Finding|Finding|SIMPLE_SEGMENT|911,917|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Finding|Sign or Symptom|SIMPLE_SEGMENT|911,917|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|911,925|false|false|false|C0002965;C0152172|Angina decubitus;Angina, Unstable|angina at rest
Finding|Functional Concept|SIMPLE_SEGMENT|918,925|false|false|false|C0443144|At rest (qualifier value)|at rest
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|921,925|false|false|false|C1742913|REST protein, human|rest
Drug|Biologically Active Substance|SIMPLE_SEGMENT|921,925|false|false|false|C1742913|REST protein, human|rest
Event|Event|SIMPLE_SEGMENT|921,925|false|false|false|||rest
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|921,925|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Gene or Genome|SIMPLE_SEGMENT|921,925|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Molecular Function|SIMPLE_SEGMENT|921,925|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|944,952|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|SIMPLE_SEGMENT|944,952|false|false|false|||baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|944,952|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Drug|Organic Chemical|SIMPLE_SEGMENT|960,973|false|false|false|C0017887|nitroglycerin|nitroglycerin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|960,973|false|false|false|C0017887|nitroglycerin|nitroglycerin
Event|Event|SIMPLE_SEGMENT|960,973|false|false|false|||nitroglycerin
Event|Event|SIMPLE_SEGMENT|1025,1034|false|false|false|||complains
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1047,1052|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|1047,1052|false|false|false|C0741025|Chest problem|chest
Finding|Sign or Symptom|SIMPLE_SEGMENT|1047,1058|false|false|false|C0008031|Chest Pain|chest pains
Event|Event|SIMPLE_SEGMENT|1053,1058|false|false|false|||pains
Finding|Sign or Symptom|SIMPLE_SEGMENT|1053,1058|false|false|false|C0030193|Pain|pains
Event|Event|SIMPLE_SEGMENT|1070,1079|false|false|false|||different
Finding|Intellectual Product|SIMPLE_SEGMENT|1089,1096|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|1089,1096|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1097,1103|false|false|false|C2926611||angina
Event|Event|SIMPLE_SEGMENT|1097,1103|false|false|false|||angina
Finding|Finding|SIMPLE_SEGMENT|1097,1103|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Finding|Sign or Symptom|SIMPLE_SEGMENT|1097,1103|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Finding|Finding|SIMPLE_SEGMENT|1111,1118|false|false|false|C3888388|Usually|usually
Event|Event|SIMPLE_SEGMENT|1119,1122|false|false|false|||ahs
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1123,1128|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|1123,1128|false|false|false|C0741025|Chest problem|chest
Event|Event|SIMPLE_SEGMENT|1130,1138|false|false|false|||pressire
Event|Event|SIMPLE_SEGMENT|1153,1158|false|false|false|||feels
Finding|Intellectual Product|SIMPLE_SEGMENT|1170,1176|false|false|false|C1546717||needle
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|1177,1183|false|false|false|C0033119|Puncture wound|pricks
Event|Event|SIMPLE_SEGMENT|1177,1183|false|false|false|||pricks
Finding|Finding|SIMPLE_SEGMENT|1177,1183|false|false|false|C0439821|Pricking sensation quality|pricks
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1186,1190|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|1186,1190|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1186,1190|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1186,1190|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|1205,1215|false|false|false|||persistent
Finding|Idea or Concept|SIMPLE_SEGMENT|1238,1249|false|true|false|C0750502|Significant|significant
Drug|Organic Chemical|SIMPLE_SEGMENT|1250,1256|true|true|false|C0723011|Relief brand of phenylephrine|relief
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1250,1256|true|true|false|C0723011|Relief brand of phenylephrine|relief
Event|Event|SIMPLE_SEGMENT|1250,1256|false|false|false|||relief
Finding|Finding|SIMPLE_SEGMENT|1250,1256|true|true|false|C0564405|Feeling relief|relief
Event|Event|SIMPLE_SEGMENT|1281,1286|false|false|false|||worse
Finding|Finding|SIMPLE_SEGMENT|1281,1286|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Idea or Concept|SIMPLE_SEGMENT|1281,1286|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1292,1296|false|false|false|C4318566|Deep Resection Margin|deep
Finding|Finding|SIMPLE_SEGMENT|1292,1306|false|false|false|C1321587;C1328799|Breathing abnormally deep;Deep breathing|deep breathing
Finding|Sign or Symptom|SIMPLE_SEGMENT|1292,1306|false|false|false|C1321587;C1328799|Breathing abnormally deep;Deep breathing|deep breathing
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1297,1306|false|false|false|C5885990||breathing
Event|Event|SIMPLE_SEGMENT|1297,1306|false|false|false|||breathing
Finding|Finding|SIMPLE_SEGMENT|1297,1306|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|SIMPLE_SEGMENT|1297,1306|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|SIMPLE_SEGMENT|1297,1306|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|SIMPLE_SEGMENT|1297,1306|false|false|false|C1160636|respiratory system process|breathing
Event|Event|SIMPLE_SEGMENT|1317,1325|false|false|false|||pressure
Finding|Finding|SIMPLE_SEGMENT|1317,1325|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|1317,1325|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|1317,1325|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|1317,1325|false|false|false|C0033095||pressure
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1329,1337|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Event|Event|SIMPLE_SEGMENT|1329,1337|false|false|false|||anterior
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1329,1343|false|false|false|C0230132|Anterior chest wall structure|anterior chest
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1338,1343|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|1338,1343|false|false|false|C0741025|Chest problem|chest
Event|Event|SIMPLE_SEGMENT|1349,1355|false|false|false|||states
Event|Event|SIMPLE_SEGMENT|1368,1372|false|false|false|||feel
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1383,1387|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|1383,1387|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1383,1387|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1383,1387|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|1407,1411|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1407,1411|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1419,1423|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|1419,1423|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1419,1423|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1419,1423|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|1436,1444|false|false|false|||remained
Event|Event|SIMPLE_SEGMENT|1446,1455|false|false|false|||continous
Event|Event|SIMPLE_SEGMENT|1464,1475|false|false|false|||accompanied
Event|Event|SIMPLE_SEGMENT|1484,1487|false|false|false|||SOB
Finding|Sign or Symptom|SIMPLE_SEGMENT|1484,1487|false|false|false|C0013404|Dyspnea|SOB
Event|Event|SIMPLE_SEGMENT|1492,1503|false|false|false|||diaphoresis
Finding|Finding|SIMPLE_SEGMENT|1492,1503|false|true|false|C0700590|Increased sweating|diaphoresis
Event|Event|SIMPLE_SEGMENT|1506,1520|false|false|false|||lighthededness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1522,1528|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|1522,1528|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1522,1528|false|false|false|C0027497|Nausea|nausea
Event|Event|SIMPLE_SEGMENT|1535,1547|false|false|false|||palpitations
Finding|Finding|SIMPLE_SEGMENT|1535,1547|false|false|false|C0030252|Palpitations|palpitations
Event|Event|SIMPLE_SEGMENT|1553,1559|false|false|false|||denies
Event|Event|SIMPLE_SEGMENT|1582,1589|false|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|1582,1589|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1582,1589|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Event|Event|SIMPLE_SEGMENT|1591,1600|false|false|false|||orthopnea
Finding|Finding|SIMPLE_SEGMENT|1591,1600|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1591,1600|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1602,1607|false|false|false|C0003086;C0003087;C4284979|Ankle;Ankle joint structure;Lower extremity>Ankle|ankle
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|1602,1607|false|false|false|C0003086;C0003087;C4284979|Ankle;Ankle joint structure;Lower extremity>Ankle|ankle
Finding|Pathologic Function|SIMPLE_SEGMENT|1602,1613|false|false|false|C0235439|Ankle edema (finding)|ankle edema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1608,1613|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|1608,1613|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|1608,1613|false|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|1615,1627|false|false|false|||palpitations
Finding|Finding|SIMPLE_SEGMENT|1615,1627|false|false|false|C0030252|Palpitations|palpitations
Event|Event|SIMPLE_SEGMENT|1629,1636|false|false|false|||syncope
Finding|Sign or Symptom|SIMPLE_SEGMENT|1629,1636|false|false|false|C0039070|Syncope|syncope
Event|Event|SIMPLE_SEGMENT|1641,1651|false|false|false|||presyncope
Finding|Sign or Symptom|SIMPLE_SEGMENT|1641,1651|false|false|false|C0700200|Presyncope|presyncope
Event|Event|SIMPLE_SEGMENT|1663,1667|false|false|false|||says
Event|Event|SIMPLE_SEGMENT|1686,1693|false|false|false|||feeling
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1699,1703|false|false|false|C0009443;C0024117|Chronic Obstructive Airway Disease;Common Cold|cold
Drug|Organic Chemical|SIMPLE_SEGMENT|1699,1703|false|false|false|C0719425|Cold brand of chlorpheniramine-phenylpropanolamine|cold
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1699,1703|false|false|false|C0719425|Cold brand of chlorpheniramine-phenylpropanolamine|cold
Event|Event|SIMPLE_SEGMENT|1699,1703|false|false|false|||cold
Finding|Organism Function|SIMPLE_SEGMENT|1699,1703|false|false|false|C0234192|Cold Sensation|cold
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|1699,1703|false|false|false|C0009264|Cold Temperature|cold
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1699,1703|false|false|false|C0010412|Cold Therapy|cold
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1725,1728|false|false|false|C0028723;C2985261|NUT Family Member 1, human;Nuts|nut
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1725,1728|false|false|false|C0028723;C2985261|NUT Family Member 1, human;Nuts|nut
Drug|Food|SIMPLE_SEGMENT|1725,1728|false|false|false|C0028723;C2985261|NUT Family Member 1, human;Nuts|nut
Event|Event|SIMPLE_SEGMENT|1725,1728|false|false|false|||nut
Finding|Gene or Genome|SIMPLE_SEGMENT|1725,1728|false|false|false|C1837033;C2985260|NUTM1 gene;NUTM1 wt Allele|nut
Event|Event|SIMPLE_SEGMENT|1729,1735|false|false|false|||denies
Event|Event|SIMPLE_SEGMENT|1740,1746|false|false|false|||fevers
Finding|Sign or Symptom|SIMPLE_SEGMENT|1740,1746|true|false|false|C0015967|Fever|fevers
Event|Event|SIMPLE_SEGMENT|1750,1756|false|false|false|||chills
Finding|Sign or Symptom|SIMPLE_SEGMENT|1750,1756|true|false|false|C0085593|Chills|chills
Finding|Intellectual Product|SIMPLE_SEGMENT|1768,1775|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|1768,1775|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Event|Event|SIMPLE_SEGMENT|1776,1786|false|false|false|||productive
Drug|Organic Chemical|SIMPLE_SEGMENT|1788,1793|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1788,1793|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|SIMPLE_SEGMENT|1788,1793|false|false|false|||cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|1788,1793|false|false|false|C0010200|Coughing|cough
Event|Event|SIMPLE_SEGMENT|1799,1805|false|false|false|||denies
Event|Event|SIMPLE_SEGMENT|1810,1812|false|false|false|||GI
Event|Event|SIMPLE_SEGMENT|1817,1827|false|false|false|||complaints
Finding|Finding|SIMPLE_SEGMENT|1817,1827|false|false|false|C5441521|Complaint (finding)|complaints
Finding|Body Substance|SIMPLE_SEGMENT|1843,1850|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1843,1850|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1843,1850|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|1867,1871|false|false|false|||work
Event|Event|SIMPLE_SEGMENT|1887,1891|false|false|false|||loss
Finding|Finding|SIMPLE_SEGMENT|1887,1891|false|false|false|C5890125|Loss (adaptation)|loss
Finding|Functional Concept|SIMPLE_SEGMENT|1897,1906|false|false|false|C1516691|Cognitive|cognitive
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1897,1917|false|false|false|C0338656|Impaired cognition|cognitive impairment
Event|Event|SIMPLE_SEGMENT|1907,1917|false|false|false|||impairment
Finding|Finding|SIMPLE_SEGMENT|1907,1917|false|false|false|C0221099;C0684336|Impaired;Impaired health|impairment
Finding|Functional Concept|SIMPLE_SEGMENT|1907,1917|false|false|false|C0221099;C0684336|Impaired;Impaired health|impairment
Event|Event|SIMPLE_SEGMENT|1972,1975|false|false|false|||EKG
Finding|Intellectual Product|SIMPLE_SEGMENT|1972,1975|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1972,1975|false|false|false|C1623258|Electrocardiography|EKG
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|1977,1982|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|1977,1982|false|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|SIMPLE_SEGMENT|1977,1982|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1977,1982|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Event|Event|SIMPLE_SEGMENT|1977,1982|false|false|false|||sinus
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1997,2008|false|false|false|C0011570|Mental Depression|depressions
Event|Event|SIMPLE_SEGMENT|1997,2008|false|false|false|||depressions
Event|Event|SIMPLE_SEGMENT|2009,2016|false|false|false|||similar
Finding|Finding|SIMPLE_SEGMENT|2030,2033|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|2030,2033|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Functional Concept|SIMPLE_SEGMENT|2035,2043|false|false|false|C0475224|Ischemic|ischemic
Event|Event|SIMPLE_SEGMENT|2044,2048|false|false|false|||chgs
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2050,2054|false|false|false|C0587081|Laboratory test finding|Labs
Event|Event|SIMPLE_SEGMENT|2055,2067|false|false|false|||unremarkable
Finding|Finding|SIMPLE_SEGMENT|2074,2077|false|false|false|C5848551|Neg - answer|neg
Event|Event|SIMPLE_SEGMENT|2082,2085|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2082,2085|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|SIMPLE_SEGMENT|2090,2095|false|false|false|||acute
Finding|Intellectual Product|SIMPLE_SEGMENT|2090,2095|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Finding|SIMPLE_SEGMENT|2101,2121|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|2106,2113|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|2106,2113|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|2106,2113|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|2106,2113|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2106,2113|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|2106,2121|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2114,2121|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2114,2121|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2114,2121|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2126,2133|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|SIMPLE_SEGMENT|2126,2133|false|false|false|C1314974|Cardiac attachment|CARDIAC
Finding|Finding|SIMPLE_SEGMENT|2126,2138|false|false|false|C3176821|CARD.RISK|CARDIAC RISK
Finding|Finding|SIMPLE_SEGMENT|2126,2146|false|false|false|C2024776|cardiac risk factors|CARDIAC RISK FACTORS
Event|Event|SIMPLE_SEGMENT|2134,2138|false|false|false|||RISK
Finding|Idea or Concept|SIMPLE_SEGMENT|2134,2138|false|false|false|C0035647|Risk|RISK
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2134,2146|false|false|false|C1830376||RISK FACTORS
Finding|Finding|SIMPLE_SEGMENT|2134,2146|false|false|false|C0035648;C0455624;C1553898|History of - risk factor;risk factors;risk factors - observation list|RISK FACTORS
Finding|Intellectual Product|SIMPLE_SEGMENT|2134,2146|false|false|false|C0035648;C0455624;C1553898|History of - risk factor;risk factors;risk factors - observation list|RISK FACTORS
Event|Event|SIMPLE_SEGMENT|2139,2146|false|false|false|||FACTORS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2151,2159|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|Diabetes
Event|Event|SIMPLE_SEGMENT|2151,2159|false|false|false|||Diabetes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2164,2176|false|false|false|C0242339|Dyslipidemias|Dyslipidemia
Event|Event|SIMPLE_SEGMENT|2164,2176|false|false|false|||Dyslipidemia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2181,2184|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|2181,2184|false|false|false|||HTN
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2190,2197|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|SIMPLE_SEGMENT|2190,2197|true|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Event|SIMPLE_SEGMENT|2198,2205|false|false|false|||HISTORY
Finding|Conceptual Entity|SIMPLE_SEGMENT|2198,2205|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|HISTORY
Finding|Finding|SIMPLE_SEGMENT|2198,2205|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|HISTORY
Finding|Functional Concept|SIMPLE_SEGMENT|2198,2205|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|HISTORY
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2210,2218|false|false|false|C0018787|Heart|Coronary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2210,2225|false|false|false|C0205042|Coronary artery|Coronary artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2210,2233|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|Coronary artery disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2219,2225|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|2219,2225|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2219,2233|false|false|false|C0852949|Arteriopathic disease|artery disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2226,2233|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|2226,2233|false|false|false|||disease
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2237,2246|false|false|false|C0012000|Diastole|Diastolic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2237,2271|false|false|false|C2183328|diastolic congestive heart failure|Diastolic congestive heart failure
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2247,2271|false|false|false|C0018802|Congestive heart failure|congestive heart failure
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2258,2263|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2258,2263|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|2258,2263|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2258,2271|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Event|Event|SIMPLE_SEGMENT|2264,2271|false|false|false|||failure
Finding|Functional Concept|SIMPLE_SEGMENT|2264,2271|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|SIMPLE_SEGMENT|2264,2271|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|SIMPLE_SEGMENT|2264,2271|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|SIMPLE_SEGMENT|2275,2279|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2275,2279|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Event|Event|SIMPLE_SEGMENT|2281,2285|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2281,2285|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2291,2322|false|false|false|C1449706|Coronary Artery Bypass, Off-Pump|Off pump coronary artery bypass
Finding|Molecular Function|SIMPLE_SEGMENT|2295,2299|false|false|false|C1150186|matrix metalloproteinase 7 activity|pump
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2300,2308|false|false|false|C0018787|Heart|coronary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2300,2315|false|false|false|C0205042|Coronary artery|coronary artery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2300,2322|false|false|false|C0010055|Coronary Artery Bypass Surgery|coronary artery bypass
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2300,2328|false|false|false|C0010055|Coronary Artery Bypass Surgery|coronary artery bypass graft
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2309,2315|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|2309,2315|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2309,2328|false|false|false|C5886769|Arterial bypass graft|artery bypass graft
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2316,2322|false|false|false|C0813207|Creation of shunt|bypass
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2316,2328|false|false|false|C0185098|Bypass graft|bypass graft
Anatomy|Tissue|SIMPLE_SEGMENT|2323,2328|false|false|false|C0332835|Transplanted tissue|graft
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2323,2328|false|false|false|C0181074;C1705210|Graft Dosage Form;Graft material|graft
Event|Event|SIMPLE_SEGMENT|2323,2328|false|false|false|||graft
Finding|Intellectual Product|SIMPLE_SEGMENT|2323,2328|false|false|false|C1546653|Graft - Specimen Source Codes|graft
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2323,2328|false|false|false|C1961139;C3683798|Graft Procedures on the Head;Grafting procedure|graft
Finding|Functional Concept|SIMPLE_SEGMENT|2333,2337|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2341,2364|false|false|false|C0226276|Structure of internal thoracic artery|internal mammary artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2350,2357|false|false|false|C0006141;C0929301|Breast;Mammary gland|mammary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2350,2364|false|false|false|C0024661|Mammary Arteries|mammary artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2358,2364|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|2358,2364|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Finding|Functional Concept|SIMPLE_SEGMENT|2368,2372|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2368,2399|false|false|false|C0226032;C1321506|Anterior descending branch of left coronary artery|left anterior descending artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2373,2381|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Finding|Functional Concept|SIMPLE_SEGMENT|2382,2392|false|false|false|C1547177|Sequencing - Descending|descending
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2393,2399|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|2393,2399|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2406,2420|false|false|false|C0036186;C0392907|Great saphenous vein structure;Saphenous Vein|saphenous vein
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2416,2420|false|false|false|C0042449|Veins|vein
Anatomy|Tissue|SIMPLE_SEGMENT|2421,2427|false|false|false|C0332835|Transplanted tissue|grafts
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2421,2427|false|false|false|C0181074|Graft material|grafts
Event|Event|SIMPLE_SEGMENT|2421,2427|false|false|false|||grafts
Finding|Finding|SIMPLE_SEGMENT|2452,2460|false|false|false|C1550517|Target Awareness - marginal|marginal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2461,2469|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Anatomy|Body System|SIMPLE_SEGMENT|2461,2469|false|false|false|C0003842;C0226004|Arterial system;Arteries|arteries
Procedure|Health Care Activity|SIMPLE_SEGMENT|2461,2469|false|false|false|C0397581|Procedure on artery|arteries
Finding|Functional Concept|SIMPLE_SEGMENT|2475,2487|false|false|false|C1522243|Percutaneous Route of Drug Administration|PERCUTANEOUS
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2475,2510|false|false|false|C1532338|Percutaneous Coronary Intervention|PERCUTANEOUS CORONARY INTERVENTIONS
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2488,2496|false|false|false|C0018787|Heart|CORONARY
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2497,2510|false|false|false|C2979881||INTERVENTIONS
Event|Event|SIMPLE_SEGMENT|2497,2510|false|false|false|||INTERVENTIONS
Procedure|Health Care Activity|SIMPLE_SEGMENT|2497,2510|false|false|false|C0886296;C1273869|Intervention regimes;Nursing interventions|INTERVENTIONS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2512,2515|false|false|false|C0006430|Burning Mouth Syndrome|BMS
Event|Event|SIMPLE_SEGMENT|2512,2515|false|false|false|||BMS
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2519,2527|false|false|false|C4489236|Proximal Resection Margin|proximal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2528,2531|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2528,2531|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|SIMPLE_SEGMENT|2528,2531|false|false|false|||LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|2528,2531|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2539,2542|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2539,2542|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2539,2542|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|SIMPLE_SEGMENT|2539,2542|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|SIMPLE_SEGMENT|2539,2542|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2539,2542|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Event|Event|SIMPLE_SEGMENT|2539,2542|false|false|false|||DES
Finding|Gene or Genome|SIMPLE_SEGMENT|2539,2542|false|false|false|C1413980|DES gene|DES
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2550,2553|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2550,2553|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|SIMPLE_SEGMENT|2550,2553|false|false|false|||LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|2550,2553|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2559,2562|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2559,2562|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2559,2562|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|SIMPLE_SEGMENT|2559,2562|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|SIMPLE_SEGMENT|2559,2562|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2559,2562|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Event|Event|SIMPLE_SEGMENT|2559,2562|false|false|false|||DES
Finding|Gene or Genome|SIMPLE_SEGMENT|2559,2562|false|false|false|C1413980|DES gene|DES
Event|Event|SIMPLE_SEGMENT|2566,2570|false|false|false|||edge
Finding|Conceptual Entity|SIMPLE_SEGMENT|2566,2570|false|false|false|C2697523|Graph Edge|edge
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2582,2585|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2582,2585|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|2582,2585|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2586,2589|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2586,2589|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2586,2589|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|SIMPLE_SEGMENT|2586,2589|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|SIMPLE_SEGMENT|2586,2589|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2586,2589|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Event|Event|SIMPLE_SEGMENT|2586,2589|false|false|false|||DES
Finding|Gene or Genome|SIMPLE_SEGMENT|2586,2589|false|false|false|C1413980|DES gene|DES
Event|Event|SIMPLE_SEGMENT|2596,2604|false|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|2596,2604|false|false|false|C1261287|Stenosis|stenosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2605,2611|false|false|false|C4522154|Distal Resection Margin|distal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2626,2629|false|false|false|C4551552|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|DES
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2626,2629|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2626,2629|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Hormone|SIMPLE_SEGMENT|2626,2629|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Organic Chemical|SIMPLE_SEGMENT|2626,2629|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2626,2629|false|false|false|C0011702;C0012203;C5441700|DES protein, human;Desmosine;diethylstilbestrol|DES
Event|Event|SIMPLE_SEGMENT|2626,2629|false|false|false|||DES
Finding|Gene or Genome|SIMPLE_SEGMENT|2626,2629|false|false|false|C1413980|DES gene|DES
Finding|Individual Behavior|SIMPLE_SEGMENT|2645,2651|false|false|false|C0562458|Pacing up and down|PACING
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2652,2655|false|false|false|C0020725;C0021122|Disruptive, Impulse Control, and Conduct Disorders;Type II Mucolipidosis|ICD
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2652,2655|false|false|false|C0020725;C0021122|Disruptive, Impulse Control, and Conduct Disorders;Type II Mucolipidosis|ICD
Event|Event|SIMPLE_SEGMENT|2652,2655|false|false|false|||ICD
Finding|Gene or Genome|SIMPLE_SEGMENT|2652,2655|false|false|false|C0870733;C5891008|GNPTAB wt Allele;International Classification of Diseases|ICD
Finding|Intellectual Product|SIMPLE_SEGMENT|2652,2655|false|false|false|C0870733;C5891008|GNPTAB wt Allele;International Classification of Diseases|ICD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2652,2655|false|false|false|C5575277|Icd Regimen|ICD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2663,2677|false|false|false|C0028756|Morbid obesity|Morbid obesity
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2670,2677|false|false|false|C0028754|Obesity|obesity
Event|Event|SIMPLE_SEGMENT|2670,2677|false|false|false|||obesity
Finding|Finding|SIMPLE_SEGMENT|2670,2677|false|false|false|C4759928|BODY MASS INDEX QUANTITATIVE TRAIT LOCUS 20|obesity
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2681,2685|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2681,2685|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|SIMPLE_SEGMENT|2681,2685|false|false|false|||COPD
Finding|Gene or Genome|SIMPLE_SEGMENT|2681,2685|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2688,2692|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|SIMPLE_SEGMENT|2688,2692|false|false|false|||GERD
Finding|Functional Concept|SIMPLE_SEGMENT|2695,2700|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2695,2713|false|false|false|C0828608|Right tendinous cuff|Right rotator cuff
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2701,2713|false|false|false|C0085515|Rotator Cuff|rotator cuff
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|2701,2720|false|false|false|C0851122|Rotator Cuff Injuries|rotator cuff injury
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2709,2713|false|false|false|C1550244|Cuff - body part|cuff
Finding|Pathologic Function|SIMPLE_SEGMENT|2709,2713|false|false|false|C3668885|Cuffing (morphologic abnormality)|cuff
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|2714,2720|false|false|false|C3263722;C3263723|Traumatic AND/OR non-traumatic injury;Traumatic injury|injury
Event|Event|SIMPLE_SEGMENT|2714,2720|false|false|false|||injury
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2721,2729|false|false|false|C0006444|Bursitis|bursitis
Event|Event|SIMPLE_SEGMENT|2721,2729|false|false|false|||bursitis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2732,2741|false|false|false|C0149931|Migraine Disorders|Migraines
Event|Event|SIMPLE_SEGMENT|2732,2741|false|false|false|||Migraines
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2744,2754|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|Depression
Event|Event|SIMPLE_SEGMENT|2744,2754|false|false|false|||Depression
Finding|Functional Concept|SIMPLE_SEGMENT|2744,2754|false|false|false|C0460137;C1579931|Depression - motion|Depression
Finding|Sign or Symptom|SIMPLE_SEGMENT|2744,2754|false|false|false|C0460137;C1579931|Depression - motion|Depression
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2757,2760|false|false|false|C0029408|Degenerative polyarthritis|DJD
Event|Event|SIMPLE_SEGMENT|2757,2760|false|false|false|||DJD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2763,2774|false|false|false|C0019112|Hemorrhoids|Hemorrhoids
Event|Event|SIMPLE_SEGMENT|2763,2774|false|false|false|||Hemorrhoids
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2777,2784|false|false|false|C0035854|Rosacea|Rosacea
Event|Event|SIMPLE_SEGMENT|2777,2784|false|false|false|||Rosacea
Finding|Functional Concept|SIMPLE_SEGMENT|2790,2796|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|2790,2804|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|2797,2804|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2797,2804|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2797,2804|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2797,2804|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|2810,2816|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2810,2816|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|2810,2816|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|2810,2816|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|2810,2824|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|2817,2824|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2817,2824|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2817,2824|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2817,2824|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Event|Event|SIMPLE_SEGMENT|2865,2869|false|false|false|||know
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2870,2880|false|true|false|C3812393|ErbB Receptors|her family
Drug|Enzyme|SIMPLE_SEGMENT|2870,2880|false|true|false|C3812393|ErbB Receptors|her family
Finding|Receptor|SIMPLE_SEGMENT|2870,2880|false|true|false|C3812393|ErbB Receptors|her family
Event|Event|SIMPLE_SEGMENT|2874,2880|false|false|false|||family
Finding|Classification|SIMPLE_SEGMENT|2874,2880|true|true|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2874,2880|true|true|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|2874,2880|true|true|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|2874,2880|true|true|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Event|Event|SIMPLE_SEGMENT|2887,2895|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|2887,2895|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|2887,2895|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2887,2895|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|2887,2900|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2887,2900|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|2896,2900|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|2896,2900|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2896,2900|false|false|false|C0582103|Medical Examination|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2902,2911|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|SIMPLE_SEGMENT|2912,2916|false|false|false|||EXAM
Finding|Functional Concept|SIMPLE_SEGMENT|2912,2916|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|2912,2916|false|false|false|C0582103|Medical Examination|EXAM
Event|Event|SIMPLE_SEGMENT|2922,2923|false|false|false|||T
Event|Event|SIMPLE_SEGMENT|2929,2931|false|false|false|||BP
Event|Event|SIMPLE_SEGMENT|2954,2957|false|false|false|||sat
Event|Event|SIMPLE_SEGMENT|2965,2972|false|false|false|||GENERAL
Finding|Classification|SIMPLE_SEGMENT|2965,2972|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|2965,2972|false|false|false|C3812897|General medical service|GENERAL
Finding|Finding|SIMPLE_SEGMENT|2974,2982|false|false|false|C1961028|Oriented to place|Oriented
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2987,2991|false|false|false|C2713234||Mood
Event|Event|SIMPLE_SEGMENT|2987,2991|false|false|false|||Mood
Finding|Conceptual Entity|SIMPLE_SEGMENT|2987,2991|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Finding|Finding|SIMPLE_SEGMENT|2987,2991|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Finding|Mental Process|SIMPLE_SEGMENT|2987,2991|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Event|Event|SIMPLE_SEGMENT|2993,2999|false|false|false|||affect
Event|Event|SIMPLE_SEGMENT|3000,3011|false|false|false|||appropriate
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3015,3020|false|false|false|C1512338|HEENT|HEENT
Event|Event|SIMPLE_SEGMENT|3022,3026|false|false|false|||NCAT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3028,3034|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3028,3034|false|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|SIMPLE_SEGMENT|3028,3034|false|false|false|||Sclera
Procedure|Health Care Activity|SIMPLE_SEGMENT|3028,3034|false|false|false|C2228481|examination of sclera|Sclera
Event|Event|SIMPLE_SEGMENT|3035,3044|false|false|false|||anicteric
Finding|Finding|SIMPLE_SEGMENT|3035,3044|false|false|false|C0205180|Anicteric|anicteric
Event|Event|SIMPLE_SEGMENT|3046,3051|false|false|false|||PERRL
Finding|Finding|SIMPLE_SEGMENT|3046,3051|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Event|Event|SIMPLE_SEGMENT|3053,3057|false|false|false|||EOMI
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3059,3070|false|false|false|C0009758;C0229274|Structure of palpebral conjunctiva;conjunctiva|Conjunctiva
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3059,3070|false|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|Conjunctiva
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3059,3070|false|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|Conjunctiva
Event|Event|SIMPLE_SEGMENT|3059,3070|false|false|false|||Conjunctiva
Finding|Body Substance|SIMPLE_SEGMENT|3059,3070|false|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|Conjunctiva
Finding|Intellectual Product|SIMPLE_SEGMENT|3059,3070|false|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|Conjunctiva
Procedure|Health Care Activity|SIMPLE_SEGMENT|3059,3070|false|false|false|C0872390;C2228431|Procedure on conjunctiva;examination of conjunctiva|Conjunctiva
Event|Event|SIMPLE_SEGMENT|3086,3092|false|false|false|||pallor
Finding|Finding|SIMPLE_SEGMENT|3086,3092|true|false|false|C0241137|Pallor of skin|pallor
Event|Event|SIMPLE_SEGMENT|3096,3104|false|false|false|||cyanosis
Finding|Sign or Symptom|SIMPLE_SEGMENT|3096,3104|true|false|false|C0010520|Cyanosis|cyanosis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|3112,3116|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3112,3116|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|3112,3116|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|3112,3116|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3112,3123|false|false|false|C0026639|Oral mucous membrane structure|oral mucosa
Anatomy|Tissue|SIMPLE_SEGMENT|3117,3123|false|false|false|C0026724|Mucous Membrane|mucosa
Finding|Intellectual Product|SIMPLE_SEGMENT|3117,3123|false|false|false|C1561514||mucosa
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3128,3139|true|false|false|C0155210;C0302314|Eyelid Xanthoma;Xanthoma|xanthelasma
Event|Event|SIMPLE_SEGMENT|3128,3139|false|false|false|||xanthelasma
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3144,3148|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|SIMPLE_SEGMENT|3144,3148|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|SIMPLE_SEGMENT|3144,3148|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|SIMPLE_SEGMENT|3150,3156|false|false|false|||Supple
Finding|Functional Concept|SIMPLE_SEGMENT|3150,3156|false|false|false|C0332254|Supple|Supple
Event|Event|SIMPLE_SEGMENT|3162,3165|false|false|false|||JVP
Finding|Finding|SIMPLE_SEGMENT|3162,3165|false|false|false|C0428897|Jugular venous pressure|JVP
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3177,3182|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|SIMPLE_SEGMENT|3177,3182|false|false|false|C0741025|Chest problem|Chest
Finding|Idea or Concept|SIMPLE_SEGMENT|3184,3195|false|false|false|C0750502|Significant|significant
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3204,3207|false|false|false|C0034155;C1268935|Congenital Thrombotic Thrombocytopenic Purpura;Purpura, Thrombotic Thrombocytopenic|TTP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3204,3207|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3204,3207|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Drug|Organic Chemical|SIMPLE_SEGMENT|3204,3207|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Drug|Vitamin|SIMPLE_SEGMENT|3204,3207|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Event|Event|SIMPLE_SEGMENT|3204,3207|false|false|false|||TTP
Finding|Gene or Genome|SIMPLE_SEGMENT|3204,3207|false|false|false|C1413036;C1421571;C3539814|ADAMTS13 gene;ZFP36 gene;ZFP36 wt Allele|TTP
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3213,3221|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3213,3227|false|false|false|C0230132|Anterior chest wall structure|anterior chest
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3213,3232|false|false|false|C0230132;C1305714|Anterior chest wall structure|anterior chest wall
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3213,3232|false|false|false|C0230132;C1305714|Anterior chest wall structure|anterior chest wall
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3222,3227|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|3222,3227|false|false|false|C0741025|Chest problem|chest
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3222,3232|false|false|false|C0205076;C4266615|Chest wall structure;Chest>Chest wall|chest wall
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3222,3232|false|false|false|C0205076;C4266615|Chest wall structure;Chest>Chest wall|chest wall
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3236,3243|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|SIMPLE_SEGMENT|3236,3243|false|false|false|C1314974|Cardiac attachment|CARDIAC
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3249,3253|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Event|Event|SIMPLE_SEGMENT|3254,3257|false|false|false|||RRR
Event|Event|SIMPLE_SEGMENT|3265,3266|false|false|false|||g
Event|Event|SIMPLE_SEGMENT|3271,3278|false|false|false|||thrills
Finding|Finding|SIMPLE_SEGMENT|3271,3278|true|false|false|C0232269|Cardiac thrill (finding)|thrills
Event|Event|SIMPLE_SEGMENT|3280,3285|false|false|false|||lifts
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3303,3308|false|false|false|C0024109|Lung|LUNGS
Finding|Functional Concept|SIMPLE_SEGMENT|3317,3321|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Event|Event|SIMPLE_SEGMENT|3330,3338|false|false|false|||crackles
Finding|Finding|SIMPLE_SEGMENT|3330,3338|false|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Event|Event|SIMPLE_SEGMENT|3352,3362|false|false|false|||consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|3352,3362|false|true|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|3352,3367|false|true|false|C0332290|Consistent with|consistent with
Anatomy|Tissue|SIMPLE_SEGMENT|3369,3376|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3369,3376|false|false|false|C0032226|Pleural Diseases|pleural
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3377,3384|false|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3377,3384|false|false|false|C1951340|Process Pharmacologic Substance|process
Event|Event|SIMPLE_SEGMENT|3377,3384|false|false|false|||process
Finding|Functional Concept|SIMPLE_SEGMENT|3377,3384|false|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|3377,3384|false|false|false|C1522240|Process|process
Event|Event|SIMPLE_SEGMENT|3385,3389|false|false|false|||seen
Event|Event|SIMPLE_SEGMENT|3393,3396|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3393,3396|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Idea or Concept|SIMPLE_SEGMENT|3408,3412|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3413,3416|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3413,3416|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|SIMPLE_SEGMENT|3413,3416|false|false|false|C0001861;C3536832|Air (substance);air|air
Finding|Finding|SIMPLE_SEGMENT|3413,3416|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|SIMPLE_SEGMENT|3413,3416|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|SIMPLE_SEGMENT|3413,3416|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3413,3425|false|false|false|C0001868|Air Movements|air movement
Event|Event|SIMPLE_SEGMENT|3417,3425|false|false|false|||movement
Finding|Organism Function|SIMPLE_SEGMENT|3417,3425|false|false|false|C0026649|Movement|movement
Event|Event|SIMPLE_SEGMENT|3435,3442|false|false|false|||wheezes
Finding|Sign or Symptom|SIMPLE_SEGMENT|3435,3442|false|false|false|C0043144|Wheezing|wheezes
Event|Event|SIMPLE_SEGMENT|3446,3453|false|false|false|||rhonchi
Finding|Finding|SIMPLE_SEGMENT|3446,3453|false|false|false|C0035508|Rhonchi|rhonchi
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3457,3464|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3457,3464|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|SIMPLE_SEGMENT|3457,3464|false|false|false|||ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|3457,3464|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3466,3470|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|SIMPLE_SEGMENT|3466,3470|false|false|false|||Soft
Event|Event|SIMPLE_SEGMENT|3472,3476|false|false|false|||NTND
Event|Event|SIMPLE_SEGMENT|3481,3484|false|false|false|||HSM
Finding|Gene or Genome|SIMPLE_SEGMENT|3481,3484|true|false|false|C1537594|LRRC4B gene|HSM
Event|Event|SIMPLE_SEGMENT|3488,3498|false|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|3488,3498|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|3488,3498|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3500,3503|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|Abd
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|3500,3503|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|Abd
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3504,3509|false|false|false|C0003483;C4037978|Aorta;Chest+Abdomen>Aorta|aorta
Procedure|Health Care Activity|SIMPLE_SEGMENT|3504,3509|false|false|false|C0869784|Procedure on aorta|aorta
Event|Event|SIMPLE_SEGMENT|3515,3523|false|false|false|||enlarged
Event|Event|SIMPLE_SEGMENT|3527,3536|false|false|false|||palpation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3527,3536|false|false|false|C0030247|Palpation|palpation
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3541,3550|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|SIMPLE_SEGMENT|3541,3557|true|false|false|C0221755|Abdominal bruit|abdominal bruits
Event|Event|SIMPLE_SEGMENT|3551,3557|false|false|false|||bruits
Finding|Finding|SIMPLE_SEGMENT|3551,3557|true|false|false|C0006318|Bruit|bruits
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3561,3572|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3587,3594|false|false|false|C0015811|Femur|femoral
Event|Event|SIMPLE_SEGMENT|3595,3601|false|false|false|||bruits
Finding|Finding|SIMPLE_SEGMENT|3595,3601|true|false|false|C0006318|Bruit|bruits
Anatomy|Body System|SIMPLE_SEGMENT|3605,3609|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3605,3609|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3605,3609|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|SIMPLE_SEGMENT|3605,3609|false|false|false|||SKIN
Finding|Body Substance|SIMPLE_SEGMENT|3605,3609|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|SIMPLE_SEGMENT|3605,3609|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Pathologic Function|SIMPLE_SEGMENT|3614,3620|false|false|false|C0333138|Stasis|stasis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3614,3631|true|false|false|C0011620|Stasis dermatitis|stasis dermatitis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3621,3631|true|false|false|C0011603|Dermatitis|dermatitis
Event|Event|SIMPLE_SEGMENT|3621,3631|false|false|false|||dermatitis
Event|Event|SIMPLE_SEGMENT|3633,3639|false|false|false|||ulcers
Finding|Pathologic Function|SIMPLE_SEGMENT|3633,3639|true|false|false|C0041582|Ulcer|ulcers
Event|Event|SIMPLE_SEGMENT|3641,3646|false|false|false|||scars
Finding|Finding|SIMPLE_SEGMENT|3641,3646|true|false|false|C0241158;C2004491|Cicatrix;Scar Tissue|scars
Finding|Pathologic Function|SIMPLE_SEGMENT|3641,3646|true|false|false|C0241158;C2004491|Cicatrix;Scar Tissue|scars
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3651,3660|true|false|false|C0302314|Xanthoma|xanthomas
Event|Event|SIMPLE_SEGMENT|3651,3660|false|false|false|||xanthomas
Drug|Food|SIMPLE_SEGMENT|3664,3670|false|false|false|C5890763||PULSES
Event|Event|SIMPLE_SEGMENT|3664,3670|false|false|false|||PULSES
Finding|Physiologic Function|SIMPLE_SEGMENT|3664,3670|false|false|false|C0391850|Physiologic pulse|PULSES
Procedure|Health Care Activity|SIMPLE_SEGMENT|3664,3670|false|false|false|C0034107|Pulse taking|PULSES
Finding|Body Substance|SIMPLE_SEGMENT|3722,3731|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|3722,3731|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|3722,3731|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|3722,3731|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|SIMPLE_SEGMENT|3732,3736|false|false|false|||EXAM
Finding|Functional Concept|SIMPLE_SEGMENT|3732,3736|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|3732,3736|false|false|false|C0582103|Medical Examination|EXAM
Event|Event|SIMPLE_SEGMENT|3742,3743|false|false|false|||T
Event|Event|SIMPLE_SEGMENT|3749,3751|false|false|false|||BP
Event|Event|SIMPLE_SEGMENT|3770,3772|false|false|false|||RR
Event|Event|SIMPLE_SEGMENT|3779,3782|false|false|false|||sat
Event|Event|SIMPLE_SEGMENT|3790,3797|false|false|false|||GENERAL
Finding|Classification|SIMPLE_SEGMENT|3790,3797|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|3790,3797|false|false|false|C3812897|General medical service|GENERAL
Finding|Finding|SIMPLE_SEGMENT|3799,3807|false|false|false|C1961028|Oriented to place|Oriented
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3812,3816|false|false|false|C2713234||Mood
Finding|Conceptual Entity|SIMPLE_SEGMENT|3812,3816|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Finding|Finding|SIMPLE_SEGMENT|3812,3816|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Finding|Mental Process|SIMPLE_SEGMENT|3812,3816|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Event|Event|SIMPLE_SEGMENT|3817,3828|false|false|false|||appropriate
Finding|Finding|SIMPLE_SEGMENT|3834,3845|false|false|false|C0233471|Flat affect|flat affect
Event|Event|SIMPLE_SEGMENT|3839,3845|false|false|false|||affect
Finding|Mental Process|SIMPLE_SEGMENT|3839,3845|false|false|false|C0001721|Affect (mental function)|affect
Procedure|Health Care Activity|SIMPLE_SEGMENT|3839,3845|false|false|false|C2237113|assessment of affect|affect
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3848,3851|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3848,3851|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3848,3851|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|3848,3851|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3848,3851|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|3848,3851|false|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|3848,3851|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3854,3859|false|false|false|C1512338|HEENT|HEENT
Event|Event|SIMPLE_SEGMENT|3861,3865|false|false|false|||NCAT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3867,3873|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3867,3873|false|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|SIMPLE_SEGMENT|3867,3873|false|false|false|||Sclera
Procedure|Health Care Activity|SIMPLE_SEGMENT|3867,3873|false|false|false|C2228481|examination of sclera|Sclera
Event|Event|SIMPLE_SEGMENT|3874,3883|false|false|false|||anicteric
Finding|Finding|SIMPLE_SEGMENT|3874,3883|false|false|false|C0205180|Anicteric|anicteric
Event|Event|SIMPLE_SEGMENT|3885,3890|false|false|false|||PERRL
Finding|Finding|SIMPLE_SEGMENT|3885,3890|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Event|Event|SIMPLE_SEGMENT|3892,3896|false|false|false|||EOMI
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3898,3909|false|false|false|C0009758;C0229274|Structure of palpebral conjunctiva;conjunctiva|Conjunctiva
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3898,3909|false|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|Conjunctiva
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3898,3909|false|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|Conjunctiva
Event|Event|SIMPLE_SEGMENT|3898,3909|false|false|false|||Conjunctiva
Finding|Body Substance|SIMPLE_SEGMENT|3898,3909|false|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|Conjunctiva
Finding|Intellectual Product|SIMPLE_SEGMENT|3898,3909|false|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|Conjunctiva
Procedure|Health Care Activity|SIMPLE_SEGMENT|3898,3909|false|false|false|C0872390;C2228431|Procedure on conjunctiva;examination of conjunctiva|Conjunctiva
Event|Event|SIMPLE_SEGMENT|3925,3931|false|false|false|||pallor
Finding|Finding|SIMPLE_SEGMENT|3925,3931|true|false|false|C0241137|Pallor of skin|pallor
Event|Event|SIMPLE_SEGMENT|3935,3943|false|false|false|||cyanosis
Finding|Sign or Symptom|SIMPLE_SEGMENT|3935,3943|true|false|false|C0010520|Cyanosis|cyanosis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|3951,3955|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3951,3955|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|3951,3955|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|3951,3955|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3951,3962|false|false|false|C0026639|Oral mucous membrane structure|oral mucosa
Anatomy|Tissue|SIMPLE_SEGMENT|3956,3962|false|false|false|C0026724|Mucous Membrane|mucosa
Finding|Intellectual Product|SIMPLE_SEGMENT|3956,3962|false|false|false|C1561514||mucosa
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3967,3978|true|false|false|C0155210;C0302314|Eyelid Xanthoma;Xanthoma|xanthelasma
Event|Event|SIMPLE_SEGMENT|3967,3978|false|false|false|||xanthelasma
Finding|Functional Concept|SIMPLE_SEGMENT|3982,3986|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3982,3993|false|false|false|C0229124|Structure of cornea of left eye|Left cornea
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3987,3993|false|false|false|C0010031|Cornea|cornea
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3987,3993|false|false|false|C0010034;C0153629;C0154026|Benign neoplasm of cornea;Corneal Diseases;Malignant neoplasm of cornea|cornea
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3987,3993|false|false|false|C0010034;C0153629;C0154026|Benign neoplasm of cornea;Corneal Diseases;Malignant neoplasm of cornea|cornea
Event|Event|SIMPLE_SEGMENT|3987,3993|false|false|false|||cornea
Finding|Body Substance|SIMPLE_SEGMENT|3987,3993|false|false|false|C1550625|SpecimenType - Cornea|cornea
Finding|Finding|SIMPLE_SEGMENT|3999,4003|false|false|false|C0241158;C1419736;C2004491|Cicatrix;RPS4X gene;Scar Tissue|scar
Finding|Gene or Genome|SIMPLE_SEGMENT|3999,4003|false|false|false|C0241158;C1419736;C2004491|Cicatrix;RPS4X gene;Scar Tissue|scar
Finding|Pathologic Function|SIMPLE_SEGMENT|3999,4003|false|false|false|C0241158;C1419736;C2004491|Cicatrix;RPS4X gene;Scar Tissue|scar
Finding|Finding|SIMPLE_SEGMENT|3999,4010|false|false|false|C0241158;C2004491|Cicatrix;Scar Tissue|scar tissue
Finding|Pathologic Function|SIMPLE_SEGMENT|3999,4010|false|false|false|C0241158;C2004491|Cicatrix;Scar Tissue|scar tissue
Anatomy|Tissue|SIMPLE_SEGMENT|4004,4010|false|false|false|C0040300|Body tissue|tissue
Finding|Intellectual Product|SIMPLE_SEGMENT|4004,4010|false|false|false|C1547928|Tissue Specimen Code|tissue
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4026,4030|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|SIMPLE_SEGMENT|4026,4030|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|SIMPLE_SEGMENT|4026,4030|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|SIMPLE_SEGMENT|4032,4038|false|false|false|||Supple
Finding|Functional Concept|SIMPLE_SEGMENT|4032,4038|false|false|false|C0332254|Supple|Supple
Event|Event|SIMPLE_SEGMENT|4049,4052|false|false|false|||JVP
Finding|Finding|SIMPLE_SEGMENT|4049,4052|false|false|false|C0428897|Jugular venous pressure|JVP
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4058,4069|true|false|false|C0018021|Goiter|thyromegaly
Event|Event|SIMPLE_SEGMENT|4058,4069|false|false|false|||thyromegaly
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4071,4076|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|CHEST
Finding|Finding|SIMPLE_SEGMENT|4071,4076|false|false|false|C0741025|Chest problem|CHEST
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4078,4081|false|false|false|C0034155;C1268935|Congenital Thrombotic Thrombocytopenic Purpura;Purpura, Thrombotic Thrombocytopenic|TTP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4078,4081|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4078,4081|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Drug|Organic Chemical|SIMPLE_SEGMENT|4078,4081|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Drug|Vitamin|SIMPLE_SEGMENT|4078,4081|false|false|false|C1506603;C4723973|ZFP36 protein, human;thiamine triphosphorate|TTP
Event|Event|SIMPLE_SEGMENT|4078,4081|false|false|false|||TTP
Finding|Gene or Genome|SIMPLE_SEGMENT|4078,4081|false|false|false|C1413036;C1421571;C3539814|ADAMTS13 gene;ZFP36 gene;ZFP36 wt Allele|TTP
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4087,4094|false|false|false|C0038293|Sternum|sternum
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4095,4102|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|SIMPLE_SEGMENT|4095,4102|false|false|false|C1314974|Cardiac attachment|CARDIAC
Finding|Pathologic Function|SIMPLE_SEGMENT|4104,4111|false|false|false|C5441917|Distant Metastasis|Distant
Finding|Finding|SIMPLE_SEGMENT|4104,4124|false|false|false|C2198873|distant heart sounds|Distant heart sounds
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4112,4117|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4112,4117|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|4112,4117|false|false|false|C0795691|HEART PROBLEM|heart
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4112,4124|false|false|false|C4050434||heart sounds
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4112,4124|false|false|false|C0018820|Heart Sounds|heart sounds
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4112,4124|false|false|false|C2230284|auscultation of heart sounds|heart sounds
Event|Event|SIMPLE_SEGMENT|4118,4124|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|4118,4124|false|false|false|C0037709||sounds
Event|Event|SIMPLE_SEGMENT|4133,4134|false|false|false|||g
Event|Event|SIMPLE_SEGMENT|4139,4146|false|false|false|||thrills
Finding|Finding|SIMPLE_SEGMENT|4139,4146|true|false|false|C0232269|Cardiac thrill (finding)|thrills
Event|Event|SIMPLE_SEGMENT|4148,4153|false|false|false|||lifts
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4171,4176|false|false|false|C0024109|Lung|LUNGS
Drug|Organic Chemical|SIMPLE_SEGMENT|4178,4182|false|false|false|C0951233|cetrimonium bromide|CTAB
Event|Event|SIMPLE_SEGMENT|4178,4182|false|false|false|||CTAB
Event|Event|SIMPLE_SEGMENT|4186,4194|false|false|false|||wheezing
Finding|Sign or Symptom|SIMPLE_SEGMENT|4186,4194|true|false|false|C0043144|Wheezing|wheezing
Event|Event|SIMPLE_SEGMENT|4196,4201|false|false|false|||rales
Finding|Finding|SIMPLE_SEGMENT|4196,4201|true|false|false|C0034642;C0240859|Basilar Rales;Rales|rales
Event|Event|SIMPLE_SEGMENT|4203,4210|false|false|false|||rhonchi
Finding|Finding|SIMPLE_SEGMENT|4203,4210|true|false|false|C0035508|Rhonchi|rhonchi
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4213,4220|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4213,4220|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|SIMPLE_SEGMENT|4213,4220|false|false|false|||ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|4213,4220|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4222,4227|false|false|false|C0028754|Obesity|Obese
Event|Event|SIMPLE_SEGMENT|4222,4227|false|false|false|||Obese
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4229,4233|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|SIMPLE_SEGMENT|4229,4233|false|false|false|||soft
Event|Event|SIMPLE_SEGMENT|4235,4239|false|false|false|||NTND
Event|Event|SIMPLE_SEGMENT|4244,4247|false|false|false|||HSM
Finding|Gene or Genome|SIMPLE_SEGMENT|4244,4247|true|false|false|C1537594|LRRC4B gene|HSM
Event|Event|SIMPLE_SEGMENT|4251,4261|false|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|4251,4261|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|4251,4261|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4263,4266|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|Abd
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|4263,4266|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|Abd
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4267,4272|false|false|false|C0003483;C4037978|Aorta;Chest+Abdomen>Aorta|aorta
Procedure|Health Care Activity|SIMPLE_SEGMENT|4267,4272|false|false|false|C0869784|Procedure on aorta|aorta
Event|Event|SIMPLE_SEGMENT|4278,4286|false|false|false|||enlarged
Event|Event|SIMPLE_SEGMENT|4290,4299|false|false|false|||palpation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4290,4299|false|false|false|C0030247|Palpation|palpation
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4304,4313|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|SIMPLE_SEGMENT|4304,4320|true|false|false|C0221755|Abdominal bruit|abdominal bruits
Event|Event|SIMPLE_SEGMENT|4314,4320|false|false|false|||bruits
Finding|Finding|SIMPLE_SEGMENT|4314,4320|true|false|false|C0006318|Bruit|bruits
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4324,4335|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4350,4357|false|false|false|C0015811|Femur|femoral
Event|Event|SIMPLE_SEGMENT|4358,4364|false|false|false|||bruits
Finding|Finding|SIMPLE_SEGMENT|4358,4364|true|false|false|C0006318|Bruit|bruits
Anatomy|Body System|SIMPLE_SEGMENT|4368,4372|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4368,4372|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4368,4372|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|SIMPLE_SEGMENT|4368,4372|false|false|false|||SKIN
Finding|Body Substance|SIMPLE_SEGMENT|4368,4372|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|SIMPLE_SEGMENT|4368,4372|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Pathologic Function|SIMPLE_SEGMENT|4377,4383|false|false|false|C0333138|Stasis|stasis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4377,4394|true|false|false|C0011620|Stasis dermatitis|stasis dermatitis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4384,4394|true|false|false|C0011603|Dermatitis|dermatitis
Event|Event|SIMPLE_SEGMENT|4384,4394|false|false|false|||dermatitis
Event|Event|SIMPLE_SEGMENT|4396,4402|false|false|false|||ulcers
Finding|Pathologic Function|SIMPLE_SEGMENT|4396,4402|true|false|false|C0041582|Ulcer|ulcers
Event|Event|SIMPLE_SEGMENT|4404,4409|false|false|false|||scars
Finding|Finding|SIMPLE_SEGMENT|4404,4409|true|false|false|C0241158;C2004491|Cicatrix;Scar Tissue|scars
Finding|Pathologic Function|SIMPLE_SEGMENT|4404,4409|true|false|false|C0241158;C2004491|Cicatrix;Scar Tissue|scars
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4414,4423|true|false|false|C0302314|Xanthoma|xanthomas
Event|Event|SIMPLE_SEGMENT|4414,4423|false|false|false|||xanthomas
Drug|Food|SIMPLE_SEGMENT|4427,4433|false|false|false|C5890763||PULSES
Event|Event|SIMPLE_SEGMENT|4427,4433|false|false|false|||PULSES
Finding|Physiologic Function|SIMPLE_SEGMENT|4427,4433|false|false|false|C0391850|Physiologic pulse|PULSES
Procedure|Health Care Activity|SIMPLE_SEGMENT|4427,4433|false|false|false|C0034107|Pulse taking|PULSES
Finding|Conceptual Entity|SIMPLE_SEGMENT|4438,4444|false|false|false|C0442038;C0920847|Circumpennate;Radial|radial
Event|Event|SIMPLE_SEGMENT|4445,4448|false|false|false|||DPP
Finding|Gene or Genome|SIMPLE_SEGMENT|4445,4448|false|false|false|C1414174;C5848994|DSPP gene;DSPP wt Allele|DPP
Event|Event|SIMPLE_SEGMENT|4472,4476|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|4472,4476|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|4472,4476|false|false|false|C0582103|Medical Examination|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|4499,4508|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|SIMPLE_SEGMENT|4509,4513|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4509,4513|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4528,4533|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4528,4533|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4528,4533|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|4534,4537|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|4542,4545|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4542,4545|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4542,4545|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4552,4555|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4552,4555|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|4552,4555|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4552,4555|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4561,4564|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4561,4564|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|4571,4574|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|4571,4574|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4571,4574|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4571,4574|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4571,4574|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|4578,4581|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4578,4581|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|4578,4581|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|4578,4581|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|4578,4581|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4578,4581|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4588,4592|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4607,4610|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4627,4632|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4627,4632|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4627,4632|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4637,4640|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|SIMPLE_SEGMENT|4637,4640|false|false|false|||PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4637,4640|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4662,4667|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4662,4667|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4662,4667|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|4662,4675|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4662,4675|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4662,4675|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4668,4675|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|4668,4675|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4668,4675|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|4668,4675|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4668,4675|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4668,4675|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4721,4725|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4721,4725|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4721,4725|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4750,4755|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4750,4755|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4750,4755|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4756,4759|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4756,4759|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|4756,4759|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|4756,4759|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|4756,4759|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|4756,4759|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|4756,4759|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4756,4759|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4763,4766|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4763,4766|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4763,4766|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4763,4766|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|4763,4766|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|4763,4766|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|4763,4766|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4770,4777|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|SIMPLE_SEGMENT|4770,4777|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4805,4810|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4805,4810|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4805,4810|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4811,4817|false|false|false|C0023764|lipase|Lipase
Drug|Enzyme|SIMPLE_SEGMENT|4811,4817|false|false|false|C0023764|lipase|Lipase
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4811,4817|false|false|false|C0023764|lipase|Lipase
Event|Event|SIMPLE_SEGMENT|4811,4817|false|false|false|||Lipase
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4811,4817|false|false|false|C0373670|Lipase measurement|Lipase
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4834,4839|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4834,4839|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4834,4839|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4866,4871|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4866,4871|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4866,4871|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4872,4877|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|SIMPLE_SEGMENT|4872,4877|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|SIMPLE_SEGMENT|4872,4877|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4872,4877|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Event|Event|SIMPLE_SEGMENT|4875,4877|false|false|false|||MB
Finding|Gene or Genome|SIMPLE_SEGMENT|4875,4879|false|false|false|C1413238;C3273407|CD79A gene;CD79A wt Allele|MB-1
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4906,4911|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4906,4911|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4906,4911|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4906,4919|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4912,4919|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4912,4919|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4912,4919|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4912,4919|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|4912,4919|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|4912,4919|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|4912,4919|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4912,4919|false|false|false|C0201925|Calcium measurement|Calcium
Event|Event|SIMPLE_SEGMENT|4941,4944|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4941,4944|false|false|false|C0039985|Plain chest X-ray|CXR
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4950,4958|false|false|false|C2926606||FINDINGS
Event|Event|SIMPLE_SEGMENT|4950,4958|false|false|false|||FINDINGS
Finding|Functional Concept|SIMPLE_SEGMENT|4950,4958|false|false|false|C2607943|findings aspects|FINDINGS
Event|Event|SIMPLE_SEGMENT|4982,4987|false|false|false|||views
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4995,5000|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|4995,5000|false|false|false|C0741025|Chest problem|chest
Event|Event|SIMPLE_SEGMENT|5024,5032|false|false|false|||blunting
Finding|Functional Concept|SIMPLE_SEGMENT|5036,5040|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5036,5059|false|false|false|C0504100|Left costodiaphragmatic recess|left costophrenic angle
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5041,5059|false|false|false|C0230151|Costophrenic angle|costophrenic angle
Event|Event|SIMPLE_SEGMENT|5070,5080|false|false|false|||suggestive
Finding|Functional Concept|SIMPLE_SEGMENT|5070,5080|false|false|false|C0332299|Suggestive of|suggestive
Finding|Functional Concept|SIMPLE_SEGMENT|5070,5083|false|false|false|C0332299|Suggestive of|suggestive of
Event|Event|SIMPLE_SEGMENT|5096,5104|false|false|false|||scarring
Finding|Pathologic Function|SIMPLE_SEGMENT|5096,5104|false|false|false|C0008767;C2004491|Cicatrix;Cicatrization|scarring
Anatomy|Tissue|SIMPLE_SEGMENT|5108,5115|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5108,5115|false|false|false|C0032226|Pleural Diseases|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5108,5126|false|false|false|C0264545|Thickening of pleura|pleural thickening
Event|Event|SIMPLE_SEGMENT|5116,5126|false|false|false|||thickening
Finding|Finding|SIMPLE_SEGMENT|5116,5126|false|false|false|C0205400|Thickened|thickening
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5133,5138|false|false|false|C0024109|Lung|lungs
Event|Event|SIMPLE_SEGMENT|5154,5159|false|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|5154,5159|false|false|false|C1550016|Remote control command - Clear|clear
Event|Event|SIMPLE_SEGMENT|5201,5207|false|false|false|||normal
Event|Event|SIMPLE_SEGMENT|5209,5215|false|false|false|||limits
Finding|Functional Concept|SIMPLE_SEGMENT|5209,5215|false|false|false|C0439801|Limited (extensiveness)|limits
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5218,5235|false|false|false|C1282959|Median Sternotomy|Median sternotomy
Event|Event|SIMPLE_SEGMENT|5225,5235|false|false|false|||sternotomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5225,5235|false|false|false|C0185792|Sternotomy (procedure)|sternotomy
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5246,5257|false|false|false|C0025066|Mediastinum|mediastinal
Event|Event|SIMPLE_SEGMENT|5258,5263|false|false|false|||clips
Event|Event|SIMPLE_SEGMENT|5271,5276|false|false|false|||noted
Event|Event|SIMPLE_SEGMENT|5280,5290|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|5280,5290|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|5280,5290|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|5297,5302|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5303,5318|false|false|false|C0553534|Cardiopulmonary|cardiopulmonary
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5303,5318|false|false|false|C4072686|Cardiovascular disease+Pulmonary disease|cardiopulmonary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5319,5326|false|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5319,5326|true|false|false|C1951340|Process Pharmacologic Substance|process
Event|Event|SIMPLE_SEGMENT|5319,5326|false|false|false|||process
Finding|Functional Concept|SIMPLE_SEGMENT|5319,5326|true|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|5319,5326|true|false|false|C1522240|Process|process
Event|Event|SIMPLE_SEGMENT|5329,5337|false|false|false|||Exercise
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|5329,5337|false|false|false|C0015259|Exercise|Exercise
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5329,5337|false|false|false|C1522704|Exercise Pain Management|Exercise
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5338,5344|false|false|false|C1718621|W stress|Stress
Drug|Organic Chemical|SIMPLE_SEGMENT|5338,5344|false|false|false|C0723460|Stress bismuth subsalicylate|Stress
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5338,5344|false|false|false|C0723460|Stress bismuth subsalicylate|Stress
Event|Event|SIMPLE_SEGMENT|5338,5344|false|false|false|||Stress
Finding|Finding|SIMPLE_SEGMENT|5338,5344|false|false|false|C0038435|Stress|Stress
Event|Event|SIMPLE_SEGMENT|5350,5360|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|5350,5360|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|5350,5360|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Finding|SIMPLE_SEGMENT|5362,5370|false|false|false|C0741302|atypia morphology|Atypical
Finding|Intellectual Product|SIMPLE_SEGMENT|5371,5383|false|false|false|C1272517|Sudden onset (contextual qualifier) (qualifier value)|sudden onset
Finding|Intellectual Product|SIMPLE_SEGMENT|5371,5386|false|false|false|C1272517|Sudden onset (contextual qualifier) (qualifier value)|sudden onset of
Event|Event|SIMPLE_SEGMENT|5378,5383|false|false|false|||onset
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5387,5392|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|5387,5392|false|false|false|C0741025|Chest problem|chest
Finding|Sign or Symptom|SIMPLE_SEGMENT|5387,5402|false|false|false|C0232292|Chest tightness|chest tightness
Event|Event|SIMPLE_SEGMENT|5393,5402|false|false|false|||tightness
Finding|Finding|SIMPLE_SEGMENT|5422,5432|false|false|false|C0429029|ST segment|ST segment
Event|Event|SIMPLE_SEGMENT|5433,5440|false|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|5433,5440|false|false|false|C0392747|Changing|changes
Event|Event|SIMPLE_SEGMENT|5444,5452|false|false|false|||achieved
Finding|Finding|SIMPLE_SEGMENT|5453,5456|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|SIMPLE_SEGMENT|5453,5456|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Event|Event|SIMPLE_SEGMENT|5457,5465|false|false|false|||workload
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|5468,5475|false|false|false|C0035253|Rest|Resting
Finding|Intellectual Product|SIMPLE_SEGMENT|5476,5480|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5481,5489|false|false|false|C0039155|Systole|systolic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5481,5502|false|false|false|C0221155|Systolic Hypertension|systolic hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5490,5502|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|SIMPLE_SEGMENT|5490,5502|false|false|false|||hypertension
Event|Event|SIMPLE_SEGMENT|5518,5529|false|false|false|||hemodynamic
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5518,5529|false|false|false|C0019010|Hemodynamics|hemodynamic
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5518,5529|false|false|false|C4281788|hemodynamics (procedure)|hemodynamic
Event|Event|SIMPLE_SEGMENT|5531,5539|false|false|false|||response
Finding|Finding|SIMPLE_SEGMENT|5531,5539|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Intellectual Product|SIMPLE_SEGMENT|5531,5539|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Mental Process|SIMPLE_SEGMENT|5531,5539|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Organism Function|SIMPLE_SEGMENT|5531,5551|false|false|false|C2265833|response to exercise|response to exercise
Event|Event|SIMPLE_SEGMENT|5543,5551|false|false|false|||exercise
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|5543,5551|false|false|false|C0015259|Exercise|exercise
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5543,5551|false|false|false|C1522704|Exercise Pain Management|exercise
Procedure|Health Care Activity|SIMPLE_SEGMENT|5553,5557|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|Echo
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5553,5557|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|Echo
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5558,5564|false|false|false|C4255046||report
Event|Event|SIMPLE_SEGMENT|5558,5564|false|false|false|||report
Finding|Intellectual Product|SIMPLE_SEGMENT|5558,5564|false|false|false|C0684224|Report (document)|report
Procedure|Health Care Activity|SIMPLE_SEGMENT|5558,5564|false|false|false|C0700287|Reporting|report
Event|Event|SIMPLE_SEGMENT|5565,5569|false|false|false|||sent
Event|Event|SIMPLE_SEGMENT|5583,5591|false|false|false|||Exercise
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|5583,5591|false|false|false|C0015259|Exercise|Exercise
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5583,5591|false|false|false|C1522704|Exercise Pain Management|Exercise
Procedure|Health Care Activity|SIMPLE_SEGMENT|5592,5596|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|Echo
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5592,5596|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|Echo
Event|Event|SIMPLE_SEGMENT|5602,5612|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|5602,5612|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|5602,5612|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|5614,5618|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|Poor
Finding|Conceptual Entity|SIMPLE_SEGMENT|5619,5629|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|functional
Finding|Functional Concept|SIMPLE_SEGMENT|5619,5629|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|functional
Event|Event|SIMPLE_SEGMENT|5630,5638|false|false|false|||exercise
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|5630,5638|false|false|false|C0015259|Exercise|exercise
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5630,5638|false|false|false|C1522704|Exercise Pain Management|exercise
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5662,5665|false|false|false|C0018064|Equine Gonadotropins|ECG
Drug|Hormone|SIMPLE_SEGMENT|5662,5665|false|false|false|C0018064|Equine Gonadotropins|ECG
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5662,5665|false|false|false|C0018064|Equine Gonadotropins|ECG
Event|Event|SIMPLE_SEGMENT|5662,5665|false|false|false|||ECG
Finding|Intellectual Product|SIMPLE_SEGMENT|5662,5665|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|ECG
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5662,5665|false|false|false|C1623258|Electrocardiography|ECG
Event|Event|SIMPLE_SEGMENT|5667,5674|false|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|5667,5674|false|false|false|C0392747|Changing|changes
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|5682,5689|false|false|false|C1689985|Absence (morphologic abnormality)|absence
Event|Event|SIMPLE_SEGMENT|5682,5689|false|false|false|||absence
Finding|Functional Concept|SIMPLE_SEGMENT|5682,5689|false|false|false|C0332197|Absent|absence
Finding|Functional Concept|SIMPLE_SEGMENT|5682,5692|false|false|false|C0332197|Absent|absence of
Event|Event|SIMPLE_SEGMENT|5714,5722|false|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|5714,5722|false|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|5714,5725|false|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Finding|Functional Concept|SIMPLE_SEGMENT|5727,5736|false|false|false|C0205263|Induce (action)|inducible
Event|Event|SIMPLE_SEGMENT|5737,5745|false|false|false|||ischemia
Finding|Pathologic Function|SIMPLE_SEGMENT|5737,5745|false|false|false|C0022116|Ischemia|ischemia
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5737,5745|false|false|false|C4321499|Ischemia Procedure|ischemia
Finding|Finding|SIMPLE_SEGMENT|5758,5761|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|SIMPLE_SEGMENT|5758,5761|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Event|Event|SIMPLE_SEGMENT|5762,5770|false|false|false|||workload
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|5772,5779|false|false|false|C0035253|Rest|Resting
Finding|Intellectual Product|SIMPLE_SEGMENT|5780,5784|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5786,5794|false|false|false|C0039155|Systole|systolic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5786,5807|false|false|false|C0221155|Systolic Hypertension|systolic hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5795,5807|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|SIMPLE_SEGMENT|5795,5807|false|false|false|||hypertension
Event|Event|SIMPLE_SEGMENT|5823,5834|false|false|false|||hemodynamic
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5823,5834|false|false|false|C0019010|Hemodynamics|hemodynamic
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5823,5834|false|false|false|C4281788|hemodynamics (procedure)|hemodynamic
Event|Event|SIMPLE_SEGMENT|5835,5843|false|false|false|||response
Finding|Finding|SIMPLE_SEGMENT|5835,5843|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Intellectual Product|SIMPLE_SEGMENT|5835,5843|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Mental Process|SIMPLE_SEGMENT|5835,5843|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Event|Event|SIMPLE_SEGMENT|5848,5859|false|false|false|||physiologic
Finding|Functional Concept|SIMPLE_SEGMENT|5848,5859|false|false|false|C0205463|Physiological|physiologic
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5860,5866|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|SIMPLE_SEGMENT|5860,5866|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5860,5866|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Event|Event|SIMPLE_SEGMENT|5860,5866|false|false|false|||stress
Finding|Finding|SIMPLE_SEGMENT|5860,5866|false|false|false|C0038435|Stress|stress
Finding|Body Substance|SIMPLE_SEGMENT|5870,5879|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|5870,5879|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|5870,5879|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|5870,5879|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|SIMPLE_SEGMENT|5880,5884|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5880,5884|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5899,5904|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5899,5904|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5899,5904|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|5905,5908|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|5913,5916|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5913,5916|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5913,5916|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5923,5926|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5923,5926|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|5923,5926|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5923,5926|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5932,5935|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5932,5935|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|5943,5946|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|5943,5946|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5943,5946|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5943,5946|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5943,5946|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|5950,5953|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5950,5953|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|5950,5953|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|5950,5953|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|5950,5953|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5950,5953|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5960,5964|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5979,5982|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5999,6004|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5999,6004|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5999,6004|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Event|SIMPLE_SEGMENT|6017,6018|false|false|false|||-
Drug|Inorganic Chemical|SIMPLE_SEGMENT|6034,6038|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6034,6038|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6034,6038|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6064,6069|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|6064,6069|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|6064,6069|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6101,6105|false|false|false|C0270724|Infantile Neuroaxonal Dystrophy|PLAN
Event|Event|SIMPLE_SEGMENT|6101,6105|false|false|false|||PLAN
Finding|Functional Concept|SIMPLE_SEGMENT|6101,6105|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|PLAN
Finding|Intellectual Product|SIMPLE_SEGMENT|6101,6105|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|PLAN
Finding|Mental Process|SIMPLE_SEGMENT|6101,6105|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|PLAN
Finding|Finding|SIMPLE_SEGMENT|6111,6114|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|pmh
Finding|Finding|SIMPLE_SEGMENT|6115,6121|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|6115,6121|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6128,6131|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6128,6131|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|6128,6131|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|6128,6131|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|6128,6131|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6128,6131|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|6128,6131|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6128,6131|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|SIMPLE_SEGMENT|6136,6140|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6136,6140|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Finding|Intellectual Product|SIMPLE_SEGMENT|6147,6154|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|6147,6154|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6156,6162|false|false|false|C2926611||angina
Event|Event|SIMPLE_SEGMENT|6156,6162|false|false|false|||angina
Finding|Finding|SIMPLE_SEGMENT|6156,6162|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Finding|Sign or Symptom|SIMPLE_SEGMENT|6156,6162|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6170,6173|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|6170,6173|false|false|false|||HTN
Event|Event|SIMPLE_SEGMENT|6182,6190|false|false|false|||presents
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6196,6201|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|6196,6201|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6196,6206|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6196,6206|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6202,6206|false|true|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|6202,6206|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|6202,6206|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6202,6206|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|6208,6218|false|false|false|||concerning
Drug|Hormone|SIMPLE_SEGMENT|6223,6232|false|false|false|C3273442|Crescendo|crescendo
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6223,6232|false|false|false|C3273442|Crescendo|crescendo
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6223,6239|false|false|false|C0002965|Angina, Unstable|crescendo angina
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6233,6239|false|false|false|C2926611||angina
Event|Event|SIMPLE_SEGMENT|6233,6239|false|false|false|||angina
Finding|Finding|SIMPLE_SEGMENT|6233,6239|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Finding|Sign or Symptom|SIMPLE_SEGMENT|6233,6239|false|false|false|C0002962;C2024883|Angina Pectoris|angina
Event|Event|SIMPLE_SEGMENT|6249,6255|false|false|false|||ISSUES
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6260,6265|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|SIMPLE_SEGMENT|6260,6265|false|false|false|C0741025|Chest problem|Chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6260,6270|false|false|false|C2926613||Chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6260,6270|false|false|false|C0008031|Chest Pain|Chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6266,6270|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|6266,6270|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|6266,6270|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6266,6270|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Body Substance|SIMPLE_SEGMENT|6272,6279|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6272,6279|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6272,6279|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|SIMPLE_SEGMENT|6285,6289|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|SIMPLE_SEGMENT|6285,6289|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|SIMPLE_SEGMENT|6285,6289|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6290,6298|false|false|false|C0018787|Heart|coronary
Event|Event|SIMPLE_SEGMENT|6299,6303|false|false|false|||risk
Finding|Idea or Concept|SIMPLE_SEGMENT|6299,6303|false|false|false|C0035647|Risk|risk
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|6320,6323|false|false|false|C0041207|Truncus Arteriosus, Persistent|cat
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6320,6323|false|false|false|C0008169;C1443200;C3530118|CAT protein, human;Cat hair antigen;Chloramphenicol O-Acetyltransferase|cat
Drug|Enzyme|SIMPLE_SEGMENT|6320,6323|false|false|false|C0008169;C1443200;C3530118|CAT protein, human;Cat hair antigen;Chloramphenicol O-Acetyltransferase|cat
Drug|Immunologic Factor|SIMPLE_SEGMENT|6320,6323|false|false|false|C0008169;C1443200;C3530118|CAT protein, human;Cat hair antigen;Chloramphenicol O-Acetyltransferase|cat
Event|Event|SIMPLE_SEGMENT|6320,6323|false|false|false|||cat
Finding|Gene or Genome|SIMPLE_SEGMENT|6320,6323|false|false|false|C1151515;C1366498;C1413138;C4050461;C4758039|CAT gene;Chloramphenicol Acetyl Transferase Gene;Chronic Obstructive Pulmonary Disease Assessment Test scale;Cutaneous Assessment Tool;catalase activity|cat
Finding|Intellectual Product|SIMPLE_SEGMENT|6320,6323|false|false|false|C1151515;C1366498;C1413138;C4050461;C4758039|CAT gene;Chloramphenicol Acetyl Transferase Gene;Chronic Obstructive Pulmonary Disease Assessment Test scale;Cutaneous Assessment Tool;catalase activity|cat
Finding|Molecular Function|SIMPLE_SEGMENT|6320,6323|false|false|false|C1151515;C1366498;C1413138;C4050461;C4758039|CAT gene;Chloramphenicol Acetyl Transferase Gene;Chronic Obstructive Pulmonary Disease Assessment Test scale;Cutaneous Assessment Tool;catalase activity|cat
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6320,6323|false|false|false|C0040405;C0280589;C2097305|X-Ray Computed Tomography;allergy testing cat;cytarabine/thioguanine protocol|cat
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6320,6323|false|false|false|C0040405;C0280589;C2097305|X-Ray Computed Tomography;allergy testing cat;cytarabine/thioguanine protocol|cat
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6320,6323|false|false|false|C0040405;C0280589;C2097305|X-Ray Computed Tomography;allergy testing cat;cytarabine/thioguanine protocol|cat
Finding|Gene or Genome|SIMPLE_SEGMENT|6334,6337|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|SIMPLE_SEGMENT|6346,6352|false|false|false|||reveal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6367,6374|true|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|6367,6374|false|false|false|||disease
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6377,6381|false|false|false|C5552605|FACT Complex|Fact
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6377,6381|false|false|false|C5552605|FACT Complex|Fact
Finding|Gene or Genome|SIMPLE_SEGMENT|6377,6381|false|false|false|C1420522;C5551287|SSRP1 wt Allele;SUPT16H gene|Fact
Event|Event|SIMPLE_SEGMENT|6402,6417|false|false|false|||reproducability
Finding|Finding|SIMPLE_SEGMENT|6421,6429|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Finding|Functional Concept|SIMPLE_SEGMENT|6421,6429|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|6421,6429|false|false|false|C0031809|Physical Examination|physical
Finding|Finding|SIMPLE_SEGMENT|6421,6434|false|false|false|C1509143|physical examination (physical finding)|physical exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|6421,6434|false|false|false|C0031809|Physical Examination|physical exam
Event|Event|SIMPLE_SEGMENT|6430,6434|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|6430,6434|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|6430,6434|false|false|false|C0582103|Medical Examination|exam
Event|Event|SIMPLE_SEGMENT|6435,6443|false|false|false|||suggests
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6449,6456|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|6449,6456|false|false|false|C1314974|Cardiac attachment|cardiac
Event|Event|SIMPLE_SEGMENT|6457,6462|false|false|false|||cause
Finding|Conceptual Entity|SIMPLE_SEGMENT|6457,6462|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Finding|Functional Concept|SIMPLE_SEGMENT|6457,6462|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Event|Event|SIMPLE_SEGMENT|6472,6480|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|6472,6480|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|6472,6480|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|SIMPLE_SEGMENT|6485,6496|false|false|false|||complicated
Finding|Body Substance|SIMPLE_SEGMENT|6500,6507|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6500,6507|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6500,6507|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|6511,6518|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|6511,6518|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|6511,6518|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|6511,6518|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|6511,6521|false|false|false|C0262926|Medical History|history of
Finding|Functional Concept|SIMPLE_SEGMENT|6522,6531|false|false|false|C1516691|Cognitive|cognitive
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|6522,6542|false|false|false|C0338656|Impaired cognition|cognitive impairment
Event|Event|SIMPLE_SEGMENT|6532,6542|false|false|false|||impairment
Finding|Finding|SIMPLE_SEGMENT|6532,6542|false|false|false|C0221099;C0684336|Impaired;Impaired health|impairment
Finding|Functional Concept|SIMPLE_SEGMENT|6532,6542|false|false|false|C0221099;C0684336|Impaired;Impaired health|impairment
Event|Event|SIMPLE_SEGMENT|6551,6556|false|false|false|||known
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6557,6560|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6557,6560|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|6557,6560|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|6557,6560|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|6557,6560|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6557,6560|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|6557,6560|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6557,6560|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|SIMPLE_SEGMENT|6571,6579|false|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|6571,6579|false|false|false|C1261287|Stenosis|stenosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6580,6586|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|SIMPLE_SEGMENT|6580,6586|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6580,6586|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Finding|Finding|SIMPLE_SEGMENT|6580,6586|false|false|false|C0038435|Stress|stress
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6580,6591|false|false|false|C0920208|Echocardiography, Stress|stress echo
Event|Event|SIMPLE_SEGMENT|6587,6591|false|false|false|||echo
Procedure|Health Care Activity|SIMPLE_SEGMENT|6587,6591|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6587,6591|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Event|Event|SIMPLE_SEGMENT|6609,6615|false|false|false|||assess
Event|Event|SIMPLE_SEGMENT|6620,6630|false|false|false|||functional
Finding|Conceptual Entity|SIMPLE_SEGMENT|6620,6630|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|functional
Finding|Functional Concept|SIMPLE_SEGMENT|6620,6630|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|functional
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|6632,6643|false|false|false|C0000768|Congenital Abnormality|abnormality
Event|Event|SIMPLE_SEGMENT|6632,6643|false|false|false|||abnormality
Finding|Finding|SIMPLE_SEGMENT|6632,6643|false|false|false|C1704258|Abnormality|abnormality
Event|Event|SIMPLE_SEGMENT|6649,6657|false|false|false|||exertion
Finding|Organism Function|SIMPLE_SEGMENT|6649,6657|false|false|false|C0015264|Exertion|exertion
Event|Event|SIMPLE_SEGMENT|6663,6667|false|false|false|||ECHO
Procedure|Health Care Activity|SIMPLE_SEGMENT|6663,6667|true|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6663,6667|true|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|6668,6681|true|false|false|C0000768|Congenital Abnormality|abnormalities
Event|Event|SIMPLE_SEGMENT|6668,6681|false|false|false|||abnormalities
Finding|Functional Concept|SIMPLE_SEGMENT|6668,6681|true|false|false|C0000769|teratologic|abnormalities
Event|Event|SIMPLE_SEGMENT|6687,6692|false|false|false|||noted
Event|Event|SIMPLE_SEGMENT|6706,6714|false|false|false|||reported
Finding|Finding|SIMPLE_SEGMENT|6715,6723|false|false|false|C0741302|atypia morphology|atypical
Finding|Sign or Symptom|SIMPLE_SEGMENT|6715,6734|false|true|false|C0262384|Atypical chest pain|atypical chest pain
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6724,6729|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|6724,6729|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6724,6734|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6724,6734|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6730,6734|false|true|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|6730,6734|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|6730,6734|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6730,6734|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6740,6746|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|SIMPLE_SEGMENT|6740,6746|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6740,6746|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Event|Event|SIMPLE_SEGMENT|6740,6746|false|false|false|||stress
Finding|Finding|SIMPLE_SEGMENT|6740,6746|false|false|false|C0038435|Stress|stress
Event|Event|SIMPLE_SEGMENT|6758,6767|false|false|false|||continued
Finding|Idea or Concept|SIMPLE_SEGMENT|6771,6775|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|6771,6775|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|6771,6775|false|false|false|C1553498|home health encounter|home
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6776,6779|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Enzyme|SIMPLE_SEGMENT|6776,6779|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Organic Chemical|SIMPLE_SEGMENT|6776,6779|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6776,6779|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Event|Event|SIMPLE_SEGMENT|6776,6779|false|false|false|||ASA
Finding|Gene or Genome|SIMPLE_SEGMENT|6776,6779|false|false|false|C1412553|ARSA gene|ASA
Drug|Organic Chemical|SIMPLE_SEGMENT|6781,6787|false|false|false|C0633084|Plavix|plavix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6781,6787|false|false|false|C0633084|Plavix|plavix
Event|Event|SIMPLE_SEGMENT|6781,6787|false|false|false|||plavix
Drug|Organic Chemical|SIMPLE_SEGMENT|6789,6795|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|statin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6789,6795|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|statin
Event|Event|SIMPLE_SEGMENT|6789,6795|false|false|false|||statin
Finding|Gene or Genome|SIMPLE_SEGMENT|6789,6795|false|false|false|C1414273|EEF1A2 gene|statin
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|6797,6804|false|false|false|C0028125;C0699857;C3848573|Nitrate;Nitrates;nitrate ion|nitrate
Drug|Inorganic Chemical|SIMPLE_SEGMENT|6797,6804|false|false|false|C0028125;C0699857;C3848573|Nitrate;Nitrates;nitrate ion|nitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6797,6804|false|false|false|C0028125;C0699857;C3848573|Nitrate;Nitrates;nitrate ion|nitrate
Event|Event|SIMPLE_SEGMENT|6797,6804|false|false|false|||nitrate
Drug|Organic Chemical|SIMPLE_SEGMENT|6809,6819|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6809,6819|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|SIMPLE_SEGMENT|6809,6819|false|false|false|||metoprolol
Finding|Idea or Concept|SIMPLE_SEGMENT|6827,6835|false|false|false|C4288901|In-House|in-house
Event|Event|SIMPLE_SEGMENT|6846,6855|false|false|false|||monitored
Event|Event|SIMPLE_SEGMENT|6859,6863|false|false|false|||tele
Finding|Gene or Genome|SIMPLE_SEGMENT|6859,6863|false|false|false|C1420621;C1515258|TCAP gene;Telephone Number|tele
Finding|Intellectual Product|SIMPLE_SEGMENT|6859,6863|false|false|false|C1420621;C1515258|TCAP gene;Telephone Number|tele
Event|Event|SIMPLE_SEGMENT|6876,6882|false|false|false|||alarms
Finding|Intellectual Product|SIMPLE_SEGMENT|6876,6882|true|false|false|C3484361|Alarms (package insert)|alarms
Event|Event|SIMPLE_SEGMENT|6894,6904|false|false|false|||discharged
Event|Event|SIMPLE_SEGMENT|6905,6909|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|6905,6909|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|6905,6909|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|6905,6909|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|6918,6926|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|6918,6926|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|6918,6926|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6918,6926|false|false|false|C5237010|Expression Negative|negative
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6927,6933|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|SIMPLE_SEGMENT|6927,6933|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6927,6933|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Event|Event|SIMPLE_SEGMENT|6927,6933|false|false|false|||stress
Finding|Finding|SIMPLE_SEGMENT|6927,6933|false|false|false|C0038435|Stress|stress
Event|Event|SIMPLE_SEGMENT|6937,6943|false|false|false|||follow
Finding|Functional Concept|SIMPLE_SEGMENT|6937,6943|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|6937,6943|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|SIMPLE_SEGMENT|6937,6946|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|SIMPLE_SEGMENT|6937,6946|false|false|false|C1522577|follow-up|follow-up
Event|Event|SIMPLE_SEGMENT|6944,6946|false|false|false|||up
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6957,6960|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|6957,6960|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6957,6960|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6957,6960|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|6957,6960|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|6957,6960|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|6957,6960|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6957,6960|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|6957,6960|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|6957,6960|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|6957,6960|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|SIMPLE_SEGMENT|6971,6978|false|false|false|||CHRONIC
Finding|Intellectual Product|SIMPLE_SEGMENT|6971,6978|false|false|false|C1547296|Chronic - Admission Level of Care Code|CHRONIC
Procedure|Health Care Activity|SIMPLE_SEGMENT|6971,6978|false|false|false|C1555457|Provision of recurring care for chronic illness|CHRONIC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6992,7001|false|false|false|C0012000|Diastole|Diastolic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6992,7005|false|false|false|C2183328|diastolic congestive heart failure|Diastolic CHF
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|7002,7005|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7002,7005|false|false|false|C0018802|Congestive heart failure|CHF
Event|Event|SIMPLE_SEGMENT|7002,7005|false|false|false|||CHF
Event|Event|SIMPLE_SEGMENT|7019,7024|false|false|false|||signs
Finding|Finding|SIMPLE_SEGMENT|7019,7024|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|7019,7024|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Drug|Substance|SIMPLE_SEGMENT|7028,7033|true|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|7028,7033|true|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Finding|SIMPLE_SEGMENT|7028,7042|true|false|false|C0546817;C5848920|Fluid Overload;Hypervolemia (finding)|fluid overload
Finding|Pathologic Function|SIMPLE_SEGMENT|7028,7042|true|false|false|C0546817;C5848920|Fluid Overload;Hypervolemia (finding)|fluid overload
Event|Event|SIMPLE_SEGMENT|7034,7042|false|false|false|||overload
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7063,7071|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|SIMPLE_SEGMENT|7063,7071|false|false|false|||baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|7063,7071|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|SIMPLE_SEGMENT|7072,7080|false|false|false|||diuresis
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|7072,7080|false|false|false|C0012797|Diuresis|diuresis
Event|Event|SIMPLE_SEGMENT|7091,7100|false|false|false|||continued
Event|Event|SIMPLE_SEGMENT|7104,7108|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|7104,7108|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|7104,7108|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|7104,7108|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|7125,7134|false|false|false|||monitored
Event|Event|SIMPLE_SEGMENT|7145,7150|false|false|false|||signs
Finding|Finding|SIMPLE_SEGMENT|7145,7150|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|7145,7150|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Event|Event|SIMPLE_SEGMENT|7154,7168|false|false|false|||decompensation
Finding|Finding|SIMPLE_SEGMENT|7154,7168|false|false|false|C0231187|Decompensation|decompensation
Event|Event|SIMPLE_SEGMENT|7173,7181|false|false|false|||required
Event|Event|SIMPLE_SEGMENT|7186,7194|false|false|false|||diuresis
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|7186,7194|false|false|false|C0012797|Diuresis|diuresis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7200,7208|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|Diabetes
Event|Event|SIMPLE_SEGMENT|7200,7208|false|false|false|||Diabetes
Event|Event|SIMPLE_SEGMENT|7211,7215|false|false|false|||HISS
Finding|Intellectual Product|SIMPLE_SEGMENT|7211,7215|false|false|false|C0019972|Hospital Information Systems|HISS
Finding|Idea or Concept|SIMPLE_SEGMENT|7216,7224|false|false|false|C4288901|In-House|in-house
Event|Event|SIMPLE_SEGMENT|7239,7248|false|false|false|||continued
Event|Event|SIMPLE_SEGMENT|7252,7256|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|7252,7256|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|7252,7256|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|7252,7256|false|false|false|C1553498|home health encounter|home
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7258,7265|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|7258,7265|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7258,7265|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|7258,7265|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|7258,7265|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7258,7265|false|false|false|C0202098|Insulin measurement|insulin
Event|Event|SIMPLE_SEGMENT|7266,7273|false|false|false|||regimen
Finding|Intellectual Product|SIMPLE_SEGMENT|7266,7273|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7266,7273|false|false|false|C0040808|Treatment Protocols|regimen
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7282,7288|false|false|false|C0876064|Lantus|lantus
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7282,7288|false|false|false|C0876064|Lantus|lantus
Event|Event|SIMPLE_SEGMENT|7289,7292|false|false|false|||QHS
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7297,7308|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7297,7308|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|7297,7308|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|7297,7308|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|7297,7321|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|SIMPLE_SEGMENT|7312,7321|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|7312,7321|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7340,7350|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|7340,7350|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|7340,7355|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|SIMPLE_SEGMENT|7351,7355|false|false|false|||list
Finding|Intellectual Product|SIMPLE_SEGMENT|7351,7355|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|SIMPLE_SEGMENT|7359,7367|false|false|false|||accurate
Drug|Organic Chemical|SIMPLE_SEGMENT|7372,7380|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7372,7380|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|7372,7380|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|SIMPLE_SEGMENT|7372,7380|false|false|false|||complete
Finding|Functional Concept|SIMPLE_SEGMENT|7372,7380|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|7372,7380|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|SIMPLE_SEGMENT|7385,7393|false|false|false|C0126174|losartan|Losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7385,7393|false|false|false|C0126174|losartan|Losartan
Event|Event|SIMPLE_SEGMENT|7385,7393|false|false|false|||Losartan
Drug|Organic Chemical|SIMPLE_SEGMENT|7385,7403|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7385,7403|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7394,7403|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7394,7403|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|SIMPLE_SEGMENT|7394,7403|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|7394,7403|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7394,7403|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Event|Event|SIMPLE_SEGMENT|7394,7403|false|false|false|||Potassium
Finding|Physiologic Function|SIMPLE_SEGMENT|7394,7403|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7394,7403|false|false|false|C0202194|Potassium measurement|Potassium
Drug|Organic Chemical|SIMPLE_SEGMENT|7423,7430|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7423,7430|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|7450,7462|false|false|false|C0007248|carisoprodol|carisoprodol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7450,7462|false|false|false|C0007248|carisoprodol|carisoprodol
Event|Event|SIMPLE_SEGMENT|7450,7462|false|false|false|||carisoprodol
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|7475,7479|false|false|false|C0226896|Oral cavity|Oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7475,7479|false|false|false|C1272919|Oral Dosage Form|Oral
Finding|Finding|SIMPLE_SEGMENT|7475,7479|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Finding|Functional Concept|SIMPLE_SEGMENT|7475,7479|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Event|Event|SIMPLE_SEGMENT|7484,7489|false|false|false|||spasm
Finding|Gene or Genome|SIMPLE_SEGMENT|7484,7489|false|false|false|C0037763;C3812627|KANTR gene;Spasm|spasm
Finding|Sign or Symptom|SIMPLE_SEGMENT|7484,7489|false|false|false|C0037763;C3812627|KANTR gene;Spasm|spasm
Event|Event|SIMPLE_SEGMENT|7491,7495|false|false|false|||Take
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7498,7504|false|false|false|C0039225|Tablet Dosage Form|tablet
Event|Event|SIMPLE_SEGMENT|7498,7504|false|false|false|||tablet
Finding|Gene or Genome|SIMPLE_SEGMENT|7519,7522|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7523,7529|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|SIMPLE_SEGMENT|7523,7529|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Finding|Sign or Symptom|SIMPLE_SEGMENT|7523,7535|false|false|false|C0037763|Spasm|muscle spasm
Event|Event|SIMPLE_SEGMENT|7530,7535|false|false|false|||spasm
Finding|Gene or Genome|SIMPLE_SEGMENT|7530,7535|false|false|false|C0037763;C3812627|KANTR gene;Spasm|spasm
Finding|Sign or Symptom|SIMPLE_SEGMENT|7530,7535|false|false|false|C0037763;C3812627|KANTR gene;Spasm|spasm
Drug|Organic Chemical|SIMPLE_SEGMENT|7540,7552|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7540,7552|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Organic Chemical|SIMPLE_SEGMENT|7571,7580|false|false|false|C0040805|trazodone|traZODONE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7571,7580|false|false|false|C0040805|trazodone|traZODONE
Drug|Organic Chemical|SIMPLE_SEGMENT|7597,7606|false|false|false|C0030049|oxycodone|Oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7597,7606|false|false|false|C0030049|oxycodone|Oxycodone
Event|Event|SIMPLE_SEGMENT|7597,7606|false|false|false|||Oxycodone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7597,7606|false|false|false|C0524222|Oxycodone measurement|Oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7597,7620|false|false|false|C0717368|acetaminophen / oxycodone|Oxycodone-Acetaminophen
Drug|Organic Chemical|SIMPLE_SEGMENT|7607,7620|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7607,7620|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|SIMPLE_SEGMENT|7607,7620|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7607,7620|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7635,7638|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|SIMPLE_SEGMENT|7635,7638|false|false|false|||TAB
Event|Event|SIMPLE_SEGMENT|7642,7645|false|false|false|||Q8H
Finding|Gene or Genome|SIMPLE_SEGMENT|7646,7649|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7650,7654|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|7650,7654|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|7650,7654|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|7650,7654|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|7659,7671|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7659,7671|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|7691,7704|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7691,7704|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Event|Event|SIMPLE_SEGMENT|7691,7704|false|false|false|||Nitroglycerin
Finding|Gene or Genome|SIMPLE_SEGMENT|7718,7721|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7722,7727|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|7722,7727|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7722,7732|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|7722,7732|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7728,7732|false|true|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|7728,7732|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|7728,7732|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|7728,7732|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|7737,7747|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7737,7747|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|7737,7757|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7737,7757|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|7748,7757|false|false|false|C0038617;C0220918|Succinates;succinate|Succinate
Event|Event|SIMPLE_SEGMENT|7748,7757|false|false|false|||Succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|7782,7792|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7782,7792|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|SIMPLE_SEGMENT|7782,7804|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7782,7804|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Event|Event|SIMPLE_SEGMENT|7793,7804|false|false|false|||Mononitrate
Finding|Finding|SIMPLE_SEGMENT|7806,7814|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|7806,7814|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|SIMPLE_SEGMENT|7815,7822|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|7815,7822|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|7815,7822|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7815,7822|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|SIMPLE_SEGMENT|7845,7856|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7845,7856|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Organic Chemical|SIMPLE_SEGMENT|7877,7888|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7877,7888|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|SIMPLE_SEGMENT|7877,7888|false|false|false|||Fluticasone
Drug|Organic Chemical|SIMPLE_SEGMENT|7877,7899|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7877,7899|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|SIMPLE_SEGMENT|7889,7899|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Event|Event|SIMPLE_SEGMENT|7909,7913|false|false|false|||PUFF
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7917,7920|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7917,7920|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7917,7920|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|7917,7920|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|7917,7920|false|false|false|C1332410|BID gene|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7949,7956|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Hormone|SIMPLE_SEGMENT|7949,7956|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7949,7956|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Event|Event|SIMPLE_SEGMENT|7949,7956|false|false|false|||Insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|7949,7956|false|false|false|C1337112|INS gene|Insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7949,7956|false|false|false|C0202098|Insulin measurement|Insulin
Event|Event|SIMPLE_SEGMENT|7960,7967|false|false|false|||Sliding
Finding|Functional Concept|SIMPLE_SEGMENT|7960,7967|false|false|false|C0332246|Sliding|Sliding
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7960,7973|false|false|false|C2937251|sliding scale|Sliding Scale
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7968,7973|false|false|false|C0222045|Integumentary scale|Scale
Event|Activity|SIMPLE_SEGMENT|7968,7973|false|false|false|C1947916|Scaling|Scale
Finding|Conceptual Entity|SIMPLE_SEGMENT|7968,7973|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|Scale
Finding|Intellectual Product|SIMPLE_SEGMENT|7968,7973|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|Scale
Event|Event|SIMPLE_SEGMENT|8000,8008|false|false|false|||Override
Finding|Functional Concept|SIMPLE_SEGMENT|8000,8008|false|false|false|C1547671|Override|Override
Event|Event|SIMPLE_SEGMENT|8010,8016|false|false|false|||Reason
Finding|Idea or Concept|SIMPLE_SEGMENT|8010,8016|false|false|false|C0392360|Indication of (contextual qualifier)|Reason
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8018,8025|false|false|false|C1314782|Levemir|Levemir
Drug|Hormone|SIMPLE_SEGMENT|8018,8025|false|false|false|C1314782|Levemir|Levemir
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8018,8025|false|false|false|C1314782|Levemir|Levemir
Event|Event|SIMPLE_SEGMENT|8040,8048|false|false|false|||pharmacy
Finding|Intellectual Product|SIMPLE_SEGMENT|8040,8048|false|false|false|C1547997;C3244303|Diagnostic Service Section ID - Pharmacy;Pharmacy domain|pharmacy
Procedure|Health Care Activity|SIMPLE_SEGMENT|8040,8048|false|false|false|C0031321|Pharmaceutical Services|pharmacy
Event|Event|SIMPLE_SEGMENT|8049,8053|false|false|false|||list
Finding|Intellectual Product|SIMPLE_SEGMENT|8049,8053|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|SIMPLE_SEGMENT|8057,8066|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|8057,8066|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8057,8066|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8057,8066|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8057,8066|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|8057,8078|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8067,8078|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8067,8078|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|8067,8078|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|8067,8078|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|8083,8090|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8083,8090|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|8110,8122|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8110,8122|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|8142,8153|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8142,8153|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Organic Chemical|SIMPLE_SEGMENT|8173,8184|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8173,8184|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|SIMPLE_SEGMENT|8173,8184|false|false|false|||Fluticasone
Drug|Organic Chemical|SIMPLE_SEGMENT|8173,8195|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8173,8195|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|SIMPLE_SEGMENT|8185,8195|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Event|Event|SIMPLE_SEGMENT|8205,8209|false|false|false|||PUFF
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8213,8216|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8213,8216|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8213,8216|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|8213,8216|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|8213,8216|false|false|false|C1332410|BID gene|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8244,8251|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Hormone|SIMPLE_SEGMENT|8244,8251|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8244,8251|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Event|Event|SIMPLE_SEGMENT|8244,8251|false|false|false|||Insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|8244,8251|false|false|false|C1337112|INS gene|Insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8244,8251|false|false|false|C0202098|Insulin measurement|Insulin
Event|Event|SIMPLE_SEGMENT|8255,8262|false|false|false|||Sliding
Finding|Functional Concept|SIMPLE_SEGMENT|8255,8262|false|false|false|C0332246|Sliding|Sliding
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8255,8268|false|false|false|C2937251|sliding scale|Sliding Scale
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8263,8268|false|false|false|C0222045|Integumentary scale|Scale
Event|Activity|SIMPLE_SEGMENT|8263,8268|false|false|false|C1947916|Scaling|Scale
Finding|Conceptual Entity|SIMPLE_SEGMENT|8263,8268|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|Scale
Finding|Intellectual Product|SIMPLE_SEGMENT|8263,8268|false|false|false|C0349674;C1522412;C2981742|Base Number;Scale - rank;Scale, LOINC Axis 5|Scale
Event|Event|SIMPLE_SEGMENT|8295,8303|false|false|false|||Override
Finding|Functional Concept|SIMPLE_SEGMENT|8295,8303|false|false|false|C1547671|Override|Override
Event|Event|SIMPLE_SEGMENT|8305,8311|false|false|false|||Reason
Finding|Idea or Concept|SIMPLE_SEGMENT|8305,8311|false|false|false|C0392360|Indication of (contextual qualifier)|Reason
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8313,8320|false|false|false|C1314782|Levemir|Levemir
Drug|Hormone|SIMPLE_SEGMENT|8313,8320|false|false|false|C1314782|Levemir|Levemir
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8313,8320|false|false|false|C1314782|Levemir|Levemir
Event|Event|SIMPLE_SEGMENT|8335,8343|false|false|false|||pharmacy
Finding|Intellectual Product|SIMPLE_SEGMENT|8335,8343|false|false|false|C1547997;C3244303|Diagnostic Service Section ID - Pharmacy;Pharmacy domain|pharmacy
Procedure|Health Care Activity|SIMPLE_SEGMENT|8335,8343|false|false|false|C0031321|Pharmaceutical Services|pharmacy
Event|Event|SIMPLE_SEGMENT|8344,8348|false|false|false|||list
Finding|Intellectual Product|SIMPLE_SEGMENT|8344,8348|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Drug|Organic Chemical|SIMPLE_SEGMENT|8353,8361|false|false|false|C0126174|losartan|Losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8353,8361|false|false|false|C0126174|losartan|Losartan
Event|Event|SIMPLE_SEGMENT|8353,8361|false|false|false|||Losartan
Drug|Organic Chemical|SIMPLE_SEGMENT|8353,8371|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8353,8371|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8362,8371|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|8362,8371|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|SIMPLE_SEGMENT|8362,8371|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|8362,8371|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8362,8371|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Event|Event|SIMPLE_SEGMENT|8362,8371|false|false|false|||Potassium
Finding|Physiologic Function|SIMPLE_SEGMENT|8362,8371|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8362,8371|false|false|false|C0202194|Potassium measurement|Potassium
Drug|Organic Chemical|SIMPLE_SEGMENT|8391,8404|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8391,8404|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Event|Event|SIMPLE_SEGMENT|8391,8404|false|false|false|||Nitroglycerin
Finding|Gene or Genome|SIMPLE_SEGMENT|8418,8421|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8422,8427|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|8422,8427|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8422,8432|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|8422,8432|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8428,8432|false|true|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|8428,8432|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|8428,8432|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|8428,8432|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|8437,8449|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8437,8449|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Organic Chemical|SIMPLE_SEGMENT|8468,8477|false|false|false|C0040805|trazodone|traZODONE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8468,8477|false|false|false|C0040805|trazodone|traZODONE
Drug|Organic Chemical|SIMPLE_SEGMENT|8495,8507|false|false|false|C0007248|carisoprodol|carisoprodol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8495,8507|false|false|false|C0007248|carisoprodol|carisoprodol
Event|Event|SIMPLE_SEGMENT|8495,8507|false|false|false|||carisoprodol
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|8520,8524|false|false|false|C0226896|Oral cavity|Oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8520,8524|false|false|false|C1272919|Oral Dosage Form|Oral
Finding|Finding|SIMPLE_SEGMENT|8520,8524|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Finding|Functional Concept|SIMPLE_SEGMENT|8520,8524|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Event|Event|SIMPLE_SEGMENT|8529,8534|false|false|false|||spasm
Finding|Gene or Genome|SIMPLE_SEGMENT|8529,8534|false|false|false|C0037763;C3812627|KANTR gene;Spasm|spasm
Finding|Sign or Symptom|SIMPLE_SEGMENT|8529,8534|false|false|false|C0037763;C3812627|KANTR gene;Spasm|spasm
Drug|Organic Chemical|SIMPLE_SEGMENT|8540,8550|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8540,8550|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|8540,8560|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8540,8560|false|false|false|C0724633|metoprolol succinate|Metoprolol Succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|8551,8560|false|false|false|C0038617;C0220918|Succinates;succinate|Succinate
Event|Event|SIMPLE_SEGMENT|8551,8560|false|false|false|||Succinate
Drug|Organic Chemical|SIMPLE_SEGMENT|8585,8594|false|false|false|C0030049|oxycodone|Oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8585,8594|false|false|false|C0030049|oxycodone|Oxycodone
Event|Event|SIMPLE_SEGMENT|8585,8594|false|false|false|||Oxycodone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8585,8594|false|false|false|C0524222|Oxycodone measurement|Oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8585,8608|false|false|false|C0717368|acetaminophen / oxycodone|Oxycodone-Acetaminophen
Drug|Organic Chemical|SIMPLE_SEGMENT|8595,8608|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8595,8608|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|SIMPLE_SEGMENT|8595,8608|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8595,8608|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8623,8626|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|SIMPLE_SEGMENT|8623,8626|false|false|false|||TAB
Event|Event|SIMPLE_SEGMENT|8630,8633|false|false|false|||Q8H
Finding|Gene or Genome|SIMPLE_SEGMENT|8634,8637|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8638,8642|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|8638,8642|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|8638,8642|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|8638,8642|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|8648,8658|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8648,8658|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|SIMPLE_SEGMENT|8648,8670|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8648,8670|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Event|Event|SIMPLE_SEGMENT|8659,8670|false|false|false|||Mononitrate
Finding|Finding|SIMPLE_SEGMENT|8672,8680|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|8672,8680|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|SIMPLE_SEGMENT|8681,8688|false|false|false|||Release
Finding|Functional Concept|SIMPLE_SEGMENT|8681,8688|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|SIMPLE_SEGMENT|8681,8688|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8681,8688|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Event|Event|SIMPLE_SEGMENT|8709,8718|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|8709,8718|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8709,8718|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8709,8718|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8709,8718|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8709,8730|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|8709,8730|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8719,8730|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|8719,8730|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|8719,8730|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|SIMPLE_SEGMENT|8732,8736|false|false|false|||Home
Finding|Idea or Concept|SIMPLE_SEGMENT|8732,8736|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|8732,8736|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|8732,8736|false|false|false|C1553498|home health encounter|Home
Event|Event|SIMPLE_SEGMENT|8739,8748|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|8739,8748|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8739,8748|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8739,8748|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8739,8748|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|8739,8758|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8749,8758|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|8749,8758|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|8749,8758|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|8749,8758|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8749,8758|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Finding|SIMPLE_SEGMENT|8760,8768|false|false|false|C0741302|atypia morphology|Atypical
Finding|Sign or Symptom|SIMPLE_SEGMENT|8760,8779|false|false|false|C0262384|Atypical chest pain|Atypical Chest Pain
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8769,8774|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|SIMPLE_SEGMENT|8769,8774|false|false|false|C0741025|Chest problem|Chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8769,8779|false|false|false|C2926613||Chest Pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|8769,8779|false|false|false|C0008031|Chest Pain|Chest Pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8775,8779|false|true|false|C2598155||Pain
Event|Event|SIMPLE_SEGMENT|8775,8779|false|false|false|||Pain
Finding|Functional Concept|SIMPLE_SEGMENT|8775,8779|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|8775,8779|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Event|Event|SIMPLE_SEGMENT|8783,8792|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|8783,8792|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8783,8792|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8783,8792|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8783,8792|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8793,8802|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8793,8802|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|8793,8802|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|8793,8802|false|false|false|C1705253|Logical Condition|Condition
Event|Event|SIMPLE_SEGMENT|8804,8809|false|false|false|||Level
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8804,8826|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|8804,8826|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|SIMPLE_SEGMENT|8813,8826|false|false|false|||Consciousness
Finding|Finding|SIMPLE_SEGMENT|8813,8826|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|8813,8826|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8828,8833|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|8828,8833|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8828,8833|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|8828,8833|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|8828,8833|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|8828,8833|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|8828,8833|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|8838,8849|false|false|false|||interactive
Finding|Functional Concept|SIMPLE_SEGMENT|8838,8849|false|false|false|C1704675|Interaction|interactive
Finding|Mental Process|SIMPLE_SEGMENT|8851,8857|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8851,8864|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|8851,8864|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8858,8864|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|8858,8864|false|false|false|C1546481|What subject filter - Status|Status
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|8866,8874|false|false|false|C0009676|Confusion|Confused
Event|Event|SIMPLE_SEGMENT|8866,8874|false|false|false|||Confused
Finding|Finding|SIMPLE_SEGMENT|8866,8874|false|false|false|C0683369;C1547301|Clouded consciousness;Precaution Code - Confused|Confused
Finding|Intellectual Product|SIMPLE_SEGMENT|8866,8874|false|false|false|C0683369;C1547301|Clouded consciousness;Precaution Code - Confused|Confused
Event|Activity|SIMPLE_SEGMENT|8888,8896|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|8888,8896|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|8888,8896|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8897,8903|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|8897,8903|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|8897,8903|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|8905,8915|false|false|false|||Ambulatory
Finding|Functional Concept|SIMPLE_SEGMENT|8905,8915|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|8905,8915|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|8905,8915|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|8905,8915|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|SIMPLE_SEGMENT|8918,8929|false|false|false|||Independent
Finding|Finding|SIMPLE_SEGMENT|8918,8929|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|SIMPLE_SEGMENT|8918,8929|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Event|Event|SIMPLE_SEGMENT|8934,8943|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|8934,8943|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8934,8943|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8934,8943|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8934,8943|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8934,8956|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|8934,8956|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|8934,8956|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8944,8956|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|8944,8956|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|8944,8956|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Event|Event|SIMPLE_SEGMENT|8972,8976|false|false|false|||came
Finding|Idea or Concept|SIMPLE_SEGMENT|8984,8992|false|false|false|C1547192|Organization unit type - Hospital|hospital
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8998,9003|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|8998,9003|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8998,9008|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|8998,9008|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9004,9008|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|9004,9008|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9004,9008|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9004,9008|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Gene or Genome|SIMPLE_SEGMENT|9019,9022|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|lab
Finding|Intellectual Product|SIMPLE_SEGMENT|9019,9022|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|lab
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9023,9029|false|false|false|C0817096|Chest|chests
Event|Event|SIMPLE_SEGMENT|9035,9038|false|false|false|||EKG
Finding|Intellectual Product|SIMPLE_SEGMENT|9035,9038|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9035,9038|false|false|false|C1623258|Electrocardiography|EKG
Event|Event|SIMPLE_SEGMENT|9051,9061|false|false|false|||reassuring
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9089,9094|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|9089,9094|false|true|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Event|Event|SIMPLE_SEGMENT|9089,9094|false|false|false|||heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|9089,9094|false|true|false|C0795691|HEART PROBLEM|heart
Event|Event|SIMPLE_SEGMENT|9096,9102|false|false|false|||attack
Finding|Finding|SIMPLE_SEGMENT|9096,9102|false|false|false|C1261512;C1304680|Attack (finding);Attack behavior|attack
Finding|Social Behavior|SIMPLE_SEGMENT|9096,9102|false|false|false|C1261512;C1304680|Attack (finding);Attack behavior|attack
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9136,9142|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|SIMPLE_SEGMENT|9136,9142|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9136,9142|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Finding|Finding|SIMPLE_SEGMENT|9136,9142|false|false|false|C0038435|Stress|stress
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9136,9147|false|false|false|C0015260;C3494508|Exercise stress test;Stress Test|stress test
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9143,9147|false|false|false|C4318744|Test - temporal region|test
Event|Event|SIMPLE_SEGMENT|9143,9147|false|false|false|||test
Finding|Functional Concept|SIMPLE_SEGMENT|9143,9147|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|SIMPLE_SEGMENT|9143,9147|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|9143,9147|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9143,9147|false|false|false|C0022885|Laboratory Procedures|test
Event|Event|SIMPLE_SEGMENT|9163,9170|false|false|false|||suggest
Event|Event|SIMPLE_SEGMENT|9175,9183|false|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|9175,9183|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|9175,9186|true|true|false|C0332120|Evidence of (contextual qualifier)|evidence of
Finding|Idea or Concept|SIMPLE_SEGMENT|9187,9196|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9197,9205|false|false|false|C0018787|Heart|coronary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9197,9212|false|false|false|C0205042|Coronary artery|coronary artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9197,9220|true|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|coronary artery disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9206,9212|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|9206,9212|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9206,9220|false|false|false|C0852949|Arteriopathic disease|artery disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9213,9220|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|9213,9220|false|false|false|||disease
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9229,9234|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|9229,9234|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9229,9239|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9229,9239|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9235,9239|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|9235,9239|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9235,9239|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9235,9239|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|9244,9256|false|false|false|||reproducible
Event|Event|SIMPLE_SEGMENT|9262,9270|false|false|false|||touching
Finding|Functional Concept|SIMPLE_SEGMENT|9262,9270|false|false|false|C2584295|Touching|touching
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9276,9281|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|9276,9281|false|false|false|C0741025|Chest problem|chest
Event|Event|SIMPLE_SEGMENT|9297,9304|false|false|false|||typical
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9308,9316|false|false|false|C0018787|Heart|coronary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9308,9323|false|false|false|C0205042|Coronary artery|coronary artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9308,9331|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|coronary artery disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9317,9323|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|9317,9323|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9317,9331|false|false|false|C0852949|Arteriopathic disease|artery disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9324,9331|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|9324,9331|false|false|false|||disease
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9332,9336|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|9332,9336|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9332,9336|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9332,9336|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|SIMPLE_SEGMENT|9344,9350|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|9344,9350|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Drug|Organic Chemical|SIMPLE_SEGMENT|9355,9362|false|false|false|C0163712|Relate - vinyl resin|related
Event|Event|SIMPLE_SEGMENT|9355,9362|false|false|false|||related
Finding|Finding|SIMPLE_SEGMENT|9355,9362|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|SIMPLE_SEGMENT|9355,9362|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9366,9381|false|false|false|C2707260||musculoskeletal
Event|Event|SIMPLE_SEGMENT|9366,9381|false|false|false|||musculoskeletal
Finding|Functional Concept|SIMPLE_SEGMENT|9366,9381|false|false|false|C0497254|Musculoskeletal|musculoskeletal
Finding|Finding|SIMPLE_SEGMENT|9366,9386|false|false|false|C0026858|Musculoskeletal Pain|musculoskeletal pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9382,9386|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|9382,9386|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|9382,9386|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|9382,9386|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|9395,9402|false|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|9395,9402|false|false|false|C0392747|Changing|changes
Event|Event|SIMPLE_SEGMENT|9413,9417|false|false|false|||made
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9426,9436|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|9426,9436|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|9426,9436|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Finding|Intellectual Product|SIMPLE_SEGMENT|9426,9441|false|false|false|C0746470|MEDICATION LIST|medication list
Event|Event|SIMPLE_SEGMENT|9437,9441|false|false|false|||list
Finding|Intellectual Product|SIMPLE_SEGMENT|9437,9441|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|SIMPLE_SEGMENT|9452,9460|false|false|false|||followup
Procedure|Health Care Activity|SIMPLE_SEGMENT|9452,9460|false|false|false|C1522577|follow-up|followup
Event|Event|SIMPLE_SEGMENT|9471,9483|false|false|false|||cardiologist
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9496,9506|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|9496,9506|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|9496,9506|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|9507,9514|false|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|9507,9514|false|false|false|C0392747|Changing|changes
Procedure|Health Care Activity|SIMPLE_SEGMENT|9518,9526|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9527,9539|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|9527,9539|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|9527,9539|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

