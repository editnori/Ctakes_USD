 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|43,52|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|43,52|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|43,57|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|77,86|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|77,86|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|77,91|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|133,136|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|144,151|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|144,151|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|SIMPLE_SEGMENT|153,165|false|false|false|||NEUROSURGERY
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|153,165|false|false|false|C0524850|Neurosurgical Procedures|NEUROSURGERY
Disorder|Injury or Poisoning|Allergies|180,191|false|false|false|C0161486;C2876539|Poisoning by penicillin;Poisoning by, adverse effect of and underdosing of penicillins|Penicillins
Drug|Antibiotic|Allergies|180,191|false|false|false|C0030842|penicillins|Penicillins
Drug|Organic Chemical|Allergies|180,191|false|false|false|C0030842|penicillins|Penicillins
Event|Event|Allergies|180,191|false|false|false|||Penicillins
Finding|Pathologic Function|Allergies|180,191|false|false|false|C0413443|Adverse reaction to penicillins|Penicillins
Event|Event|Allergies|194,203|false|false|false|||Attending
Finding|Functional Concept|Allergies|194,203|false|false|false|C1999232|Attending (action)|Attending
Finding|Functional Concept|Chief Complaint|228,232|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|Chief Complaint|228,237|false|false|false|C0230371|Structure of left hand|Left hand
Anatomy|Body Part, Organ, or Organ Component|Chief Complaint|233,237|false|false|false|C0018563;C4285005|Hand;Upper extremity>Hand|hand
Finding|Finding|Chief Complaint|233,237|false|false|false|C0741992|Hand problem|hand
Anatomy|Body Location or Region|Chief Complaint|242,246|false|false|false|C0015450;C4266571|Face;Head>Face|face
Disorder|Disease or Syndrome|Chief Complaint|242,246|false|false|false|C3160739|FANCONI ANEMIA, COMPLEMENTATION GROUP E|face
Finding|Gene or Genome|Chief Complaint|242,246|false|false|false|C1414531;C1423759;C2828055|ELOVL6 gene;FANCE gene;FANCE wt Allele|face
Finding|Sign or Symptom|Chief Complaint|242,255|false|false|false|C0239511|Numbness of face|face numbness
Event|Event|Chief Complaint|247,255|false|false|false|||numbness
Finding|Finding|Chief Complaint|247,255|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|Chief Complaint|247,255|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Functional Concept|Chief Complaint|257,261|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Chief Complaint|257,266|false|false|false|C0230371|Structure of left hand|left hand
Finding|Finding|Chief Complaint|257,275|false|false|false|C2141892|left hand weakness|left hand weakness
Anatomy|Body Part, Organ, or Organ Component|Chief Complaint|262,266|false|false|false|C0018563;C4285005|Hand;Upper extremity>Hand|hand
Finding|Finding|Chief Complaint|262,266|false|false|false|C0741992|Hand problem|hand
Finding|Finding|Chief Complaint|262,275|false|false|false|C0575810|Weakness of hand|hand weakness
Event|Event|Chief Complaint|267,275|false|false|false|||weakness
Finding|Sign or Symptom|Chief Complaint|267,275|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Event|Event|Chief Complaint|280,290|false|false|false|||clumsiness
Finding|Sign or Symptom|Chief Complaint|280,290|false|false|false|C0233844|Clumsiness|clumsiness
Event|Event|Chief Complaint|293,298|false|false|false|||fever
Finding|Finding|Chief Complaint|293,298|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|Chief Complaint|293,298|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|Chief Complaint|304,312|false|false|false|||headache
Finding|Sign or Symptom|Chief Complaint|304,312|false|false|false|C0018681|Headache|headache
Finding|Classification|Chief Complaint|316,321|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|322,330|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|322,330|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|334,352|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|343,352|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|343,352|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|343,352|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|343,352|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|343,352|false|false|false|C0184661|Interventional procedure|Procedure
Finding|Functional Concept|Chief Complaint|354,359|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Event|Event|Chief Complaint|369,379|false|false|false|||craniotomy
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|369,379|false|false|false|C0010280|Craniotomy|craniotomy
Disorder|Disease or Syndrome|Chief Complaint|384,391|false|false|false|C0000833|Abscess|abscess
Finding|Intellectual Product|Chief Complaint|384,391|false|false|false|C1546533||abscess
Anatomy|Body Location or Region|Chief Complaint|392,400|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Chief Complaint|392,400|false|false|false|C0332803|Surgical wound|incision
Event|Event|Chief Complaint|392,400|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|392,400|false|false|false|C0184898|Surgical incisions|incision
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|392,413|false|false|false|C0152277|Incision and drainage|incision and drainage
Event|Event|Chief Complaint|405,413|false|false|false|||drainage
Finding|Body Substance|Chief Complaint|405,413|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|Chief Complaint|405,413|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|405,413|false|false|false|C0013103|Drainage procedure|drainage
Event|Event|History of Present Illness|483,490|false|false|false|||history
Finding|Conceptual Entity|History of Present Illness|483,490|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|483,490|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|483,490|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|483,493|false|false|false|C0262926|Medical History|history of
Event|Event|History of Present Illness|498,506|false|false|false|||presents
Event|Event|History of Present Illness|512,521|false|false|false|||headaches
Finding|Sign or Symptom|History of Present Illness|512,521|false|false|false|C0018681|Headache|headaches
Finding|Functional Concept|History of Present Illness|526,530|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|526,535|false|false|false|C0230371|Structure of left hand|left hand
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|531,535|false|false|false|C0018563;C4285005|Hand;Upper extremity>Hand|hand
Finding|Finding|History of Present Illness|531,535|false|false|false|C0741992|Hand problem|hand
Event|Event|History of Present Illness|536,546|false|false|false|||clumsiness
Finding|Sign or Symptom|History of Present Illness|536,546|false|false|false|C0233844|Clumsiness|clumsiness
Finding|Body Substance|History of Present Illness|548,555|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|548,555|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|548,555|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|History of Present Illness|556,562|false|false|false|||states
Event|Event|History of Present Illness|573,582|false|false|false|||headaches
Finding|Sign or Symptom|History of Present Illness|573,582|false|false|false|C0018681|Headache|headaches
Event|Event|History of Present Illness|589,598|false|false|false|||presented
Finding|Intellectual Product|History of Present Illness|614,618|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|History of Present Illness|647,651|true|false|false|||much
Finding|Finding|History of Present Illness|647,651|true|false|false|C4281574|Much|much
Event|Event|History of Present Illness|678,682|false|false|false|||left
Finding|Functional Concept|History of Present Illness|678,682|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|684,688|false|false|false|C0018563;C4285005|Hand;Upper extremity>Hand|hand
Finding|Finding|History of Present Illness|684,688|false|false|false|C0741992|Hand problem|hand
Event|Event|History of Present Illness|689,699|false|false|false|||clumsiness
Finding|Sign or Symptom|History of Present Illness|689,699|false|false|false|C0233844|Clumsiness|clumsiness
Event|Event|History of Present Illness|705,711|false|false|false|||states
Event|Event|History of Present Illness|725,735|false|false|false|||difficulty
Finding|Finding|History of Present Illness|725,735|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Finding|Finding|History of Present Illness|725,740|false|false|false|C0332218|Difficult (qualifier value)|difficulty with
Finding|Organism Function|History of Present Illness|742,750|false|false|false|C0220843|grasp|grasping
Event|Event|History of Present Illness|751,758|false|false|false|||objects
Event|Event|History of Present Illness|763,768|false|false|false|||using
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|773,780|false|false|false|C0016129|Fingers|fingers
Event|Event|History of Present Illness|791,799|false|false|false|||reported
Event|Event|History of Present Illness|800,804|false|false|false|||some
Event|Event|History of Present Illness|806,814|false|false|false|||numbness
Finding|Finding|History of Present Illness|806,814|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|History of Present Illness|806,814|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|822,826|false|false|false|C0018563;C4285005|Hand;Upper extremity>Hand|hand
Finding|Finding|History of Present Illness|822,826|false|false|false|C0741992|Hand problem|hand
Event|Event|History of Present Illness|839,848|false|false|false|||presented
Event|Event|History of Present Illness|876,881|false|false|false|||found
Event|Event|History of Present Illness|892,903|false|false|false|||temperature
Procedure|Health Care Activity|History of Present Illness|892,903|false|false|false|C0886414|Body temperature measurement|temperature
Drug|Organic Chemical|History of Present Illness|932,939|false|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|History of Present Illness|932,939|false|false|false|C0699142|Tylenol|Tylenol
Event|Event|History of Present Illness|961,966|false|false|false|||after
Finding|Intellectual Product|History of Present Illness|968,972|false|false|false|C1720092|Once - dosing instruction fragment|Once
Finding|Body Substance|History of Present Illness|984,991|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|984,991|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|984,991|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|997,1001|false|false|false|||seen
Event|Event|History of Present Illness|1019,1030|false|false|false|||recommended
Event|Event|History of Present Illness|1034,1037|false|false|false|||MRI
Finding|Gene or Genome|History of Present Illness|1034,1037|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|History of Present Illness|1034,1037|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|History of Present Illness|1034,1037|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Diagnostic Procedure|History of Present Illness|1034,1042|false|false|false|C0412674|MRI of head|MRI head
Anatomy|Body Location or Region|History of Present Illness|1038,1042|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1038,1042|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|History of Present Illness|1038,1042|false|false|false|C0362076|Problems with head|head
Event|Event|History of Present Illness|1038,1042|false|false|false|||head
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1038,1042|false|false|false|C0876917|Procedure on head|head
Event|Event|History of Present Illness|1044,1047|false|false|false|||MRI
Finding|Gene or Genome|History of Present Illness|1044,1047|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|History of Present Illness|1044,1047|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|History of Present Illness|1044,1047|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Diagnostic Procedure|History of Present Illness|1044,1052|false|false|false|C0412674|MRI of head|MRI head
Anatomy|Body Location or Region|History of Present Illness|1048,1052|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1048,1052|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|History of Present Illness|1048,1052|false|false|false|C0362076|Problems with head|head
Event|Event|History of Present Illness|1048,1052|false|false|false|||head
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1048,1052|false|false|false|C0876917|Procedure on head|head
Event|Event|History of Present Illness|1053,1061|false|false|false|||revealed
Event|Event|History of Present Illness|1076,1082|false|false|false|||lesion
Finding|Finding|History of Present Illness|1076,1082|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|History of Present Illness|1076,1082|false|false|false|C0221198;C1546698|Lesion|lesion
Event|Event|History of Present Illness|1083,1093|false|false|false|||concerning
Finding|Functional Concept|History of Present Illness|1102,1112|false|false|false|C0036525;C1522484|Metastatic to;metastatic qualifier|metastatic
Disorder|Neoplastic Process|History of Present Illness|1102,1120|false|false|false|C0027627;C2939419;C2939420|Metastatic Neoplasm;Metastatic malignant neoplasm;Neoplasm Metastasis|metastatic disease
Finding|Finding|History of Present Illness|1102,1120|false|false|false|C1513183|Metastatic Lesion|metastatic disease
Disorder|Disease or Syndrome|History of Present Illness|1113,1120|false|false|false|C0012634|Disease|disease
Event|Event|History of Present Illness|1113,1120|false|false|false|||disease
Disorder|Disease or Syndrome|History of Present Illness|1126,1133|false|false|false|C0000833|Abscess|abscess
Event|Event|History of Present Illness|1126,1133|false|false|false|||abscess
Finding|Intellectual Product|History of Present Illness|1126,1133|false|false|false|C1546533||abscess
Event|Event|History of Present Illness|1135,1147|false|false|false|||Neurosurgery
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1135,1147|false|false|false|C0524850|Neurosurgical Procedures|Neurosurgery
Event|Event|History of Present Illness|1152,1161|false|false|false|||consulted
Event|Event|History of Present Illness|1174,1184|false|false|false|||evaluation
Finding|Idea or Concept|History of Present Illness|1174,1184|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|History of Present Illness|1174,1184|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Event|Event|History of Present Illness|1191,1198|false|false|false|||reports
Finding|Intellectual Product|History of Present Illness|1201,1205|false|false|false|C1547225|Mild Severity of Illness Code|mild
Event|Event|History of Present Illness|1206,1214|false|false|false|||headache
Finding|Sign or Symptom|History of Present Illness|1206,1214|false|false|false|C0018681|Headache|headache
Event|Event|History of Present Illness|1216,1224|false|false|false|||numbness
Finding|Finding|History of Present Illness|1216,1224|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|History of Present Illness|1216,1224|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Functional Concept|History of Present Illness|1232,1236|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|History of Present Illness|1232,1249|false|false|false|C0230026|Left side of face|left side of face
Anatomy|Body Location or Region|History of Present Illness|1237,1249|false|false|false|C4322912|Side of face|side of face
Anatomy|Body Location or Region|History of Present Illness|1245,1249|false|false|false|C0015450;C4266571|Face;Head>Face|face
Disorder|Disease or Syndrome|History of Present Illness|1245,1249|false|false|false|C3160739|FANCONI ANEMIA, COMPLEMENTATION GROUP E|face
Event|Event|History of Present Illness|1245,1249|false|false|false|||face
Finding|Gene or Genome|History of Present Illness|1245,1249|false|false|false|C1414531;C1423759;C2828055|ELOVL6 gene;FANCE gene;FANCE wt Allele|face
Event|Event|History of Present Illness|1255,1265|false|false|false|||difficulty
Finding|Finding|History of Present Illness|1255,1265|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Finding|Functional Concept|History of Present Illness|1276,1280|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1276,1285|false|false|false|C0230371|Structure of left hand|left hand
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1281,1285|false|false|false|C0018563;C4285005|Hand;Upper extremity>Hand|hand
Finding|Finding|History of Present Illness|1281,1285|false|false|false|C0741992|Hand problem|hand
Event|Event|History of Present Illness|1291,1297|true|false|false|||denies
Event|Event|History of Present Illness|1309,1315|true|false|false|||travel
Finding|Daily or Recreational Activity|History of Present Illness|1309,1315|true|false|false|C0040802|travel|travel
Procedure|Health Care Activity|History of Present Illness|1309,1315|true|false|false|C1555670|travel charge|travel
Event|Event|History of Present Illness|1348,1357|true|false|false|||ingesting
Event|Event|History of Present Illness|1362,1365|true|false|false|||raw
Procedure|Diagnostic Procedure|History of Present Illness|1362,1365|true|false|false|C0001884|Airway Resistance Test|raw
Event|Event|History of Present Illness|1369,1377|true|false|false|||uncooked
Drug|Food|History of Present Illness|1379,1384|true|false|false|C0025017|Meat|meats
Event|Event|History of Present Illness|1379,1384|true|false|false|||meats
Event|Event|History of Present Illness|1395,1401|true|false|false|||denies
Event|Event|History of Present Illness|1406,1413|true|false|false|||changes
Finding|Functional Concept|History of Present Illness|1406,1413|true|false|false|C0392747|Changing|changes
Attribute|Clinical Attribute|History of Present Illness|1417,1423|true|false|false|C2707266||vision
Event|Event|History of Present Illness|1417,1423|true|false|false|||vision
Finding|Organism Function|History of Present Illness|1417,1423|true|false|false|C0042789|Vision|vision
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|1425,1435|true|false|false|C0013362|Dysarthria|dysarthria
Event|Event|History of Present Illness|1425,1435|true|false|false|||dysarthria
Event|Event|History of Present Illness|1438,1446|false|false|false|||weakness
Finding|Sign or Symptom|History of Present Illness|1438,1446|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Attribute|Clinical Attribute|History of Present Illness|1448,1454|false|false|false|C4255480||nausea
Event|Event|History of Present Illness|1448,1454|false|false|false|||nausea
Finding|Sign or Symptom|History of Present Illness|1448,1454|false|false|false|C0027497|Nausea|nausea
Event|Event|History of Present Illness|1456,1465|false|false|false|||vomitting
Event|Event|History of Present Illness|1467,1475|false|false|false|||diarrhea
Finding|Finding|History of Present Illness|1467,1475|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|History of Present Illness|1467,1475|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Drug|Organic Chemical|History of Present Illness|1477,1482|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|1477,1482|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|History of Present Illness|1477,1482|false|false|false|||cough
Finding|Sign or Symptom|History of Present Illness|1477,1482|false|false|false|C0010200|Coughing|cough
Event|Event|History of Present Illness|1487,1493|false|false|false|||chills
Finding|Sign or Symptom|History of Present Illness|1487,1493|true|false|false|C0085593|Chills|chills
Disorder|Disease or Syndrome|Past Medical History|1520,1538|false|false|false|C0026769|Multiple Sclerosis|Multiple sclerosis
Event|Event|Past Medical History|1529,1538|false|false|false|||sclerosis
Finding|Pathologic Function|Past Medical History|1529,1538|false|false|false|C0036429|Sclerosis|sclerosis
Event|Event|Family Medical History|1577,1583|false|false|false|||Mother
Finding|Idea or Concept|Family Medical History|1577,1583|false|false|false|C1546508|Relationship - Mother|Mother
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1589,1599|false|false|false|C0030274|Pancreas|pancreatic
Drug|Amino Acid, Peptide, or Protein|Family Medical History|1589,1599|false|false|false|C0030292|Pancreatic Hormones|pancreatic
Drug|Hormone|Family Medical History|1589,1599|false|false|false|C0030292|Pancreatic Hormones|pancreatic
Drug|Pharmacologic Substance|Family Medical History|1589,1599|false|false|false|C0030292|Pancreatic Hormones|pancreatic
Disorder|Neoplastic Process|Family Medical History|1589,1606|false|false|false|C0235974;C0346647|Malignant neoplasm of pancreas;Pancreatic carcinoma|pancreatic cancer
Disorder|Neoplastic Process|Family Medical History|1600,1606|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Family Medical History|1600,1606|false|false|false|||cancer
Finding|Conceptual Entity|Family Medical History|1608,1615|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|brother
Finding|Idea or Concept|Family Medical History|1608,1615|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|brother
Anatomy|Body Location or Region|Family Medical History|1616,1620|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1616,1620|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Family Medical History|1616,1620|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Family Medical History|1616,1620|false|false|false|C0740941|Lung Problem|lung
Disorder|Neoplastic Process|Family Medical History|1616,1627|false|false|false|C0242379;C0684249|Carcinoma of lung;Malignant neoplasm of lung|lung cancer
Disorder|Neoplastic Process|Family Medical History|1621,1627|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Family Medical History|1621,1627|false|false|false|||cancer
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1647,1652|false|false|false|C0006104;C4266577|Brain;Head>Brain|brain
Disorder|Disease or Syndrome|Family Medical History|1647,1652|false|false|false|C0006111|Brain Diseases|brain
Disorder|Neoplastic Process|Family Medical History|1647,1659|false|false|false|C0006118;C0153633|Brain Neoplasms;Malignant neoplasm of brain|brain cancer
Disorder|Neoplastic Process|Family Medical History|1653,1659|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Family Medical History|1653,1659|false|false|false|||cancer
Event|Event|General Exam|1679,1687|false|false|false|||PHYSICAL
Finding|Finding|General Exam|1679,1687|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|General Exam|1679,1687|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|General Exam|1679,1687|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|General Exam|1679,1692|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|General Exam|1679,1692|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Event|Event|General Exam|1688,1692|false|false|false|||EXAM
Finding|Functional Concept|General Exam|1688,1692|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|1688,1692|false|false|false|C0582103|Medical Examination|EXAM
Procedure|Health Care Activity|General Exam|1696,1705|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|General Exam|1762,1765|false|false|false|||Gen
Finding|Classification|General Exam|1762,1765|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Finding|Gene or Genome|General Exam|1762,1765|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Event|Event|General Exam|1774,1785|false|false|false|||comfortable
Finding|Finding|General Exam|1774,1785|false|false|false|C5546696|Feeling comfortable|comfortable
Disorder|Disease or Syndrome|General Exam|1787,1790|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|1787,1790|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|1787,1790|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|1787,1790|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|1787,1790|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|General Exam|1787,1790|false|false|false|||NAD
Finding|Finding|General Exam|1787,1790|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|General Exam|1792,1797|false|false|false|C1512338|HEENT|HEENT
Event|Event|General Exam|1799,1809|false|false|false|||atraumatic
Event|Event|General Exam|1811,1824|false|false|false|||normocephalic
Anatomy|Body Part, Organ, or Organ Component|General Exam|1825,1831|false|false|false|C0034121|Pupil|Pupils
Event|Event|General Exam|1859,1863|false|false|false|||EOMs
Finding|Functional Concept|General Exam|1859,1863|false|false|false|C0241886|Extraocular|EOMs
Event|Event|General Exam|1865,1871|false|false|false|||intact
Finding|Finding|General Exam|1865,1871|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Mental Process|General Exam|1880,1886|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|General Exam|1880,1893|false|false|false|C0488568;C0488569||Mental status
Finding|Finding|General Exam|1880,1893|false|false|false|C0278060|Mental state|Mental status
Attribute|Clinical Attribute|General Exam|1887,1893|false|false|false|C5889824||status
Event|Event|General Exam|1887,1893|false|false|false|||status
Finding|Idea or Concept|General Exam|1887,1893|false|false|false|C1546481|What subject filter - Status|status
Event|Event|General Exam|1895,1900|false|false|false|||Awake
Attribute|Clinical Attribute|General Exam|1905,1910|false|false|false|C5890168||alert
Drug|Organic Chemical|General Exam|1905,1910|false|false|false|C0718338|Alert brand of caffeine|alert
Drug|Pharmacologic Substance|General Exam|1905,1910|false|false|false|C0718338|Alert brand of caffeine|alert
Event|Event|General Exam|1905,1910|false|false|false|||alert
Finding|Finding|General Exam|1905,1910|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Functional Concept|General Exam|1905,1910|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Intellectual Product|General Exam|1905,1910|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Event|Event|General Exam|1912,1923|false|false|false|||cooperative
Event|Event|General Exam|1929,1933|false|false|false|||exam
Finding|Functional Concept|General Exam|1929,1933|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|General Exam|1929,1933|false|false|false|C0582103|Medical Examination|exam
Event|Event|General Exam|1935,1941|false|false|false|||normal
Event|Event|General Exam|1942,1948|false|false|false|||affect
Finding|Mental Process|General Exam|1942,1948|false|false|false|C0001721|Affect (mental function)|affect
Procedure|Health Care Activity|General Exam|1942,1948|false|false|false|C2237113|assessment of affect|affect
Event|Event|General Exam|1950,1961|false|false|false|||Orientation
Finding|Mental Process|General Exam|1950,1961|false|false|false|C0029266|Mental Orientation|Orientation
Event|Event|General Exam|1963,1971|false|false|false|||Oriented
Finding|Finding|General Exam|1963,1971|false|false|false|C1961028|Oriented to place|Oriented
Finding|Finding|General Exam|1963,1981|false|false|false|C1961030|Oriented to person|Oriented to person
Attribute|Clinical Attribute|General Exam|1975,1981|false|false|false|C5890614||person
Event|Event|General Exam|1975,1981|false|false|false|||person
Finding|Intellectual Product|General Exam|1975,1981|false|false|false|C1522390|Person Info|person
Event|Activity|General Exam|1983,1988|false|false|false|C1882509|put - instruction imperative|place
Event|Event|General Exam|1983,1988|false|false|false|||place
Finding|Functional Concept|General Exam|1983,1988|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|General Exam|1983,1988|false|false|false|C1533810||place
Event|Event|General Exam|2000,2006|false|false|false|||Recall
Event|Governmental or Regulatory Activity|General Exam|2000,2006|false|false|false|C1705180|Recall (activity)|Recall
Finding|Mental Process|General Exam|2000,2006|false|false|false|C0034770|Mental Recall|Recall
Event|Event|General Exam|2012,2019|false|false|false|||objects
Procedure|Therapeutic or Preventive Procedure|General Exam|2023,2032|false|false|false|C0886384|5 minutes Office visit|5 minutes
Event|Event|General Exam|2025,2032|false|false|false|||minutes
Attribute|Clinical Attribute|General Exam|2034,2042|false|false|false|C2706915||Language
Event|Event|General Exam|2034,2042|false|false|false|||Language
Finding|Intellectual Product|General Exam|2034,2042|false|false|false|C0033348|Programming Languages|Language
Event|Event|General Exam|2044,2050|false|false|false|||Speech
Finding|Organism Function|General Exam|2044,2050|false|false|false|C0037817|Speech|Speech
Procedure|Diagnostic Procedure|General Exam|2044,2050|false|false|false|C0846595|Speech assessment|Speech
Finding|Idea or Concept|General Exam|2063,2067|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Event|Event|General Exam|2068,2081|false|false|false|||comprehension
Finding|Mental Process|General Exam|2068,2081|false|false|false|C0162340|Comprehension|comprehension
Event|Event|General Exam|2086,2096|false|false|false|||repetition
Finding|Finding|General Exam|2086,2096|false|false|false|C0205341;C2018025|Repeat;speech fluency repetition (physical finding)|repetition
Finding|Functional Concept|General Exam|2086,2096|false|false|false|C0205341;C2018025|Repeat;speech fluency repetition (physical finding)|repetition
Event|Event|General Exam|2098,2104|false|false|false|||Naming
Finding|Mental Process|General Exam|2098,2104|false|false|false|C0233735|Naming (function)|Naming
Event|Event|General Exam|2105,2111|false|false|false|||intact
Finding|Finding|General Exam|2105,2111|false|false|false|C1554187|Gender Status - Intact|intact
Disorder|Mental or Behavioral Dysfunction|General Exam|2116,2126|true|false|false|C0013362|Dysarthria|dysarthria
Event|Event|General Exam|2116,2126|true|false|false|||dysarthria
Event|Event|General Exam|2141,2147|true|false|false|||errors
Anatomy|Body Part, Organ, or Organ Component|General Exam|2150,2157|false|false|false|C0037303|Bone structure of cranium|Cranial
Anatomy|Body Part, Organ, or Organ Component|General Exam|2150,2164|false|false|false|C0010268|Cranial Nerves|Cranial Nerves
Disorder|Neoplastic Process|General Exam|2150,2164|false|false|false|C0004992;C0496937|Benign neoplasm of cranial nerves;Neoplasm of uncertain or unknown behavior of cranial nerves|Cranial Nerves
Anatomy|Body Part, Organ, or Organ Component|General Exam|2158,2164|false|false|false|C0027740|Nerve|Nerves
Event|Event|General Exam|2173,2179|true|false|false|||tested
Anatomy|Body Part, Organ, or Organ Component|General Exam|2184,2190|false|false|false|C0034121|Pupil|Pupils
Event|Event|General Exam|2199,2204|false|false|false|||round
Event|Event|General Exam|2209,2217|false|false|false|||reactive
Procedure|Therapeutic or Preventive Procedure|General Exam|2209,2217|false|false|false|C4722408|Reactive Therapy|reactive
Finding|Finding|General Exam|2209,2226|false|false|false|C4068744|Reactive to light|reactive to light
Drug|Amino Acid, Peptide, or Protein|General Exam|2221,2226|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|General Exam|2221,2226|false|false|false|C1570446|TNFSF14 protein, human|light
Event|Event|General Exam|2221,2226|false|false|false|||light
Finding|Finding|General Exam|2221,2226|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|General Exam|2221,2226|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|General Exam|2221,2226|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|General Exam|2221,2226|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|General Exam|2221,2226|false|false|false|C0031765|Phototherapy|light
Finding|Functional Concept|General Exam|2251,2257|false|false|false|C0234621|Visual|Visual
Event|Event|General Exam|2258,2264|false|false|false|||fields
Event|Event|General Exam|2269,2273|false|false|false|||full
Event|Event|General Exam|2277,2290|false|false|false|||confrontation
Finding|Finding|General Exam|2277,2290|false|false|false|C0518608|Social confrontation skill|confrontation
Procedure|Diagnostic Procedure|General Exam|2277,2290|false|false|false|C0700282;C1444674|Confrontation;Confrontation visual field test|confrontation
Procedure|Therapeutic or Preventive Procedure|General Exam|2277,2290|false|false|false|C0700282;C1444674|Confrontation;Confrontation visual field test|confrontation
Finding|Functional Concept|General Exam|2305,2316|true|false|false|C0241886|Extraocular|Extraocular
Procedure|Diagnostic Procedure|General Exam|2305,2326|true|false|false|C2228439|examination of extraocular movements|Extraocular movements
Event|Event|General Exam|2317,2326|true|false|false|||movements
Finding|Organism Function|General Exam|2317,2326|true|false|false|C0026649|Movement|movements
Event|Event|General Exam|2327,2333|true|false|false|||intact
Finding|Finding|General Exam|2327,2333|true|false|false|C1554187|Gender Status - Intact|intact
Disorder|Disease or Syndrome|General Exam|2354,2363|true|false|false|C0028738|Nystagmus|nystagmus
Event|Event|General Exam|2354,2363|true|false|false|||nystagmus
Anatomy|Body Part, Organ, or Organ Component|General Exam|2368,2371|false|false|false|C2338708;C3496273;C3496274|Lamina VII of gray matter of spinal cord;layer VII (Cajal);lobule VII|VII
Finding|Intellectual Product|General Exam|2368,2371|false|false|false|C0445385|Roman numeral VII|VII
Anatomy|Body Location or Region|General Exam|2373,2379|false|false|false|C0015450|Face|Facial
Event|Event|General Exam|2380,2388|false|false|false|||strength
Finding|Idea or Concept|General Exam|2380,2388|false|false|false|C0808080|Strength (attribute)|strength
Event|Event|General Exam|2393,2402|false|false|false|||sensation
Finding|Finding|General Exam|2393,2402|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|General Exam|2393,2402|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|General Exam|2393,2402|false|false|false|C2229507|sensory exam|sensation
Event|Event|General Exam|2403,2409|false|false|false|||intact
Finding|Finding|General Exam|2403,2409|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|General Exam|2414,2423|false|false|false|||symmetric
Finding|Conceptual Entity|General Exam|2414,2423|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|General Exam|2414,2423|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Anatomy|Body Part, Organ, or Organ Component|General Exam|2425,2429|false|false|false|C0228488;C2327388|Cerebellar pyramis;Lamina VIII of gray matter of spinal cord|VIII
Finding|Gene or Genome|General Exam|2425,2429|false|false|false|C0445599;C1413661|COX8A gene;Roman numeral VIII|VIII
Finding|Intellectual Product|General Exam|2425,2429|false|false|false|C0445599;C1413661|COX8A gene;Roman numeral VIII|VIII
Event|Event|General Exam|2431,2438|false|false|false|||Hearing
Finding|Finding|General Exam|2431,2438|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|Hearing
Finding|Physiologic Function|General Exam|2431,2438|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|Hearing
Event|Event|General Exam|2439,2445|false|false|false|||intact
Finding|Finding|General Exam|2439,2445|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|General Exam|2449,2454|false|false|false|||voice
Finding|Idea or Concept|General Exam|2449,2454|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Intellectual Product|General Exam|2449,2454|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Organism Function|General Exam|2449,2454|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Anatomy|Body Part, Organ, or Organ Component|General Exam|2463,2470|false|false|false|C0700374|Palate|Palatal
Event|Event|General Exam|2471,2480|false|false|false|||elevation
Procedure|Therapeutic or Preventive Procedure|General Exam|2471,2480|false|false|false|C0439775|Elevation procedure|elevation
Event|Event|General Exam|2481,2492|false|false|false|||symmetrical
Finding|Finding|General Exam|2481,2492|false|false|false|C0332516|Symmetrical|symmetrical
Anatomy|Body Part, Organ, or Organ Component|General Exam|2498,2517|false|false|false|C0224153|Structure of sternocleidomastoid muscle|Sternocleidomastoid
Anatomy|Body Part, Organ, or Organ Component|General Exam|2522,2531|false|false|false|C0224361|Structure of trapezius muscle|trapezius
Event|Event|General Exam|2532,2538|false|false|false|||normal
Anatomy|Body Part, Organ, or Organ Component|General Exam|2557,2563|true|false|false|C0040408|Tongue|Tongue
Disorder|Neoplastic Process|General Exam|2557,2563|true|false|false|C0153933|Benign neoplasm of tongue|Tongue
Procedure|Health Care Activity|General Exam|2557,2563|true|false|false|C0872394|Procedure on tongue|Tongue
Finding|Finding|General Exam|2557,2571|true|false|false|C3693372|tongue midline|Tongue midline
Anatomy|Cell Component|General Exam|2564,2571|true|false|false|C1660780|midline cell component|midline
Event|Event|General Exam|2580,2594|true|false|false|||fasciculations
Finding|Sign or Symptom|General Exam|2580,2594|true|false|false|C0015644|Muscular fasciculation|fasciculations
Event|Event|General Exam|2597,2602|false|false|false|||Motor
Finding|Functional Concept|General Exam|2597,2602|false|false|false|C1513492|motor movement|Motor
Drug|Biomedical or Dental Material|General Exam|2611,2615|false|false|false|C0012173;C1337615|Bulk (conceptual);Dietary Fiber|bulk
Drug|Food|General Exam|2611,2615|false|false|false|C0012173;C1337615|Bulk (conceptual);Dietary Fiber|bulk
Event|Event|General Exam|2611,2615|false|false|false|||bulk
Event|Event|General Exam|2620,2624|false|false|false|||tone
Finding|Finding|General Exam|2641,2649|true|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Finding|Idea or Concept|General Exam|2641,2649|true|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Disorder|Disease or Syndrome|General Exam|2641,2659|true|false|false|C0013384|Dyskinetic syndrome|abnormal movements
Finding|Finding|General Exam|2641,2659|true|false|false|C0558189|Abnormal movement|abnormal movements
Event|Event|General Exam|2650,2659|true|false|false|||movements
Finding|Organism Function|General Exam|2650,2659|true|false|false|C0026649|Movement|movements
Event|Event|General Exam|2661,2668|true|false|false|||tremors
Finding|Sign or Symptom|General Exam|2661,2668|true|false|false|C0040822|Tremor|tremors
Event|Event|General Exam|2670,2678|false|false|false|||Strength
Finding|Idea or Concept|General Exam|2670,2678|false|false|false|C0808080|Strength (attribute)|Strength
Event|Event|General Exam|2704,2709|false|false|false|||power
Finding|Social Behavior|General Exam|2704,2709|false|false|false|C0032863|Power (Psychology)|power
Finding|Pathologic Function|General Exam|2730,2744|true|false|false|C1504476|Pronator drift|pronator drift
Event|Event|General Exam|2739,2744|true|false|false|||drift
Event|Event|General Exam|2746,2755|true|false|false|||Sensation
Finding|Finding|General Exam|2746,2755|true|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Finding|Organ or Tissue Function|General Exam|2746,2755|true|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Procedure|Health Care Activity|General Exam|2746,2755|true|false|false|C2229507|sensory exam|Sensation
Event|Event|General Exam|2757,2763|false|false|false|||Intact
Finding|Finding|General Exam|2757,2763|false|false|false|C1554187|Gender Status - Intact|Intact
Drug|Amino Acid, Peptide, or Protein|General Exam|2767,2772|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|General Exam|2767,2772|false|false|false|C1570446|TNFSF14 protein, human|light
Event|Event|General Exam|2767,2772|false|false|false|||light
Finding|Finding|General Exam|2767,2772|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|General Exam|2767,2772|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|General Exam|2767,2772|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|General Exam|2767,2772|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|General Exam|2767,2772|false|false|false|C0031765|Phototherapy|light
Finding|Physiologic Function|General Exam|2767,2778|false|false|false|C0423553|Light touch|light touch
Event|Event|General Exam|2773,2778|false|false|false|||touch
Finding|Mental Process|General Exam|2773,2778|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Finding|Organ or Tissue Function|General Exam|2773,2778|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Procedure|Therapeutic or Preventive Procedure|General Exam|2773,2778|false|false|false|C0152054|Therapeutic Touch|touch
Event|Event|General Exam|2780,2788|false|false|false|||PHYSICAL
Finding|Finding|General Exam|2780,2788|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|General Exam|2780,2788|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|General Exam|2780,2788|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|General Exam|2780,2793|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|General Exam|2780,2793|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Event|Event|General Exam|2789,2793|false|false|false|||EXAM
Finding|Functional Concept|General Exam|2789,2793|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|2789,2793|false|false|false|C0582103|Medical Examination|EXAM
Event|Event|General Exam|2797,2806|false|false|false|||DISCHARGE
Finding|Body Substance|General Exam|2797,2806|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|2797,2806|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|2797,2806|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|2797,2806|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|General Exam|2857,2860|false|false|false|||Gen
Finding|Classification|General Exam|2857,2860|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Finding|Gene or Genome|General Exam|2857,2860|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Event|Event|General Exam|2869,2880|false|false|false|||comfortable
Finding|Finding|General Exam|2869,2880|false|false|false|C5546696|Feeling comfortable|comfortable
Disorder|Disease or Syndrome|General Exam|2882,2885|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|2882,2885|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|2882,2885|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|2882,2885|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|2882,2885|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|General Exam|2882,2885|false|false|false|||NAD
Finding|Finding|General Exam|2882,2885|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|General Exam|2887,2892|false|false|false|C1512338|HEENT|HEENT
Event|Event|General Exam|2894,2904|false|false|false|||atraumatic
Event|Event|General Exam|2906,2919|false|false|false|||normocephalic
Finding|Functional Concept|General Exam|2926,2931|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Event|Event|General Exam|2932,2942|false|false|false|||craniotomy
Procedure|Therapeutic or Preventive Procedure|General Exam|2932,2942|false|false|false|C0010280|Craniotomy|craniotomy
Anatomy|Body Location or Region|General Exam|2944,2952|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|General Exam|2944,2952|false|false|false|C0332803|Surgical wound|incision
Event|Event|General Exam|2944,2952|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|General Exam|2944,2952|false|false|false|C0184898|Surgical incisions|incision
Anatomy|Body Part, Organ, or Organ Component|General Exam|2954,2960|false|false|false|C0034121|Pupil|Pupils
Event|Event|General Exam|2981,2985|false|false|false|||EOMs
Finding|Functional Concept|General Exam|2981,2985|false|false|false|C0241886|Extraocular|EOMs
Event|Event|General Exam|2987,2993|false|false|false|||intact
Finding|Finding|General Exam|2987,2993|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Mental Process|General Exam|3002,3008|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|General Exam|3002,3015|false|false|false|C0488568;C0488569||Mental status
Finding|Finding|General Exam|3002,3015|false|false|false|C0278060|Mental state|Mental status
Attribute|Clinical Attribute|General Exam|3009,3015|false|false|false|C5889824||status
Event|Event|General Exam|3009,3015|false|false|false|||status
Finding|Idea or Concept|General Exam|3009,3015|false|false|false|C1546481|What subject filter - Status|status
Event|Event|General Exam|3017,3022|false|false|false|||Awake
Attribute|Clinical Attribute|General Exam|3027,3032|false|false|false|C5890168||alert
Drug|Organic Chemical|General Exam|3027,3032|false|false|false|C0718338|Alert brand of caffeine|alert
Drug|Pharmacologic Substance|General Exam|3027,3032|false|false|false|C0718338|Alert brand of caffeine|alert
Event|Event|General Exam|3027,3032|false|false|false|||alert
Finding|Finding|General Exam|3027,3032|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Functional Concept|General Exam|3027,3032|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Intellectual Product|General Exam|3027,3032|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Event|Event|General Exam|3034,3045|false|false|false|||cooperative
Event|Event|General Exam|3051,3055|false|false|false|||exam
Finding|Functional Concept|General Exam|3051,3055|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|General Exam|3051,3055|false|false|false|C0582103|Medical Examination|exam
Event|Event|General Exam|3057,3063|false|false|false|||normal
Event|Event|General Exam|3064,3070|false|false|false|||affect
Finding|Mental Process|General Exam|3064,3070|false|false|false|C0001721|Affect (mental function)|affect
Procedure|Health Care Activity|General Exam|3064,3070|false|false|false|C2237113|assessment of affect|affect
Event|Event|General Exam|3072,3083|false|false|false|||Orientation
Finding|Mental Process|General Exam|3072,3083|false|false|false|C0029266|Mental Orientation|Orientation
Event|Event|General Exam|3085,3093|false|false|false|||Oriented
Finding|Finding|General Exam|3085,3093|false|false|false|C1961028|Oriented to place|Oriented
Finding|Finding|General Exam|3085,3103|false|false|false|C1961030|Oriented to person|Oriented to person
Attribute|Clinical Attribute|General Exam|3097,3103|false|false|false|C5890614||person
Event|Event|General Exam|3097,3103|false|false|false|||person
Finding|Intellectual Product|General Exam|3097,3103|false|false|false|C1522390|Person Info|person
Event|Activity|General Exam|3105,3110|false|false|false|C1882509|put - instruction imperative|place
Event|Event|General Exam|3105,3110|false|false|false|||place
Finding|Functional Concept|General Exam|3105,3110|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|General Exam|3105,3110|false|false|false|C1533810||place
Event|Event|General Exam|3122,3128|false|false|false|||Recall
Event|Governmental or Regulatory Activity|General Exam|3122,3128|false|false|false|C1705180|Recall (activity)|Recall
Finding|Mental Process|General Exam|3122,3128|false|false|false|C0034770|Mental Recall|Recall
Event|Event|General Exam|3134,3141|false|false|false|||objects
Procedure|Therapeutic or Preventive Procedure|General Exam|3145,3154|false|false|false|C0886384|5 minutes Office visit|5 minutes
Event|Event|General Exam|3147,3154|false|false|false|||minutes
Attribute|Clinical Attribute|General Exam|3156,3164|false|false|false|C2706915||Language
Event|Event|General Exam|3156,3164|false|false|false|||Language
Finding|Intellectual Product|General Exam|3156,3164|false|false|false|C0033348|Programming Languages|Language
Event|Event|General Exam|3166,3172|false|false|false|||Speech
Finding|Organism Function|General Exam|3166,3172|false|false|false|C0037817|Speech|Speech
Procedure|Diagnostic Procedure|General Exam|3166,3172|false|false|false|C0846595|Speech assessment|Speech
Finding|Idea or Concept|General Exam|3185,3189|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Event|Event|General Exam|3190,3203|false|false|false|||comprehension
Finding|Mental Process|General Exam|3190,3203|false|false|false|C0162340|Comprehension|comprehension
Event|Event|General Exam|3208,3218|false|false|false|||repetition
Finding|Finding|General Exam|3208,3218|false|false|false|C0205341;C2018025|Repeat;speech fluency repetition (physical finding)|repetition
Finding|Functional Concept|General Exam|3208,3218|false|false|false|C0205341;C2018025|Repeat;speech fluency repetition (physical finding)|repetition
Event|Event|General Exam|3220,3226|false|false|false|||Naming
Finding|Mental Process|General Exam|3220,3226|false|false|false|C0233735|Naming (function)|Naming
Event|Event|General Exam|3227,3233|false|false|false|||intact
Finding|Finding|General Exam|3227,3233|false|false|false|C1554187|Gender Status - Intact|intact
Disorder|Mental or Behavioral Dysfunction|General Exam|3238,3248|true|false|false|C0013362|Dysarthria|dysarthria
Event|Event|General Exam|3238,3248|true|false|false|||dysarthria
Event|Event|General Exam|3263,3269|true|false|false|||errors
Anatomy|Body Part, Organ, or Organ Component|General Exam|3272,3279|false|false|false|C0037303|Bone structure of cranium|Cranial
Anatomy|Body Part, Organ, or Organ Component|General Exam|3272,3286|false|false|false|C0010268|Cranial Nerves|Cranial Nerves
Disorder|Neoplastic Process|General Exam|3272,3286|false|false|false|C0004992;C0496937|Benign neoplasm of cranial nerves;Neoplasm of uncertain or unknown behavior of cranial nerves|Cranial Nerves
Anatomy|Body Part, Organ, or Organ Component|General Exam|3280,3286|false|false|false|C0027740|Nerve|Nerves
Event|Event|General Exam|3295,3301|true|false|false|||tested
Anatomy|Body Part, Organ, or Organ Component|General Exam|3306,3312|false|false|false|C0034121|Pupil|Pupils
Event|Event|General Exam|3321,3326|false|false|false|||round
Event|Event|General Exam|3331,3339|false|false|false|||reactive
Procedure|Therapeutic or Preventive Procedure|General Exam|3331,3339|false|false|false|C4722408|Reactive Therapy|reactive
Finding|Finding|General Exam|3331,3348|false|false|false|C4068744|Reactive to light|reactive to light
Drug|Amino Acid, Peptide, or Protein|General Exam|3343,3348|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|General Exam|3343,3348|false|false|false|C1570446|TNFSF14 protein, human|light
Event|Event|General Exam|3343,3348|false|false|false|||light
Finding|Finding|General Exam|3343,3348|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|General Exam|3343,3348|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|General Exam|3343,3348|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|General Exam|3343,3348|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|General Exam|3343,3348|false|false|false|C0031765|Phototherapy|light
Finding|Functional Concept|General Exam|3374,3380|false|false|false|C0234621|Visual|Visual
Event|Event|General Exam|3381,3387|false|false|false|||fields
Event|Event|General Exam|3392,3396|false|false|false|||full
Event|Event|General Exam|3400,3413|false|false|false|||confrontation
Finding|Finding|General Exam|3400,3413|false|false|false|C0518608|Social confrontation skill|confrontation
Procedure|Diagnostic Procedure|General Exam|3400,3413|false|false|false|C0700282;C1444674|Confrontation;Confrontation visual field test|confrontation
Procedure|Therapeutic or Preventive Procedure|General Exam|3400,3413|false|false|false|C0700282;C1444674|Confrontation;Confrontation visual field test|confrontation
Finding|Functional Concept|General Exam|3428,3439|true|false|false|C0241886|Extraocular|Extraocular
Procedure|Diagnostic Procedure|General Exam|3428,3449|true|false|false|C2228439|examination of extraocular movements|Extraocular movements
Event|Event|General Exam|3440,3449|true|false|false|||movements
Finding|Organism Function|General Exam|3440,3449|true|false|false|C0026649|Movement|movements
Event|Event|General Exam|3450,3456|true|false|false|||intact
Finding|Finding|General Exam|3450,3456|true|false|false|C1554187|Gender Status - Intact|intact
Disorder|Disease or Syndrome|General Exam|3477,3486|true|false|false|C0028738|Nystagmus|nystagmus
Event|Event|General Exam|3477,3486|true|false|false|||nystagmus
Anatomy|Body Part, Organ, or Organ Component|General Exam|3491,3494|false|false|false|C2338708;C3496273;C3496274|Lamina VII of gray matter of spinal cord;layer VII (Cajal);lobule VII|VII
Finding|Intellectual Product|General Exam|3491,3494|false|false|false|C0445385|Roman numeral VII|VII
Anatomy|Body Location or Region|General Exam|3496,3502|false|false|false|C0015450|Face|Facial
Event|Event|General Exam|3503,3511|false|false|false|||strength
Finding|Idea or Concept|General Exam|3503,3511|false|false|false|C0808080|Strength (attribute)|strength
Event|Event|General Exam|3516,3525|false|false|false|||sensation
Finding|Finding|General Exam|3516,3525|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|General Exam|3516,3525|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|General Exam|3516,3525|false|false|false|C2229507|sensory exam|sensation
Event|Event|General Exam|3526,3532|false|false|false|||intact
Finding|Finding|General Exam|3526,3532|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|General Exam|3537,3546|false|false|false|||symmetric
Finding|Conceptual Entity|General Exam|3537,3546|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|General Exam|3537,3546|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Anatomy|Body Part, Organ, or Organ Component|General Exam|3548,3552|false|false|false|C0228488;C2327388|Cerebellar pyramis;Lamina VIII of gray matter of spinal cord|VIII
Finding|Gene or Genome|General Exam|3548,3552|false|false|false|C0445599;C1413661|COX8A gene;Roman numeral VIII|VIII
Finding|Intellectual Product|General Exam|3548,3552|false|false|false|C0445599;C1413661|COX8A gene;Roman numeral VIII|VIII
Event|Event|General Exam|3554,3561|false|false|false|||Hearing
Finding|Finding|General Exam|3554,3561|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|Hearing
Finding|Physiologic Function|General Exam|3554,3561|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|Hearing
Event|Event|General Exam|3562,3568|false|false|false|||intact
Finding|Finding|General Exam|3562,3568|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|General Exam|3572,3577|false|false|false|||voice
Finding|Idea or Concept|General Exam|3572,3577|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Intellectual Product|General Exam|3572,3577|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Organism Function|General Exam|3572,3577|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Anatomy|Body Part, Organ, or Organ Component|General Exam|3586,3593|false|false|false|C0700374|Palate|Palatal
Event|Event|General Exam|3594,3603|false|false|false|||elevation
Procedure|Therapeutic or Preventive Procedure|General Exam|3594,3603|false|false|false|C0439775|Elevation procedure|elevation
Event|Event|General Exam|3604,3615|false|false|false|||symmetrical
Finding|Finding|General Exam|3604,3615|false|false|false|C0332516|Symmetrical|symmetrical
Anatomy|Body Part, Organ, or Organ Component|General Exam|3621,3640|false|false|false|C0224153|Structure of sternocleidomastoid muscle|Sternocleidomastoid
Anatomy|Body Part, Organ, or Organ Component|General Exam|3645,3654|false|false|false|C0224361|Structure of trapezius muscle|trapezius
Event|Event|General Exam|3655,3661|false|false|false|||normal
Anatomy|Body Part, Organ, or Organ Component|General Exam|3680,3686|true|false|false|C0040408|Tongue|Tongue
Disorder|Neoplastic Process|General Exam|3680,3686|true|false|false|C0153933|Benign neoplasm of tongue|Tongue
Procedure|Health Care Activity|General Exam|3680,3686|true|false|false|C0872394|Procedure on tongue|Tongue
Finding|Finding|General Exam|3680,3694|true|false|false|C3693372|tongue midline|Tongue midline
Anatomy|Cell Component|General Exam|3687,3694|true|false|false|C1660780|midline cell component|midline
Event|Event|General Exam|3703,3717|true|false|false|||fasciculations
Finding|Sign or Symptom|General Exam|3703,3717|true|false|false|C0015644|Muscular fasciculation|fasciculations
Event|Event|General Exam|3720,3725|false|false|false|||Motor
Finding|Functional Concept|General Exam|3720,3725|false|false|false|C1513492|motor movement|Motor
Drug|Biomedical or Dental Material|General Exam|3734,3738|false|false|false|C0012173;C1337615|Bulk (conceptual);Dietary Fiber|bulk
Drug|Food|General Exam|3734,3738|false|false|false|C0012173;C1337615|Bulk (conceptual);Dietary Fiber|bulk
Event|Event|General Exam|3734,3738|false|false|false|||bulk
Event|Event|General Exam|3743,3747|false|false|false|||tone
Event|Event|General Exam|3764,3772|true|false|false|||abnormal
Finding|Finding|General Exam|3764,3772|true|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Finding|Idea or Concept|General Exam|3764,3772|true|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Event|Event|General Exam|3774,3783|true|false|false|||movements
Finding|Organism Function|General Exam|3774,3783|true|false|false|C0026649|Movement|movements
Event|Event|General Exam|3784,3791|true|false|false|||tremors
Finding|Sign or Symptom|General Exam|3784,3791|true|false|false|C0040822|Tremor|tremors
Event|Event|General Exam|3793,3801|false|false|false|||Strength
Finding|Idea or Concept|General Exam|3793,3801|false|false|false|C0808080|Strength (attribute)|Strength
Event|Event|General Exam|3827,3832|false|false|false|||power
Finding|Social Behavior|General Exam|3827,3832|false|false|false|C0032863|Power (Psychology)|power
Finding|Pathologic Function|General Exam|3853,3867|true|false|false|C1504476|Pronator drift|pronator drift
Event|Event|General Exam|3862,3867|true|false|false|||drift
Event|Event|General Exam|3869,3878|true|false|false|||Sensation
Finding|Finding|General Exam|3869,3878|true|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Finding|Organ or Tissue Function|General Exam|3869,3878|true|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Procedure|Health Care Activity|General Exam|3869,3878|true|false|false|C2229507|sensory exam|Sensation
Event|Event|General Exam|3880,3886|false|false|false|||Intact
Finding|Finding|General Exam|3880,3886|false|false|false|C1554187|Gender Status - Intact|Intact
Drug|Amino Acid, Peptide, or Protein|General Exam|3890,3895|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|General Exam|3890,3895|false|false|false|C1570446|TNFSF14 protein, human|light
Event|Event|General Exam|3890,3895|false|false|false|||light
Finding|Finding|General Exam|3890,3895|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|General Exam|3890,3895|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|General Exam|3890,3895|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|General Exam|3890,3895|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|General Exam|3890,3895|false|false|false|C0031765|Phototherapy|light
Finding|Physiologic Function|General Exam|3890,3901|false|false|false|C0423553|Light touch|light touch
Event|Event|General Exam|3896,3901|false|false|false|||touch
Finding|Mental Process|General Exam|3896,3901|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Finding|Organ or Tissue Function|General Exam|3896,3901|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Procedure|Therapeutic or Preventive Procedure|General Exam|3896,3901|false|false|false|C0152054|Therapeutic Touch|touch
Event|Event|General Exam|3928,3931|false|false|false|||MRI
Finding|Gene or Genome|General Exam|3928,3931|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|General Exam|3928,3931|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|General Exam|3928,3931|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Diagnostic Procedure|General Exam|3928,3936|false|false|false|C0412674|MRI of head|MRI HEAD
Anatomy|Body Location or Region|General Exam|3932,3936|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|HEAD
Anatomy|Body Part, Organ, or Organ Component|General Exam|3932,3936|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|HEAD
Disorder|Disease or Syndrome|General Exam|3932,3936|false|false|false|C0362076|Problems with head|HEAD
Event|Event|General Exam|3932,3936|false|false|false|||HEAD
Procedure|Therapeutic or Preventive Procedure|General Exam|3932,3936|false|false|false|C0876917|Procedure on head|HEAD
Event|Event|General Exam|3938,3939|false|false|false|||/
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|3942,3950|false|false|false|C0009924|Contrast Media|CONTRAST
Event|Event|General Exam|3942,3950|false|false|false|||CONTRAST
Drug|Biomedical or Dental Material|Impression|3972,3976|false|false|false|C1882953|Ring Dosage Form|Ring
Event|Event|Impression|3987,3993|false|false|false|||lesion
Finding|Finding|Impression|3987,3993|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|Impression|3987,3993|false|false|false|C0221198;C1546698|Lesion|lesion
Event|Event|Impression|3994,4004|false|false|false|||identified
Event|Governmental or Regulatory Activity|Impression|4012,4016|false|false|false|C1510751|Academic Research Enhancement Awards|area
Finding|Functional Concept|Impression|4024,4029|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Space or Junction|Impression|4043,4049|false|false|false|C1184482;C3893558|Groove;dinoflagellate sulcus|sulcus
Anatomy|Cell Component|Impression|4043,4049|false|false|false|C1184482;C3893558|Groove;dinoflagellate sulcus|sulcus
Anatomy|Body Part, Organ, or Organ Component|Impression|4050,4062|false|false|false|C0016733|frontal lobe|frontal lobe
Disorder|Neoplastic Process|Impression|4050,4062|false|false|false|C0153635|malignant neoplasm of frontal lobe|frontal lobe
Anatomy|Body Part, Organ, or Organ Component|Impression|4058,4062|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|Impression|4058,4062|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Finding|Finding|Impression|4080,4095|false|false|false|C2825502|Vasogenic Edema|vasogenic edema
Attribute|Clinical Attribute|Impression|4090,4095|false|false|false|C1717255||edema
Event|Event|Impression|4090,4095|false|false|false|||edema
Finding|Pathologic Function|Impression|4090,4095|false|false|false|C0013604|Edema|edema
Event|Event|Impression|4097,4107|false|false|false|||restricted
Finding|Functional Concept|Impression|4097,4107|false|false|false|C0443288;C1548390;C1549594;C1610594|Confidentiality - restricted;Confidentiality code - Restricted;Document Confidentiality Status - Restricted;Restricted|restricted
Finding|Idea or Concept|Impression|4097,4107|false|false|false|C0443288;C1548390;C1549594;C1610594|Confidentiality - restricted;Confidentiality code - Restricted;Document Confidentiality Status - Restricted;Restricted|restricted
Finding|Intellectual Product|Impression|4097,4107|false|false|false|C0443288;C1548390;C1549594;C1610594|Confidentiality - restricted;Confidentiality code - Restricted;Document Confidentiality Status - Restricted;Restricted|restricted
Event|Event|Impression|4109,4118|false|false|false|||diffusion
Finding|Functional Concept|Impression|4109,4118|false|false|false|C1696141|Diffusion - RouteOfAdministration|diffusion
Phenomenon|Natural Phenomenon or Process|Impression|4109,4118|false|false|false|C0012222|Diffusion|diffusion
Finding|Finding|Impression|4120,4128|false|false|false|C0332149|Possible|possibly
Event|Event|Impression|4129,4139|false|false|false|||consistent
Finding|Idea or Concept|Impression|4129,4139|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|Impression|4129,4144|false|false|false|C0332290|Consistent with|consistent with
Disorder|Disease or Syndrome|Impression|4148,4155|true|false|false|C0000833|Abscess|abscess
Event|Event|Impression|4148,4155|true|false|false|||abscess
Finding|Intellectual Product|Impression|4148,4155|true|false|false|C1546533||abscess
Event|Event|Impression|4163,4171|true|false|false|||entities
Finding|Intellectual Product|Impression|4183,4193|true|true|false|C4554154|Completely - dosing instruction fragment|completely
Event|Event|Impression|4194,4199|true|false|false|||ruled
Disorder|Neoplastic Process|Impression|4212,4222|true|true|false|C0027627;C2939419|Metastatic malignant neoplasm;Neoplasm Metastasis|metastases
Event|Event|Impression|4212,4222|true|false|false|||metastases
Finding|Finding|Impression|4212,4222|true|true|false|C1513183|Metastatic Lesion|metastases
Anatomy|Body Part, Organ, or Organ Component|Impression|4235,4240|false|false|false|C0006104;C4266577|Brain;Head>Brain|brain
Disorder|Disease or Syndrome|Impression|4235,4240|false|false|false|C0006111|Brain Diseases|brain
Disorder|Neoplastic Process|Impression|4235,4249|false|false|false|C0006118|Brain Neoplasms|brain neoplasm
Disorder|Neoplastic Process|Impression|4241,4249|false|false|false|C0027651;C1882062|Neoplasms;Neoplastic disease|neoplasm
Event|Event|Impression|4241,4249|false|false|false|||neoplasm
Drug|Organic Chemical|Impression|4268,4273|false|false|false|C0309093|FLAIR (product)|FLAIR
Drug|Pharmacologic Substance|Impression|4268,4273|false|false|false|C0309093|FLAIR (product)|FLAIR
Event|Event|Impression|4268,4273|false|false|false|||FLAIR
Procedure|Diagnostic Procedure|Impression|4268,4273|false|false|false|C2826145|Fluid Attenuated Inversion Recovery|FLAIR
Event|Event|Impression|4294,4301|false|false|false|||lesions
Finding|Finding|Impression|4294,4301|false|false|false|C0221198|Lesion|lesions
Anatomy|Body Location or Region|Impression|4310,4321|false|false|false|C0815275|Subcortical|subcortical
Anatomy|Tissue|Impression|4322,4334|false|false|false|C0682708|White matter|white matter
Drug|Amino Acid Sequence|Impression|4359,4365|false|false|false|C1514562|Protein Domain|region
Event|Event|Impression|4368,4378|false|false|false|||consistent
Finding|Idea or Concept|Impression|4368,4378|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|Impression|4368,4383|false|false|false|C0332290|Consistent with|consistent with
Disorder|Disease or Syndrome|Impression|4390,4408|false|false|false|C0026769|Multiple Sclerosis|multiple sclerosis
Finding|Pathologic Function|Impression|4399,4408|false|false|false|C0036429|Sclerosis|sclerosis
Disorder|Disease or Syndrome|Impression|4409,4416|false|true|false|C0012634|Disease|disease
Event|Event|Impression|4409,4416|false|false|false|||disease
Event|Event|Impression|4424,4427|false|false|false|||MRI
Finding|Gene or Genome|Impression|4424,4427|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|Impression|4424,4427|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|Impression|4424,4427|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Diagnostic Procedure|Impression|4424,4432|false|false|false|C0412674|MRI of head|MRI HEAD
Anatomy|Body Location or Region|Impression|4428,4432|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|HEAD
Anatomy|Body Part, Organ, or Organ Component|Impression|4428,4432|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|HEAD
Disorder|Disease or Syndrome|Impression|4428,4432|false|false|false|C0362076|Problems with head|HEAD
Event|Event|Impression|4428,4432|false|false|false|||HEAD
Procedure|Therapeutic or Preventive Procedure|Impression|4428,4432|false|false|false|C0876917|Procedure on head|HEAD
Drug|Indicator, Reagent, or Diagnostic Aid|Impression|4436,4444|false|false|false|C0009924|Contrast Media|CONTRAST
Event|Event|Impression|4436,4444|false|false|false|||CONTRAST
Event|Event|Impression|4446,4456|false|false|false|||IMPRESSION
Finding|Intellectual Product|Impression|4446,4456|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|Impression|4446,4456|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Finding|Impression|4459,4468|false|false|false|C0442739||Unchanged
Drug|Biomedical or Dental Material|Impression|4469,4473|false|false|false|C1882953|Ring Dosage Form|ring
Event|Event|Impression|4474,4483|false|false|false|||enhancing
Event|Event|Impression|4484,4490|false|false|false|||lesion
Finding|Finding|Impression|4484,4490|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|Impression|4484,4490|false|false|false|C0221198;C1546698|Lesion|lesion
Event|Event|Impression|4491,4501|false|false|false|||identified
Event|Governmental or Regulatory Activity|Impression|4510,4514|false|false|false|C1510751|Academic Research Enhancement Awards|area
Finding|Functional Concept|Impression|4523,4528|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Space or Junction|Impression|4523,4546|false|false|false|C2953689|Right precentral sulcus|right precentral sulcus
Anatomy|Body Space or Junction|Impression|4529,4546|false|false|false|C0228201|Structure of precentral sulcus|precentral sulcus
Anatomy|Body Space or Junction|Impression|4540,4546|false|false|false|C1184482;C3893558|Groove;dinoflagellate sulcus|sulcus
Anatomy|Cell Component|Impression|4540,4546|false|false|false|C1184482;C3893558|Groove;dinoflagellate sulcus|sulcus
Anatomy|Body Part, Organ, or Organ Component|Impression|4554,4566|false|false|false|C0016733|frontal lobe|frontal lobe
Disorder|Neoplastic Process|Impression|4554,4566|false|false|false|C0153635|malignant neoplasm of frontal lobe|frontal lobe
Anatomy|Body Part, Organ, or Organ Component|Impression|4562,4566|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|Impression|4562,4566|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Finding|Finding|Impression|4585,4600|false|false|false|C2825502|Vasogenic Edema|vasogenic edema
Attribute|Clinical Attribute|Impression|4595,4600|false|false|false|C1717255||edema
Event|Event|Impression|4595,4600|false|false|false|||edema
Finding|Pathologic Function|Impression|4595,4600|false|false|false|C0013604|Edema|edema
Finding|Idea or Concept|Impression|4607,4619|false|false|false|C1549478|Amount type - Differential|differential
Attribute|Clinical Attribute|Impression|4607,4629|false|false|false|C4760371||differential diagnosis
Procedure|Diagnostic Procedure|Impression|4607,4629|false|false|false|C0011906|Differential Diagnosis|differential diagnosis
Attribute|Clinical Attribute|Impression|4620,4629|false|false|false|C0945731||diagnosis
Event|Event|Impression|4620,4629|false|false|false|||diagnosis
Finding|Classification|Impression|4620,4629|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|Impression|4620,4629|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|Impression|4620,4629|false|false|false|C0011900|Diagnosis|diagnosis
Finding|Functional Concept|Impression|4636,4644|false|false|false|C0332257|Including (qualifier)|includes
Finding|Finding|Impression|4646,4654|false|false|false|C0332149|Possible|possible
Disorder|Disease or Syndrome|Impression|4655,4662|false|false|false|C0000833|Abscess|abscess
Event|Event|Impression|4655,4662|false|false|false|||abscess
Finding|Intellectual Product|Impression|4655,4662|false|false|false|C1546533||abscess
Event|Event|Impression|4670,4678|false|false|false|||entities
Finding|Intellectual Product|Impression|4699,4709|true|true|false|C4554154|Completely - dosing instruction fragment|completely
Event|Event|Impression|4711,4719|true|false|false|||excluded
Drug|Indicator, Reagent, or Diagnostic Aid|Impression|4731,4739|false|false|false|C0009924|Contrast Media|CONTRAST
Procedure|Diagnostic Procedure|Impression|4731,4747|false|false|false|C1275583|Computerized axial tomography of brain with radiopaque contrast|CONTRAST HEAD CT
Anatomy|Body Location or Region|Impression|4740,4744|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|HEAD
Anatomy|Body Part, Organ, or Organ Component|Impression|4740,4744|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|HEAD
Disorder|Disease or Syndrome|Impression|4740,4744|false|false|false|C0362076|Problems with head|HEAD
Procedure|Therapeutic or Preventive Procedure|Impression|4740,4744|false|false|false|C0876917|Procedure on head|HEAD
Procedure|Diagnostic Procedure|Impression|4740,4747|false|false|false|C0202691|CAT scan of head|HEAD CT
Event|Event|Impression|4745,4747|false|false|false|||CT
Attribute|Clinical Attribute|Impression|4769,4775|false|false|false|C5889824||Status
Event|Event|Impression|4769,4775|false|false|false|||Status
Finding|Idea or Concept|Impression|4769,4775|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|Impression|4781,4786|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Event|Event|Impression|4796,4806|false|false|false|||craniotomy
Procedure|Therapeutic or Preventive Procedure|Impression|4796,4806|false|false|false|C0010280|Craniotomy|craniotomy
Event|Event|Impression|4818,4825|false|false|false|||density
Event|Event|Impression|4827,4833|false|false|false|||lesion
Finding|Finding|Impression|4827,4833|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|Impression|4827,4833|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Functional Concept|Impression|4842,4847|true|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Space or Junction|Impression|4842,4865|true|false|false|C2953689|Right precentral sulcus|right precentral sulcus
Anatomy|Body Space or Junction|Impression|4848,4865|true|false|false|C0228201|Structure of precentral sulcus|precentral sulcus
Anatomy|Body Space or Junction|Impression|4859,4865|true|false|false|C1184482;C3893558|Groove;dinoflagellate sulcus|sulcus
Anatomy|Cell Component|Impression|4859,4865|true|false|false|C1184482;C3893558|Groove;dinoflagellate sulcus|sulcus
Attribute|Clinical Attribute|Impression|4882,4887|true|false|false|C1717255||edema
Event|Event|Impression|4882,4887|true|false|false|||edema
Finding|Pathologic Function|Impression|4882,4887|true|false|false|C0013604|Edema|edema
Event|Event|Impression|4907,4914|true|false|false|||changed
Event|Event|Impression|4936,4944|false|false|false|||allowing
Event|Event|Impression|4950,4960|false|false|false|||difference
Event|Event|Impression|4964,4973|false|false|false|||technique
Finding|Functional Concept|Impression|4964,4973|false|false|false|C0449851|Techniques|technique
Finding|Intellectual Product|Impression|4987,4992|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Location or Region|Impression|4993,5005|true|false|false|C0524466|Intracranial|intracranial
Finding|Functional Concept|Impression|4993,5005|true|false|false|C1522213|Intracranial Route of Administration|intracranial
Finding|Pathologic Function|Impression|4993,5016|true|false|false|C0151699|Intracranial Hemorrhage|intracranial hemorrhage
Event|Event|Impression|5006,5016|true|false|false|||hemorrhage
Finding|Pathologic Function|Impression|5006,5016|true|false|false|C0019080|Hemorrhage|hemorrhage
Finding|Classification|Impression|5020,5025|true|true|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|major
Anatomy|Body Part, Organ, or Organ Component|Impression|5026,5034|true|false|false|C0005847|Blood Vessel|vascular
Event|Event|Impression|5048,5055|false|false|false|||infarct
Finding|Pathologic Function|Impression|5048,5055|false|false|false|C0021308|Infarction|infarct
Anatomy|Body Location or Region|Impression|5076,5087|false|false|false|C0815275|Subcortical|subcortical
Anatomy|Tissue|Impression|5088,5100|false|false|false|C0682708|White matter|white matter
Event|Event|Impression|5115,5125|false|false|false|||compatible
Finding|Idea or Concept|Impression|5115,5125|false|false|false|C0332290|Consistent with|compatible
Disorder|Disease or Syndrome|Impression|5144,5162|false|false|false|C0026769|Multiple Sclerosis|multiple sclerosis
Event|Event|Impression|5153,5162|false|false|false|||sclerosis
Finding|Pathologic Function|Impression|5153,5162|false|false|false|C0036429|Sclerosis|sclerosis
Disorder|Congenital Abnormality|Impression|5179,5182|false|false|false|C5889736|Isolated femoral agenesis/hypoplasia|CSF
Drug|Amino Acid, Peptide, or Protein|Impression|5179,5182|false|false|false|C0009392;C0376561;C5197246|CSF2 protein, human;Colony-Stimulating Factors;Recombinant Colony-Stimulating Factors|CSF
Drug|Biologically Active Substance|Impression|5179,5182|false|false|false|C0009392;C0376561;C5197246|CSF2 protein, human;Colony-Stimulating Factors;Recombinant Colony-Stimulating Factors|CSF
Drug|Immunologic Factor|Impression|5179,5182|false|false|false|C0009392;C0376561;C5197246|CSF2 protein, human;Colony-Stimulating Factors;Recombinant Colony-Stimulating Factors|CSF
Drug|Pharmacologic Substance|Impression|5179,5182|false|false|false|C0009392;C0376561;C5197246|CSF2 protein, human;Colony-Stimulating Factors;Recombinant Colony-Stimulating Factors|CSF
Event|Event|Impression|5179,5182|false|false|false|||CSF
Finding|Body Substance|Impression|5179,5182|false|false|false|C0007806;C0007807;C3889436|Cerebrospinal Fluid;In Cerebrospinal Fluid;LAMC2 wt Allele|CSF
Finding|Functional Concept|Impression|5179,5182|false|false|false|C0007806;C0007807;C3889436|Cerebrospinal Fluid;In Cerebrospinal Fluid;LAMC2 wt Allele|CSF
Finding|Gene or Genome|Impression|5179,5182|false|false|false|C0007806;C0007807;C3889436|Cerebrospinal Fluid;In Cerebrospinal Fluid;LAMC2 wt Allele|CSF
Procedure|Therapeutic or Preventive Procedure|Impression|5179,5182|false|false|false|C3540512|Circumferential Supracrestal Fiberotomy|CSF
Finding|Body Substance|Impression|5183,5195|false|false|false|C0007806|Cerebrospinal Fluid|SPINAL FLUID
Drug|Substance|Impression|5190,5195|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|FLUID
Event|Event|Impression|5190,5195|false|false|false|||FLUID
Finding|Intellectual Product|Impression|5190,5195|false|false|false|C1546638|Fluid Specimen Code|FLUID
Event|Event|Impression|5201,5205|false|false|false|||TUBE
Finding|Functional Concept|Impression|5201,5205|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|TUBE
Finding|Gene or Genome|Impression|5201,5205|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|TUBE
Drug|Indicator, Reagent, or Diagnostic Aid|Impression|5215,5225|false|false|false|C0061856|Gram's stain|GRAM STAIN
Drug|Organic Chemical|Impression|5215,5225|false|false|false|C0061856|Gram's stain|GRAM STAIN
Procedure|Laboratory Procedure|Impression|5215,5225|false|false|false|C0200966|Bacterial stain, routine|GRAM STAIN
Drug|Indicator, Reagent, or Diagnostic Aid|Impression|5220,5225|false|false|false|C0038128|Stains|STAIN
Event|Event|Impression|5220,5225|false|false|false|||STAIN
Procedure|Laboratory Procedure|Impression|5220,5225|false|false|false|C0487602|Staining method|STAIN
Finding|Idea or Concept|Impression|5227,5232|false|false|false|C1546485|Diagnosis Type - Final|Final
Anatomy|Cell|Impression|5248,5276|true|false|false|C0018183;C0027950|granulocyte;neutrophil|POLYMORPHONUCLEAR LEUKOCYTES
Anatomy|Cell|Impression|5266,5276|true|false|false|C0023516|Leukocytes|LEUKOCYTES
Finding|Body Substance|Impression|5266,5276|true|false|false|C1547962;C1550647|Specimen Type - Leukocytes|LEUKOCYTES
Finding|Intellectual Product|Impression|5266,5276|true|false|false|C1547962;C1550647|Specimen Type - Leukocytes|LEUKOCYTES
Event|Event|Impression|5277,5281|true|false|false|||SEEN
Finding|Finding|Impression|5293,5312|true|false|false|C2924473|Microorganisms seen|MICROORGANISMS SEEN
Event|Event|Impression|5308,5312|true|false|false|||SEEN
Event|Activity|Impression|5344,5349|false|false|false|C1947932|Smear - instruction imperative|smear
Event|Event|Impression|5344,5349|false|false|false|||smear
Finding|Functional Concept|Impression|5344,5349|false|false|false|C3872789|Smearing technique|smear
Procedure|Diagnostic Procedure|Impression|5344,5349|false|false|false|C0444186|Smear test|smear
Event|Event|Impression|5367,5373|false|false|false|||method
Finding|Functional Concept|Impression|5367,5373|false|false|false|C0025663;C0449851;C2828387|Method, LOINC Axis 6;Methods;Techniques|method
Finding|Intellectual Product|Impression|5367,5373|false|false|false|C0025663;C0449851;C2828387|Method, LOINC Axis 6;Methods;Techniques|method
Event|Event|Impression|5398,5408|false|false|false|||hematology
Finding|Intellectual Product|Impression|5398,5408|false|false|false|C1547985|Diagnostic Service Section ID - Hematology|hematology
Procedure|Laboratory Procedure|Impression|5398,5408|false|false|false|C0018941;C0200627;C2183233|Hematologic Tests;Hematology procedure;diagnostic service sources hematology (procedure)|hematology
Anatomy|Cell|Impression|5428,5444|false|false|false|C0023516|Leukocytes|white blood cell
Lab|Laboratory or Test Result|Impression|5428,5450|false|false|false|C0427512||white blood cell count
Procedure|Laboratory Procedure|Impression|5428,5450|false|false|false|C0023508|White Blood Cell Count procedure|white blood cell count
Disorder|Disease or Syndrome|Impression|5434,5439|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|Impression|5434,5439|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Anatomy|Cell|Impression|5434,5444|false|false|false|C0005773|Blood Cells|blood cell
Procedure|Laboratory Procedure|Impression|5434,5450|false|false|false|C0005771;C0009555|Blood Cell Count;Complete Blood Count|blood cell count
Anatomy|Cell|Impression|5440,5444|false|false|false|C0007634|Cells|cell
Finding|Gene or Genome|Impression|5440,5444|false|false|false|C1413336;C1413337|CEL gene;CELP gene|cell
Procedure|Laboratory Procedure|Impression|5440,5450|false|false|false|C0007584|Cell Count|cell count
Event|Event|Impression|5445,5450|false|false|false|||count
Drug|Substance|Impression|5458,5463|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|FLUID
Finding|Intellectual Product|Impression|5458,5463|false|false|false|C1546638|Fluid Specimen Code|FLUID
Drug|Biomedical or Dental Material|Impression|5464,5471|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|Impression|5464,5471|false|false|false|||CULTURE
Finding|Functional Concept|Impression|5464,5471|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|Impression|5464,5471|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|Impression|5464,5471|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|Impression|5493,5499|true|false|false|||GROWTH
Finding|Finding|Impression|5493,5499|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organ or Tissue Function|Impression|5493,5499|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organism Function|Impression|5493,5499|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Physiologic Function|Impression|5493,5499|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Phenomenon|Phenomenon or Process|Impression|5493,5499|true|false|false|C2911660|Growth action|GROWTH
Event|Event|Hospital Course|5536,5545|false|false|false|||presented
Finding|Finding|Hospital Course|5557,5566|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Idea or Concept|Hospital Course|5557,5566|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Intellectual Product|Hospital Course|5557,5566|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Pathologic Function|Hospital Course|5557,5566|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Phenomenon|Phenomenon or Process|Hospital Course|5557,5566|false|false|false|C0013956|Emergency Situation|Emergency
Procedure|Health Care Activity|Hospital Course|5557,5566|false|false|false|C1553500|emergency encounter|Emergency
Finding|Idea or Concept|Hospital Course|5567,5577|false|false|false|C1547537;C1548283;C1549615|Department - Charge type;Department - No suggested values defined;Organization Unit Type - Department|Department
Finding|Functional Concept|Hospital Course|5591,5595|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Event|Event|Hospital Course|5602,5610|false|false|false|||numbness
Finding|Finding|Hospital Course|5602,5610|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|Hospital Course|5602,5610|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5618,5622|false|false|false|C0018563;C4285005|Hand;Upper extremity>Hand|hand
Finding|Finding|Hospital Course|5618,5622|false|false|false|C0741992|Hand problem|hand
Anatomy|Body Location or Region|Hospital Course|5627,5631|false|false|false|C0015450;C4266571|Face;Head>Face|face
Disorder|Disease or Syndrome|Hospital Course|5627,5631|false|false|false|C3160739|FANCONI ANEMIA, COMPLEMENTATION GROUP E|face
Event|Event|Hospital Course|5627,5631|false|false|false|||face
Finding|Gene or Genome|Hospital Course|5627,5631|false|false|false|C1414531;C1423759;C2828055|ELOVL6 gene;FANCE gene;FANCE wt Allele|face
Event|Event|Hospital Course|5636,5640|false|false|false|||left
Finding|Functional Concept|Hospital Course|5636,5640|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5642,5646|false|false|false|C0018563;C4285005|Hand;Upper extremity>Hand|hand
Finding|Finding|Hospital Course|5642,5646|false|false|false|C0741992|Hand problem|hand
Event|Event|Hospital Course|5647,5657|false|false|false|||clumsiness
Finding|Sign or Symptom|Hospital Course|5647,5657|false|false|false|C0233844|Clumsiness|clumsiness
Event|Event|Hospital Course|5668,5677|false|false|false|||evaluated
Event|Event|Hospital Course|5703,5711|false|false|false|||believed
Event|Event|Hospital Course|5726,5731|false|false|false|||flare
Finding|Finding|Hospital Course|5726,5731|false|false|false|C1517205;C3540542|Exacerbation of cGVHD;Flare|flare
Finding|Sign or Symptom|Hospital Course|5726,5731|false|false|false|C1517205;C3540542|Exacerbation of cGVHD;Flare|flare
Event|Event|Hospital Course|5744,5752|false|false|false|||evaluted
Event|Occupational Activity|Hospital Course|5767,5774|false|false|false|C0557854|Services|service
Finding|Idea or Concept|Hospital Course|5767,5774|false|false|false|C3245478|ActInformationPrivacyReason - service|service
Event|Event|Hospital Course|5781,5789|false|false|false|||resulted
Event|Event|Hospital Course|5797,5811|false|false|false|||recommendation
Finding|Idea or Concept|Hospital Course|5797,5811|false|false|false|C0034866|Recommendation|recommendation
Event|Event|Hospital Course|5819,5822|false|false|false|||MRI
Finding|Gene or Genome|Hospital Course|5819,5822|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|Hospital Course|5819,5822|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|Hospital Course|5819,5822|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Diagnostic Procedure|Hospital Course|5819,5828|false|false|false|C4028269|Nuclear magnetic resonance imaging brain|MRI brain
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5823,5828|false|false|false|C0006104;C4266577|Brain;Head>Brain|brain
Disorder|Disease or Syndrome|Hospital Course|5823,5828|false|false|false|C0006111|Brain Diseases|brain
Event|Event|Hospital Course|5823,5828|false|false|false|||brain
Event|Event|Hospital Course|5836,5839|false|false|false|||MRI
Finding|Gene or Genome|Hospital Course|5836,5839|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|Hospital Course|5836,5839|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|Hospital Course|5836,5839|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Event|Event|Hospital Course|5844,5848|false|false|false|||read
Event|Event|Hospital Course|5852,5863|false|false|false|||demonstrate
Finding|Functional Concept|Hospital Course|5866,5871|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Event|Event|Hospital Course|5881,5887|false|false|false|||lesion
Finding|Finding|Hospital Course|5881,5887|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|Hospital Course|5881,5887|false|false|false|C0221198;C1546698|Lesion|lesion
Event|Event|Hospital Course|5889,5899|false|false|false|||concerning
Finding|Functional Concept|Hospital Course|5908,5918|false|false|false|C0036525;C1522484|Metastatic to;metastatic qualifier|metastatic
Disorder|Neoplastic Process|Hospital Course|5908,5926|false|false|false|C0027627;C2939419;C2939420|Metastatic Neoplasm;Metastatic malignant neoplasm;Neoplasm Metastasis|metastatic disease
Finding|Finding|Hospital Course|5908,5926|false|false|false|C1513183|Metastatic Lesion|metastatic disease
Disorder|Disease or Syndrome|Hospital Course|5919,5926|false|false|false|C0012634|Disease|disease
Event|Event|Hospital Course|5919,5926|false|false|false|||disease
Disorder|Disease or Syndrome|Hospital Course|5930,5937|false|true|false|C0000833|Abscess|abscess
Event|Event|Hospital Course|5930,5937|false|false|false|||abscess
Finding|Intellectual Product|Hospital Course|5930,5937|false|true|false|C1546533||abscess
Event|Event|Hospital Course|5948,5956|false|false|false|||admitted
Event|Event|Hospital Course|5960,5972|false|false|false|||Neurosurgery
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5960,5972|false|false|false|C0524850|Neurosurgical Procedures|Neurosurgery
Event|Event|Hospital Course|5985,5995|false|false|false|||evaluation
Finding|Idea or Concept|Hospital Course|5985,5995|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|Hospital Course|5985,5995|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Event|Event|Hospital Course|6000,6009|false|false|false|||treatment
Finding|Conceptual Entity|Hospital Course|6000,6009|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Hospital Course|6000,6009|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Hospital Course|6000,6009|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6000,6009|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Event|Event|Hospital Course|6035,6040|false|false|false|||taken
Finding|Functional Concept|Hospital Course|6057,6062|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Event|Event|Hospital Course|6073,6083|false|false|false|||craniotomy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6073,6083|false|false|false|C0010280|Craniotomy|craniotomy
Event|Event|Hospital Course|6103,6111|false|false|false|||drainage
Finding|Body Substance|Hospital Course|6103,6111|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|Hospital Course|6103,6111|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6103,6111|false|false|false|C0013103|Drainage procedure|drainage
Event|Event|Hospital Course|6116,6126|false|false|false|||irrigation
Finding|Functional Concept|Hospital Course|6116,6126|false|false|false|C1521919;C2314883|Irrigation Route of Administration;Irrigation [MoA]|irrigation
Finding|Molecular Function|Hospital Course|6116,6126|false|false|false|C1521919;C2314883|Irrigation Route of Administration;Irrigation [MoA]|irrigation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6116,6126|false|false|false|C0022100|Irrigation|irrigation
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6131,6136|false|false|false|C0006104;C4266577|Brain;Head>Brain|brain
Disorder|Disease or Syndrome|Hospital Course|6131,6136|false|false|false|C0006111|Brain Diseases|brain
Disorder|Disease or Syndrome|Hospital Course|6131,6144|false|false|false|C0006105;C1510428|Brain Abscess;Cerebral abscess|brain abscess
Disorder|Disease or Syndrome|Hospital Course|6137,6144|false|false|false|C0000833|Abscess|abscess
Event|Event|Hospital Course|6137,6144|false|false|false|||abscess
Finding|Intellectual Product|Hospital Course|6137,6144|false|false|false|C1546533||abscess
Event|Event|Hospital Course|6150,6159|false|false|false|||tolerated
Attribute|Clinical Attribute|Hospital Course|6164,6173|false|false|false|C0945766||procedure
Event|Event|Hospital Course|6164,6173|false|false|false|||procedure
Event|Occupational Activity|Hospital Course|6164,6173|false|false|false|C1546467|Act Class - procedure|procedure
Finding|Functional Concept|Hospital Course|6164,6173|false|false|false|C2700391|Procedure (set of actions)|procedure
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6164,6173|false|false|false|C0184661|Interventional procedure|procedure
Finding|Finding|Hospital Course|6174,6178|false|false|false|C5575035|Well (answer to question)|well
Event|Event|Hospital Course|6189,6194|false|false|false|||taken
Event|Event|Hospital Course|6198,6202|false|false|false|||PACU
Event|Event|Hospital Course|6206,6213|false|false|false|||recover
Finding|Intellectual Product|Hospital Course|6214,6218|false|false|false|C1720594|Then - dosing instruction fragment|then
Anatomy|Body Space or Junction|Hospital Course|6226,6229|false|false|false|C0228479|Structure of intraculminate fissure|ICU
Finding|Intellectual Product|Hospital Course|6226,6229|false|false|false|C4554035|Inventory of Callous-Unemotional Traits|ICU
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6246,6256|false|false|false|C0042313|vancomycin|Vancomycin
Drug|Antibiotic|Hospital Course|6246,6256|false|false|false|C0042313|vancomycin|Vancomycin
Event|Event|Hospital Course|6246,6256|false|false|false|||Vancomycin
Procedure|Laboratory Procedure|Hospital Course|6246,6256|false|false|false|C0489941|Vancomycin measurement|Vancomycin
Drug|Antibiotic|Hospital Course|6261,6270|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|Meropenem
Drug|Clinical Drug|Hospital Course|6261,6270|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|Meropenem
Drug|Organic Chemical|Hospital Course|6261,6270|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|Meropenem
Event|Event|Hospital Course|6261,6270|false|false|false|||Meropenem
Drug|Indicator, Reagent, or Diagnostic Aid|Hospital Course|6272,6282|false|false|false|C0061856|Gram's stain|Gram stain
Drug|Organic Chemical|Hospital Course|6272,6282|false|false|false|C0061856|Gram's stain|Gram stain
Procedure|Laboratory Procedure|Hospital Course|6272,6282|false|false|false|C0200966|Bacterial stain, routine|Gram stain
Drug|Indicator, Reagent, or Diagnostic Aid|Hospital Course|6277,6282|false|false|false|C0038128|Stains|stain
Event|Event|Hospital Course|6277,6282|false|false|false|||stain
Procedure|Laboratory Procedure|Hospital Course|6277,6282|false|false|false|C0487602|Staining method|stain
Finding|Classification|Hospital Course|6296,6304|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|6296,6304|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|6296,6304|false|false|false|C5237010|Expression Negative|negative
Anatomy|Cell|Hospital Course|6305,6309|false|false|false|C0206427|Rod Photoreceptors|rods
Disorder|Cell or Molecular Dysfunction|Hospital Course|6320,6328|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Event|Event|Hospital Course|6320,6328|false|false|false|||positive
Finding|Classification|Hospital Course|6320,6328|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|Hospital Course|6320,6328|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Event|Event|Hospital Course|6329,6334|false|false|false|||cocci
Event|Event|Hospital Course|6348,6354|false|false|false|||chains
Finding|Gene or Genome|Hospital Course|6356,6360|false|false|false|C3469826;C3470073|DESI1 gene;SLC35G1 gene|Post
Finding|Finding|Hospital Course|6356,6370|false|false|false|C0241311|post operative (finding)|Post operative
Anatomy|Body Location or Region|Hospital Course|6371,6375|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6371,6375|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|Hospital Course|6371,6375|false|false|false|C0362076|Problems with head|head
Event|Event|Hospital Course|6371,6375|false|false|false|||head
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6371,6375|false|false|false|C0876917|Procedure on head|head
Event|Event|Hospital Course|6380,6386|false|false|false|||showed
Finding|Gene or Genome|Hospital Course|6387,6391|false|false|false|C3469826;C3470073|DESI1 gene;SLC35G1 gene|post
Finding|Finding|Hospital Course|6387,6401|false|false|false|C0241311|post operative (finding)|post operative
Event|Event|Hospital Course|6402,6409|false|false|false|||changes
Finding|Functional Concept|Hospital Course|6402,6409|false|false|false|C0392747|Changing|changes
Finding|Finding|Hospital Course|6414,6428|false|false|false|C0241311|post operative (finding)|post operative
Event|Event|Hospital Course|6429,6433|false|false|false|||exam
Finding|Functional Concept|Hospital Course|6429,6433|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|Hospital Course|6429,6433|false|false|false|C0582103|Medical Examination|exam
Finding|Functional Concept|Hospital Course|6443,6447|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6443,6451|false|false|false|C0230347;C5779993|Left arm;Left upper arm structure|left arm
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6448,6451|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|Hospital Course|6448,6451|false|false|false|C3495676|Anorectal Malformations|arm
Event|Event|Hospital Course|6448,6451|false|false|false|||arm
Finding|Gene or Genome|Hospital Course|6448,6451|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|Hospital Course|6448,6451|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|Hospital Course|6448,6451|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6448,6451|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Finding|Sign or Symptom|Hospital Course|6448,6460|false|false|false|C0751409|Upper Extremity Paresis|arm weakness
Event|Event|Hospital Course|6452,6460|false|false|false|||weakness
Finding|Sign or Symptom|Hospital Course|6452,6460|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Finding|Body Substance|Hospital Course|6475,6482|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|6475,6482|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|6475,6482|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|6483,6492|false|false|false|||continued
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6496,6506|false|false|false|C0042313|vancomycin|vancomycin
Drug|Antibiotic|Hospital Course|6496,6506|false|false|false|C0042313|vancomycin|vancomycin
Event|Event|Hospital Course|6496,6506|false|false|false|||vancomycin
Procedure|Laboratory Procedure|Hospital Course|6496,6506|false|false|false|C0489941|Vancomycin measurement|vancomycin
Drug|Antibiotic|Hospital Course|6511,6520|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|Meropenem
Drug|Clinical Drug|Hospital Course|6511,6520|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|Meropenem
Drug|Organic Chemical|Hospital Course|6511,6520|false|false|false|C0066005;C1314417|INJECTION, MEROPENEM, 100 MG ADMINISTERED;meropenem|Meropenem
Event|Event|Hospital Course|6511,6520|false|false|false|||Meropenem
Anatomy|Cell|Hospital Course|6523,6526|false|false|false|C0023516|Leukocytes|WBC
Event|Event|Hospital Course|6531,6539|false|false|false|||elevated
Event|Event|Hospital Course|6575,6586|false|false|false|||transferred
Anatomy|Anatomical Structure|Hospital Course|6594,6599|false|false|false|C3714591|Floor (anatomic)|floor
Finding|Functional Concept|Hospital Course|6601,6605|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6601,6609|false|false|false|C0230347;C5779993|Left arm;Left upper arm structure|Left arm
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6606,6609|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|Hospital Course|6606,6609|false|false|false|C3495676|Anorectal Malformations|arm
Event|Event|Hospital Course|6606,6609|false|false|false|||arm
Finding|Gene or Genome|Hospital Course|6606,6609|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|Hospital Course|6606,6609|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|Hospital Course|6606,6609|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6606,6609|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Finding|Sign or Symptom|Hospital Course|6606,6618|false|false|false|C0751409|Upper Extremity Paresis|arm weakness
Event|Event|Hospital Course|6610,6618|false|false|false|||weakness
Finding|Sign or Symptom|Hospital Course|6610,6618|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Finding|Body Substance|Hospital Course|6647,6654|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|6647,6654|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|6647,6654|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|6655,6663|false|false|false|||reported
Event|Event|Hospital Course|6664,6672|false|false|false|||lethargy
Finding|Sign or Symptom|Hospital Course|6664,6672|false|false|false|C0023380|Lethargy|lethargy
Finding|Functional Concept|Hospital Course|6677,6681|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6677,6685|false|false|false|C0230416;C0230443|Left lower extremity;Structure of left lower leg|left leg
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6682,6685|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Finding|Hospital Course|6682,6694|false|false|false|C0427068;C1836296|Monoparesis of lower limb;Muscle Weakness Lower Limb|leg weakness
Event|Event|Hospital Course|6686,6694|false|false|false|||weakness
Finding|Sign or Symptom|Hospital Course|6686,6694|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Event|Event|Hospital Course|6700,6704|false|false|false|||exam
Finding|Functional Concept|Hospital Course|6700,6704|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|Hospital Course|6700,6704|false|false|false|C0582103|Medical Examination|exam
Finding|Body Substance|Hospital Course|6709,6716|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|6709,6716|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|6709,6716|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|6721,6727|false|false|false|||sleepy
Finding|Finding|Hospital Course|6721,6727|false|false|false|C0013144|Drowsiness|sleepy
Event|Event|Hospital Course|6732,6737|false|false|false|||awake
Finding|Finding|Hospital Course|6732,6737|false|false|false|C0234422|Awake (finding)|awake
Event|Event|Hospital Course|6748,6756|false|false|false|||oriented
Attribute|Clinical Attribute|Hospital Course|6761,6767|false|false|false|C5890614||person
Finding|Intellectual Product|Hospital Course|6761,6767|false|false|false|C1522390|Person Info|person
Event|Activity|Hospital Course|6768,6773|false|false|false|C1882509|put - instruction imperative|place
Event|Event|Hospital Course|6768,6773|false|false|false|||place
Finding|Functional Concept|Hospital Course|6768,6773|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|Hospital Course|6768,6773|false|false|false|C1533810||place
Finding|Finding|Hospital Course|6778,6782|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Hospital Course|6778,6782|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Hospital Course|6778,6782|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Functional Concept|Hospital Course|6785,6790|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Event|Event|Hospital Course|6797,6805|false|false|false|||strength
Finding|Idea or Concept|Hospital Course|6797,6805|false|false|false|C0808080|Strength (attribute)|strength
Finding|Functional Concept|Hospital Course|6818,6822|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6824,6839|false|false|false|C1140618|Upper Extremity|upper extremity
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6830,6839|false|false|false|C0015385|Limb structure|extremity
Finding|Functional Concept|Hospital Course|6852,6856|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6852,6872|false|false|false|C0230416|Left lower extremity|left lower extremity
Anatomy|Body Location or Region|Hospital Course|6857,6862|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|Hospital Course|6857,6862|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6857,6872|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6863,6872|false|false|false|C0015385|Limb structure|extremity
Event|Event|Hospital Course|6882,6888|false|false|false|||except
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6913,6917|false|false|false|C1366753|STAT protein|stat
Drug|Biologically Active Substance|Hospital Course|6913,6917|false|false|false|C1366753|STAT protein|stat
Finding|Gene or Genome|Hospital Course|6913,6917|false|false|false|C1335960;C1420304;C1547583;C1548425;C1561443|Extended Priority Codes - Stat;Referral priority - STAT;Report priority - Stat;SOAT1 gene;STAT family gene|stat
Finding|Idea or Concept|Hospital Course|6913,6917|false|false|false|C1335960;C1420304;C1547583;C1548425;C1561443|Extended Priority Codes - Stat;Referral priority - STAT;Report priority - Stat;SOAT1 gene;STAT family gene|stat
Finding|Intellectual Product|Hospital Course|6913,6917|false|false|false|C1335960;C1420304;C1547583;C1548425;C1561443|Extended Priority Codes - Stat;Referral priority - STAT;Report priority - Stat;SOAT1 gene;STAT family gene|stat
Event|Event|Hospital Course|6918,6923|false|false|false|||NCHCT
Event|Event|Hospital Course|6949,6955|false|false|false|||stable
Finding|Intellectual Product|Hospital Course|6949,6955|false|false|false|C1547311|Patient Condition Code - Stable|stable
Attribute|Clinical Attribute|Hospital Course|6966,6973|false|false|false|C2923685||consent
Event|Event|Hospital Course|6966,6973|false|false|false|||consent
Finding|Idea or Concept|Hospital Course|6966,6973|false|false|false|C1511481;C1554192;C5702721|ActClass - consent;Consent;Consent (record artifact)|consent
Finding|Intellectual Product|Hospital Course|6966,6973|false|false|false|C1511481;C1554192;C5702721|ActClass - consent;Consent;Consent (record artifact)|consent
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6978,6982|false|false|false|C2049629|Peripherally Inserted Central Catheter Line Insertion|picc
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6978,6997|false|false|false|C2049629|Peripherally Inserted Central Catheter Line Insertion|picc line placement
Drug|Biologically Active Substance|Hospital Course|6983,6987|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Hospital Course|6983,6987|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Substance|Hospital Course|6983,6987|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Event|Event|Hospital Course|6983,6987|false|false|false|||line
Finding|Intellectual Product|Hospital Course|6983,6987|false|false|false|C1546701|line source specimen code|line
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6983,6997|false|false|false|C1519955|Vascular Access Device Placement|line placement
Event|Event|Hospital Course|6988,6997|false|false|false|||placement
Procedure|Health Care Activity|Hospital Course|6988,6997|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6988,6997|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Event|Event|Hospital Course|6998,7006|false|false|false|||obtained
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7008,7012|false|false|false|C2049629|Peripherally Inserted Central Catheter Line Insertion|picc
Drug|Biologically Active Substance|Hospital Course|7013,7017|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Hospital Course|7013,7017|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Substance|Hospital Course|7013,7017|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Event|Event|Hospital Course|7013,7017|false|false|false|||line
Finding|Intellectual Product|Hospital Course|7013,7017|false|false|false|C1546701|line source specimen code|line
Event|Event|Hospital Course|7019,7025|false|false|false|||placed
Event|Event|Hospital Course|7048,7056|false|false|false|||continue
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7062,7067|false|false|false|C0042313|vancomycin|vanco
Drug|Antibiotic|Hospital Course|7062,7067|false|false|false|C0042313|vancomycin|vanco
Event|Event|Hospital Course|7062,7067|false|false|false|||vanco
Event|Event|Hospital Course|7072,7081|false|false|false|||meropenum
Finding|Idea or Concept|Hospital Course|7087,7092|false|false|false|C1546485|Diagnosis Type - Final|Final
Event|Event|Hospital Course|7093,7099|false|false|false|||abcess
Finding|Body Substance|Hospital Course|7093,7099|false|false|false|C1550609|Specimen Type - Abscess|abcess
Drug|Biomedical or Dental Material|Hospital Course|7100,7107|false|false|false|C1706355|Culture Dose Form|culture
Event|Event|Hospital Course|7100,7107|false|false|false|||culture
Finding|Functional Concept|Hospital Course|7100,7107|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Finding|Idea or Concept|Hospital Course|7100,7107|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Procedure|Laboratory Procedure|Hospital Course|7100,7107|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|culture
Lab|Laboratory or Test Result|Hospital Course|7100,7114|false|false|false|C2061903|culture result|culture result
Event|Event|Hospital Course|7108,7114|false|false|false|||result
Finding|Finding|Hospital Course|7108,7114|false|false|false|C1274040;C1546471;C2825142|Experimental Result;Result;What subject filter - Result|result
Finding|Functional Concept|Hospital Course|7108,7114|false|false|false|C1274040;C1546471;C2825142|Experimental Result;Result;What subject filter - Result|result
Finding|Idea or Concept|Hospital Course|7108,7114|false|false|false|C1274040;C1546471;C2825142|Experimental Result;Result;What subject filter - Result|result
Disorder|Disease or Syndrome|Hospital Course|7118,7123|false|false|false|C1410088|Still|still
Event|Event|Hospital Course|7124,7131|false|false|false|||pending
Finding|Idea or Concept|Hospital Course|7124,7131|false|false|false|C1691786;C1704475|Pending - Allergy Clinical Status;Pending - referral status|pending
Finding|Functional Concept|Hospital Course|7133,7137|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|Hospital Course|7133,7137|false|false|false|C0582103|Medical Examination|Exam
Event|Event|Hospital Course|7147,7153|false|false|false|||stable
Finding|Intellectual Product|Hospital Course|7147,7153|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|Hospital Course|7168,7177|false|false|false|||evaluated
Finding|Body Substance|Hospital Course|7182,7189|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|7182,7189|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|7182,7189|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|7194,7199|false|false|false|||found
Event|Event|Hospital Course|7209,7218|false|false|false|||continues
Finding|Finding|Hospital Course|7231,7244|true|false|false|C0231686|Gait, Unsteady|unsteady gait
Event|Event|Hospital Course|7240,7244|true|false|false|||gait
Finding|Finding|Hospital Course|7240,7244|true|false|false|C0016928|Gait|gait
Event|Event|Hospital Course|7262,7266|true|false|false|||safe
Finding|Intellectual Product|Hospital Course|7262,7266|true|true|true|C4684764|SAFE-Biopharma Standard|safe
Event|Event|Hospital Course|7273,7277|true|false|false|||home
Finding|Idea or Concept|Hospital Course|7273,7277|true|false|true|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|7273,7277|true|false|true|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|7273,7277|true|false|true|C1553498|home health encounter|home
Event|Event|Hospital Course|7286,7293|false|false|false|||planned
Event|Event|Hospital Course|7297,7302|false|false|false|||visit
Event|Event|Hospital Course|7324,7337|false|false|false|||re-evaluation
Procedure|Research Activity|Hospital Course|7324,7337|false|false|false|C0681840|re-evaluation|re-evaluation
Event|Event|Hospital Course|7360,7369|false|false|false|||maneuvers
Finding|Idea or Concept|Hospital Course|7384,7389|false|false|false|C1546485|Diagnosis Type - Final|final
Event|Event|Hospital Course|7390,7397|false|false|false|||results
Finding|Body Substance|Hospital Course|7406,7412|false|false|false|C1550609|Specimen Type - Abscess|abcess
Drug|Biomedical or Dental Material|Hospital Course|7413,7420|false|false|false|C1706355|Culture Dose Form|culture
Event|Event|Hospital Course|7413,7420|false|false|false|||culture
Finding|Functional Concept|Hospital Course|7413,7420|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Finding|Idea or Concept|Hospital Course|7413,7420|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Procedure|Laboratory Procedure|Hospital Course|7413,7420|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|culture
Event|Event|Hospital Course|7439,7446|false|false|false|||Milleri
Finding|Finding|Hospital Course|7448,7451|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Finding|Idea or Concept|Hospital Course|7448,7451|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Event|Event|Hospital Course|7455,7470|false|false|false|||recommendations
Finding|Idea or Concept|Hospital Course|7455,7470|false|false|false|C0034866|Recommendation|recommendations
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7492,7497|false|false|false|C0042313|vancomycin|Vanco
Drug|Antibiotic|Hospital Course|7492,7497|false|false|false|C0042313|vancomycin|Vanco
Event|Event|Hospital Course|7492,7497|false|false|false|||Vanco
Event|Event|Hospital Course|7502,7511|false|false|false|||Meropenum
Event|Event|Hospital Course|7521,7528|false|false|false|||started
Drug|Antibiotic|Hospital Course|7533,7544|false|false|false|C0007561|ceftriaxone|Ceftriaxone
Drug|Organic Chemical|Hospital Course|7533,7544|false|false|false|C0007561|ceftriaxone|Ceftriaxone
Drug|Organic Chemical|Hospital Course|7561,7567|false|false|false|C0699678|Flagyl|Flagyl
Drug|Pharmacologic Substance|Hospital Course|7561,7567|false|false|false|C0699678|Flagyl|Flagyl
Finding|Body Substance|Hospital Course|7583,7590|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|7583,7590|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|7583,7590|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|7595,7607|false|false|false|||re-evaluated
Event|Event|Hospital Course|7626,7633|false|false|false|||cleared
Event|Event|Hospital Course|7641,7651|false|false|false|||discharged
Event|Event|Hospital Course|7652,7656|false|false|false|||home
Finding|Idea or Concept|Hospital Course|7652,7656|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|7652,7656|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|7652,7656|false|false|false|C1553498|home health encounter|home
Event|Event|Hospital Course|7666,7676|false|false|false|||assistance
Finding|Social Behavior|Hospital Course|7666,7676|false|false|false|C0018896|Helping Behavior|assistance
Event|Event|Hospital Course|7699,7708|false|false|false|||recommend
Event|Event|Hospital Course|7709,7717|false|false|false|||services
Event|Occupational Activity|Hospital Course|7709,7717|false|false|false|C0557854|Services|services
Procedure|Health Care Activity|Hospital Course|7709,7717|false|false|false|C1704289|Clinical Service|services
Finding|Body Substance|Hospital Course|7724,7731|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|7724,7731|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|7724,7731|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|Hospital Course|7735,7742|false|false|false|C4534363|At home|at home
Event|Event|Hospital Course|7738,7742|false|false|false|||home
Finding|Idea or Concept|Hospital Course|7738,7742|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|7738,7742|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|7738,7742|false|false|false|C1553498|home health encounter|home
Event|Event|Hospital Course|7748,7756|false|false|false|||remained
Event|Event|Hospital Course|7757,7763|false|false|false|||stable
Finding|Intellectual Product|Hospital Course|7757,7763|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Activity|Hospital Course|7768,7779|false|false|false|C4321457|Examination|examination
Event|Event|Hospital Course|7768,7779|false|false|false|||examination
Procedure|Health Care Activity|Hospital Course|7768,7779|false|false|false|C0031809;C0582103|Medical Examination;Physical Examination|examination
Event|Event|Hospital Course|7803,7807|false|false|false|||seen
Event|Event|Hospital Course|7812,7821|false|false|false|||evaluated
Event|Event|Hospital Course|7828,7838|false|false|false|||complained
Event|Event|Hospital Course|7842,7850|false|false|false|||headache
Finding|Sign or Symptom|Hospital Course|7842,7850|false|false|false|C0018681|Headache|headache
Anatomy|Body Location or Region|Hospital Course|7870,7874|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7870,7874|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|Hospital Course|7870,7874|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7870,7874|false|false|false|C0876917|Procedure on head|head
Procedure|Diagnostic Procedure|Hospital Course|7870,7877|false|false|false|C0202691|CAT scan of head|head CT
Event|Event|Hospital Course|7875,7877|false|false|false|||CT
Event|Event|Hospital Course|7882,7889|false|false|false|||ordered
Event|Event|Hospital Course|7897,7903|false|false|false|||showed
Finding|Intellectual Product|Hospital Course|7908,7914|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|Hospital Course|7930,7937|false|false|false|||changes
Finding|Functional Concept|Hospital Course|7930,7937|false|false|false|C0392747|Changing|changes
Finding|Idea or Concept|Hospital Course|7940,7944|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|7940,7944|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|7940,7944|false|false|false|C1553498|home health encounter|Home
Procedure|Health Care Activity|Hospital Course|7940,7953|false|false|false|C0020043|Home visit (procedure)|Home services
Event|Event|Hospital Course|7945,7953|false|false|false|||services
Event|Occupational Activity|Hospital Course|7945,7953|false|false|false|C0557854|Services|services
Procedure|Health Care Activity|Hospital Course|7945,7953|false|false|false|C1704289|Clinical Service|services
Event|Event|Hospital Course|7960,7971|false|false|false|||established
Finding|Body Substance|Hospital Course|7980,7987|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|7980,7987|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|7980,7987|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|7992,8002|false|false|false|||discharged
Attribute|Clinical Attribute|Hospital Course|8007,8018|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|8007,8018|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|8007,8018|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|8007,8018|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|8007,8031|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|8022,8031|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|8022,8031|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Organic Chemical|Hospital Course|8033,8042|false|false|false|C0020740|ibuprofen|Ibuprofen
Drug|Pharmacologic Substance|Hospital Course|8033,8042|false|false|false|C0020740|ibuprofen|Ibuprofen
Event|Event|Hospital Course|8045,8054|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|8045,8054|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|8045,8054|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|8045,8054|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|8045,8054|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|8045,8066|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|8055,8066|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|8055,8066|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|8055,8066|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|8055,8066|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|8071,8084|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|8071,8084|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Hospital Course|8071,8084|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|8071,8084|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|Hospital Course|8103,8106|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|8107,8111|false|false|false|C2598155||pain
Event|Event|Hospital Course|8107,8111|false|false|false|||pain
Finding|Functional Concept|Hospital Course|8107,8111|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|8107,8111|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|8117,8130|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Drug|Pharmacologic Substance|Hospital Course|8117,8130|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Event|Event|Hospital Course|8117,8130|false|false|false|||acetaminophen
Procedure|Laboratory Procedure|Hospital Course|8117,8130|false|false|false|C0373527|Acetaminophen measurement|acetaminophen
Drug|Biomedical or Dental Material|Hospital Course|8142,8148|false|false|false|C0039225|Tablet Dosage Form|tablet
Event|Event|Hospital Course|8142,8148|false|false|false|||tablet
Finding|Functional Concept|Hospital Course|8152,8160|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|8155,8160|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|8155,8160|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Biomedical or Dental Material|Hospital Course|8193,8199|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|8200,8207|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|8200,8207|false|false|false|C0807726|refill|Refills
Drug|Antibiotic|Hospital Course|8214,8225|false|false|false|C0007561|ceftriaxone|CeftriaXONE
Drug|Organic Chemical|Hospital Course|8214,8225|false|false|false|C0007561|ceftriaxone|CeftriaXONE
Event|Event|Hospital Course|8240,8242|false|false|false|||RX
Drug|Antibiotic|Hospital Course|8244,8255|false|false|false|C0007561|ceftriaxone|ceftriaxone
Drug|Organic Chemical|Hospital Course|8244,8255|false|false|false|C0007561|ceftriaxone|ceftriaxone
Event|Event|Hospital Course|8244,8255|false|false|false|||ceftriaxone
Event|Event|Hospital Course|8311,8318|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|8311,8318|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|8325,8333|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|8325,8333|false|false|false|C1692318|docusate|Docusate
Event|Event|Hospital Course|8325,8333|false|false|false|||Docusate
Drug|Organic Chemical|Hospital Course|8325,8340|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|Hospital Course|8325,8340|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|Hospital Course|8334,8340|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|8334,8340|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|8334,8340|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|8334,8340|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|8334,8340|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|8334,8340|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8351,8354|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8351,8354|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8351,8354|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|8351,8354|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|8351,8354|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|8360,8368|false|false|false|C1692318|docusate|docusate
Drug|Pharmacologic Substance|Hospital Course|8360,8368|false|false|false|C1692318|docusate|docusate
Drug|Organic Chemical|Hospital Course|8360,8375|false|false|false|C0243237|docusate sodium|docusate sodium
Drug|Pharmacologic Substance|Hospital Course|8360,8375|false|false|false|C0243237|docusate sodium|docusate sodium
Drug|Biologically Active Substance|Hospital Course|8369,8375|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|Hospital Course|8369,8375|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|Hospital Course|8369,8375|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Event|Event|Hospital Course|8369,8375|false|false|false|||sodium
Finding|Physiologic Function|Hospital Course|8369,8375|false|false|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|Hospital Course|8369,8375|false|false|false|C0337443|Sodium measurement|sodium
Drug|Organic Chemical|Hospital Course|8377,8383|false|false|false|C0282139|Colace|Colace
Drug|Pharmacologic Substance|Hospital Course|8377,8383|false|false|false|C0282139|Colace|Colace
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8394,8401|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|Hospital Course|8394,8401|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|Hospital Course|8394,8401|false|false|false|C0006935|capsule (pharmacologic)|capsule
Finding|Functional Concept|Hospital Course|8405,8413|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|8408,8413|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|8408,8413|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|Hospital Course|8423,8426|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|8423,8426|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8437,8444|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|8437,8444|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|8437,8444|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Event|Event|Hospital Course|8445,8452|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|8445,8452|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|8459,8472|false|false|false|C0377265|levetiracetam|LeVETiracetam
Drug|Pharmacologic Substance|Hospital Course|8459,8472|false|false|false|C0377265|levetiracetam|LeVETiracetam
Event|Event|Hospital Course|8459,8472|false|false|false|||LeVETiracetam
Procedure|Laboratory Procedure|Hospital Course|8459,8472|false|false|false|C3693636|Measurement of levetiracetam|LeVETiracetam
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8484,8487|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8484,8487|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8484,8487|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|8484,8487|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|8484,8487|false|false|false|C1332410|BID gene|BID
Event|Event|Hospital Course|8489,8491|false|false|false|||RX
Drug|Organic Chemical|Hospital Course|8493,8506|false|false|false|C0377265|levetiracetam|levetiracetam
Drug|Pharmacologic Substance|Hospital Course|8493,8506|false|false|false|C0377265|levetiracetam|levetiracetam
Event|Event|Hospital Course|8493,8506|false|false|false|||levetiracetam
Procedure|Laboratory Procedure|Hospital Course|8493,8506|false|false|false|C3693636|Measurement of levetiracetam|levetiracetam
Drug|Organic Chemical|Hospital Course|8508,8514|false|false|false|C0876060|Keppra|Keppra
Drug|Pharmacologic Substance|Hospital Course|8508,8514|false|false|false|C0876060|Keppra|Keppra
Drug|Biomedical or Dental Material|Hospital Course|8527,8533|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|8537,8545|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|8540,8545|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|8540,8545|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|Hospital Course|8555,8558|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|8555,8558|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biomedical or Dental Material|Hospital Course|8569,8575|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|8576,8583|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|8576,8583|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|8590,8603|true|false|false|C0025872|metronidazole|MetRONIDAZOLE
Drug|Pharmacologic Substance|Hospital Course|8590,8603|true|false|false|C0025872|metronidazole|MetRONIDAZOLE
Drug|Organic Chemical|Hospital Course|8605,8611|false|false|false|C0699678|Flagyl|FLagyl
Drug|Pharmacologic Substance|Hospital Course|8605,8611|false|false|false|C0699678|Flagyl|FLagyl
Event|Event|Hospital Course|8623,8626|false|false|false|||TID
Event|Event|Hospital Course|8628,8630|false|false|false|||RX
Drug|Organic Chemical|Hospital Course|8632,8645|false|false|false|C0025872|metronidazole|metronidazole
Drug|Pharmacologic Substance|Hospital Course|8632,8645|false|false|false|C0025872|metronidazole|metronidazole
Event|Event|Hospital Course|8632,8645|false|false|false|||metronidazole
Drug|Organic Chemical|Hospital Course|8647,8653|false|false|false|C0699678|Flagyl|Flagyl
Drug|Pharmacologic Substance|Hospital Course|8647,8653|false|false|false|C0699678|Flagyl|Flagyl
Drug|Biomedical or Dental Material|Hospital Course|8664,8670|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|8674,8682|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|8677,8682|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|8677,8682|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Disorder|Disease or Syndrome|Hospital Course|8690,8695|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|Hospital Course|8698,8701|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|8698,8701|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biomedical or Dental Material|Hospital Course|8713,8719|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|8720,8727|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|8720,8727|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|8734,8743|false|false|false|C0030049|oxycodone|OxycoDONE
Drug|Pharmacologic Substance|Hospital Course|8734,8743|false|false|false|C0030049|oxycodone|OxycoDONE
Event|Event|Hospital Course|8734,8743|false|false|false|||OxycoDONE
Procedure|Laboratory Procedure|Hospital Course|8734,8743|false|false|false|C0524222|Oxycodone measurement|OxycoDONE
Finding|Idea or Concept|Hospital Course|8745,8754|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Finding|Intellectual Product|Hospital Course|8745,8754|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Drug|Biomedical or Dental Material|Hospital Course|8745,8762|false|false|false|C1708470|Immediate Release Dosage Form|Immediate Release
Event|Event|Hospital Course|8755,8762|false|false|false|||Release
Finding|Functional Concept|Hospital Course|8755,8762|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|8755,8762|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8755,8762|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Finding|Gene or Genome|Hospital Course|8777,8780|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|8781,8785|false|false|false|C2598155||pain
Event|Event|Hospital Course|8781,8785|false|false|false|||pain
Finding|Functional Concept|Hospital Course|8781,8785|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|8781,8785|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|8787,8789|false|false|false|||RX
Drug|Organic Chemical|Hospital Course|8791,8800|false|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|Hospital Course|8791,8800|false|false|false|C0030049|oxycodone|oxycodone
Event|Event|Hospital Course|8791,8800|false|false|false|||oxycodone
Procedure|Laboratory Procedure|Hospital Course|8791,8800|false|false|false|C0524222|Oxycodone measurement|oxycodone
Drug|Organic Chemical|Hospital Course|8802,8808|false|false|false|C3160522|Oxecta|Oxecta
Drug|Pharmacologic Substance|Hospital Course|8802,8808|false|false|false|C3160522|Oxecta|Oxecta
Event|Event|Hospital Course|8802,8808|false|false|false|||Oxecta
Drug|Biomedical or Dental Material|Hospital Course|8817,8823|false|false|false|C0039225|Tablet Dosage Form|tablet
Event|Event|Hospital Course|8817,8823|false|false|false|||tablet
Drug|Biomedical or Dental Material|Hospital Course|8817,8834|false|false|false|C3473439|TABLET, ORAL ONLY|tablet, oral only
Anatomy|Body Space or Junction|Hospital Course|8825,8829|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|8825,8829|false|false|false|C1272919|Oral Dosage Form|oral
Event|Event|Hospital Course|8825,8829|false|false|false|||oral
Finding|Finding|Hospital Course|8825,8829|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|8825,8829|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|8838,8846|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|8841,8846|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|8841,8846|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Biomedical or Dental Material|Hospital Course|8879,8885|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|8886,8893|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|8886,8893|false|false|false|C0807726|refill|Refills
Drug|Biologically Active Substance|Hospital Course|8900,8907|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Drug|Organic Chemical|Hospital Course|8900,8907|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Drug|Pharmacologic Substance|Hospital Course|8900,8907|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Drug|Organic Chemical|Hospital Course|8900,8913|false|false|false|C0354589|heparin flush|Heparin Flush
Drug|Pharmacologic Substance|Hospital Course|8900,8913|false|false|false|C0354589|heparin flush|Heparin Flush
Event|Event|Hospital Course|8908,8913|false|false|false|||Flush
Finding|Functional Concept|Hospital Course|8908,8913|false|false|false|C0016382;C1696091|Flush - RouteOfAdministration;Flushing|Flush
Finding|Sign or Symptom|Hospital Course|8908,8913|false|false|false|C0016382;C1696091|Flush - RouteOfAdministration;Flushing|Flush
Disorder|Disease or Syndrome|Hospital Course|8930,8935|false|false|false|C0238286|Mucolipidosis Type IV|mL IV
Finding|Gene or Genome|Hospital Course|8946,8949|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Biologically Active Substance|Hospital Course|8951,8955|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Hospital Course|8951,8955|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Substance|Hospital Course|8951,8955|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Finding|Intellectual Product|Hospital Course|8951,8955|false|false|false|C1546701|line source specimen code|line
Attribute|Clinical Attribute|Hospital Course|8951,8961|false|false|false|C4036660||line flush
Event|Event|Hospital Course|8956,8961|false|false|false|||flush
Finding|Functional Concept|Hospital Course|8956,8961|false|false|false|C0016382;C1696091|Flush - RouteOfAdministration;Flushing|flush
Finding|Sign or Symptom|Hospital Course|8956,8961|false|false|false|C0016382;C1696091|Flush - RouteOfAdministration;Flushing|flush
Drug|Biologically Active Substance|Hospital Course|8968,8975|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|Hospital Course|8968,8975|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|Hospital Course|8968,8975|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|Hospital Course|8968,8986|false|false|false|C0720846|Heparin Lock Flush|heparin lock flush
Drug|Pharmacologic Substance|Hospital Course|8968,8986|false|false|false|C0720846|Heparin Lock Flush|heparin lock flush
Finding|Idea or Concept|Hospital Course|8976,8980|false|false|false|C1550024|Lock - Remote control command|lock
Event|Event|Hospital Course|8981,8986|false|false|false|||flush
Finding|Functional Concept|Hospital Course|8981,8986|false|false|false|C0016382;C1696091|Flush - RouteOfAdministration;Flushing|flush
Finding|Sign or Symptom|Hospital Course|8981,8986|false|false|false|C0016382;C1696091|Flush - RouteOfAdministration;Flushing|flush
Event|Event|Hospital Course|8988,8995|false|false|false|||porcine
Finding|Finding|Hospital Course|8988,8995|false|false|false|C4554819|Porcine prosthetic valve|porcine
Drug|Biologically Active Substance|Hospital Course|8998,9005|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|Hospital Course|8998,9005|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|Hospital Course|8998,9005|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|Hospital Course|8998,9016|false|false|false|C0720846|Heparin Lock Flush|heparin lock flush
Drug|Pharmacologic Substance|Hospital Course|8998,9016|false|false|false|C0720846|Heparin Lock Flush|heparin lock flush
Finding|Idea or Concept|Hospital Course|9006,9010|false|false|false|C1550024|Lock - Remote control command|lock
Event|Event|Hospital Course|9011,9016|false|false|false|||flush
Finding|Functional Concept|Hospital Course|9011,9016|false|false|false|C0016382;C1696091|Flush - RouteOfAdministration;Flushing|flush
Finding|Sign or Symptom|Hospital Course|9011,9016|false|false|false|C0016382;C1696091|Flush - RouteOfAdministration;Flushing|flush
Disorder|Disease or Syndrome|Hospital Course|9032,9037|false|false|false|C0238286|Mucolipidosis Type IV|ml IV
Event|Event|Hospital Course|9076,9083|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|9076,9083|false|false|false|C0807726|refill|Refills
Drug|Biologically Active Substance|Hospital Course|9090,9096|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|9090,9096|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|9090,9096|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|9090,9096|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|9090,9096|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|9090,9096|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Inorganic Chemical|Hospital Course|9090,9105|false|false|false|C0037494|sodium chloride|Sodium Chloride
Drug|Element, Ion, or Isotope|Hospital Course|9097,9105|false|false|false|C0008203;C0596019|Chlorides;chloride ion|Chloride
Event|Event|Hospital Course|9097,9105|false|false|false|||Chloride
Finding|Physiologic Function|Hospital Course|9097,9105|false|false|false|C4553021|Chloride metabolic function|Chloride
Procedure|Laboratory Procedure|Hospital Course|9097,9105|false|false|false|C0201952|Chloride measurement|Chloride
Event|Event|Hospital Course|9112,9117|false|false|false|||Flush
Finding|Functional Concept|Hospital Course|9112,9117|false|false|false|C0016382;C1696091|Flush - RouteOfAdministration;Flushing|Flush
Finding|Sign or Symptom|Hospital Course|9112,9117|false|false|false|C0016382;C1696091|Flush - RouteOfAdministration;Flushing|Flush
Disorder|Disease or Syndrome|Hospital Course|9121,9126|false|false|false|C0238286|Mucolipidosis Type IV|mL IV
Finding|Gene or Genome|Hospital Course|9135,9138|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Biologically Active Substance|Hospital Course|9140,9144|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Hospital Course|9140,9144|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Substance|Hospital Course|9140,9144|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Finding|Intellectual Product|Hospital Course|9140,9144|false|false|false|C1546701|line source specimen code|line
Attribute|Clinical Attribute|Hospital Course|9140,9150|false|false|false|C4036660||line flush
Event|Event|Hospital Course|9145,9150|false|false|false|||flush
Finding|Functional Concept|Hospital Course|9145,9150|false|false|false|C0016382;C1696091|Flush - RouteOfAdministration;Flushing|flush
Finding|Sign or Symptom|Hospital Course|9145,9150|false|false|false|C0016382;C1696091|Flush - RouteOfAdministration;Flushing|flush
Event|Event|Hospital Course|9152,9157|false|false|false|||Flush
Finding|Functional Concept|Hospital Course|9152,9157|false|false|false|C0016382;C1696091|Flush - RouteOfAdministration;Flushing|Flush
Finding|Sign or Symptom|Hospital Course|9152,9157|false|false|false|C0016382;C1696091|Flush - RouteOfAdministration;Flushing|Flush
Event|Event|Hospital Course|9180,9188|false|false|false|||infusion
Finding|Functional Concept|Hospital Course|9180,9188|false|false|false|C1827465|Infusion route|infusion
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9180,9188|false|false|false|C0574032|Infusion procedures|infusion
Drug|Antibiotic|Hospital Course|9192,9203|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|Hospital Course|9192,9203|false|false|false|||antibiotics
Drug|Biologically Active Substance|Hospital Course|9210,9216|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|Hospital Course|9210,9216|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|Hospital Course|9210,9216|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Finding|Physiologic Function|Hospital Course|9210,9216|false|false|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|Hospital Course|9210,9216|false|false|false|C0337443|Sodium measurement|sodium
Drug|Inorganic Chemical|Hospital Course|9210,9225|false|false|false|C0037494|sodium chloride|sodium chloride
Drug|Element, Ion, or Isotope|Hospital Course|9217,9225|false|false|false|C0008203;C0596019|Chlorides;chloride ion|chloride
Event|Event|Hospital Course|9217,9225|false|false|false|||chloride
Finding|Physiologic Function|Hospital Course|9217,9225|false|false|false|C4553021|Chloride metabolic function|chloride
Procedure|Laboratory Procedure|Hospital Course|9217,9225|false|false|false|C0201952|Chloride measurement|chloride
Drug|Inorganic Chemical|Hospital Course|9240,9246|false|false|false|C0036082|Saline Solution|Saline
Drug|Pharmacologic Substance|Hospital Course|9240,9246|false|false|false|C0036082|Saline Solution|Saline
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9240,9246|false|false|false|C0450082|Saline method|Saline
Event|Event|Hospital Course|9240,9252|false|false|false|||Saline Flush
Procedure|Health Care Activity|Hospital Course|9240,9252|false|false|false|C3828271|Saline Flush|Saline Flush
Finding|Functional Concept|Hospital Course|9247,9252|false|false|false|C0016382;C1696091|Flush - RouteOfAdministration;Flushing|Flush
Finding|Sign or Symptom|Hospital Course|9247,9252|false|false|false|C0016382;C1696091|Flush - RouteOfAdministration;Flushing|Flush
Disorder|Disease or Syndrome|Hospital Course|9263,9268|false|false|false|C0238286|Mucolipidosis Type IV|ml IV
Event|Event|Hospital Course|9270,9273|false|false|false|||q12
Event|Event|Hospital Course|9293,9300|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|9293,9300|false|false|false|C0807726|refill|Refills
Event|Event|Hospital Course|9307,9316|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|9307,9316|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|9307,9316|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|9307,9316|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|9307,9316|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|9307,9328|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|9307,9328|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|9317,9328|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|9317,9328|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|9317,9328|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|Hospital Course|9330,9334|false|false|false|||Home
Finding|Idea or Concept|Hospital Course|9330,9334|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|9330,9334|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|9330,9334|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|Hospital Course|9340,9347|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|Hospital Course|9340,9347|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|Hospital Course|9350,9358|false|false|false|||Facility
Finding|Intellectual Product|Hospital Course|9350,9358|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|Hospital Course|9366,9375|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|9366,9375|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|9366,9375|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|9366,9375|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|9366,9375|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|9366,9385|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|9376,9385|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|9376,9385|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|9376,9385|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|9376,9385|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|9376,9385|false|false|false|C0011900|Diagnosis|Diagnosis
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9387,9392|false|false|false|C0006104;C4266577|Brain;Head>Brain|Brain
Disorder|Disease or Syndrome|Hospital Course|9387,9392|false|false|false|C0006111|Brain Diseases|Brain
Disorder|Disease or Syndrome|Hospital Course|9387,9400|false|false|false|C0006105;C1510428|Brain Abscess;Cerebral abscess|Brain abscess
Disorder|Disease or Syndrome|Hospital Course|9393,9400|false|false|false|C0000833|Abscess|abscess
Event|Event|Hospital Course|9393,9400|false|false|false|||abscess
Finding|Intellectual Product|Hospital Course|9393,9400|false|false|false|C1546533||abscess
Finding|Mental Process|Discharge Condition|9425,9431|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|9425,9438|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|9425,9438|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|9432,9438|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|9432,9438|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|9440,9445|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|9440,9445|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|9450,9458|false|false|false|||coherent
Finding|Finding|Discharge Condition|9450,9458|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|9460,9465|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|9460,9482|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|9460,9482|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|9469,9482|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|9469,9482|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|9469,9482|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|9484,9489|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|9484,9489|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|9484,9489|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|9484,9489|false|false|false|||Alert
Finding|Finding|Discharge Condition|9484,9489|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|9484,9489|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|9484,9489|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|9494,9505|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|9494,9505|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|9507,9515|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|9507,9515|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|9507,9515|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|9516,9522|false|false|false|C5889824||Status
Event|Event|Discharge Condition|9516,9522|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|9516,9522|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|Discharge Condition|9524,9534|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|9524,9534|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|9524,9534|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|9524,9534|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|9537,9545|false|false|false|||requires
Event|Event|Discharge Condition|9546,9556|false|false|false|||assistance
Finding|Social Behavior|Discharge Condition|9546,9556|false|false|false|C0018896|Helping Behavior|assistance
Drug|Amino Acid, Peptide, or Protein|Discharge Condition|9560,9563|false|false|false|C1454018|AICDA protein, human|aid
Drug|Enzyme|Discharge Condition|9560,9563|false|false|false|C1454018|AICDA protein, human|aid
Event|Event|Discharge Condition|9560,9563|false|false|false|||aid
Finding|Gene or Genome|Discharge Condition|9560,9563|false|false|false|C1421876;C3540469|AICDA gene;AICDA wt Allele|aid
Procedure|Therapeutic or Preventive Procedure|Discharge Condition|9560,9563|false|false|false|C0021588;C0280108|AID - Artificial insemination by donor;dacarbazine/doxorubicin/ifosfamide protocol|aid
Event|Event|Discharge Condition|9565,9571|false|false|false|||walker
Event|Event|Discharge Instructions|9618,9624|false|false|false|||friend
Finding|Idea or Concept|Discharge Instructions|9618,9624|false|false|false|C1546502|Relationship - Friend|friend
Finding|Classification|Discharge Instructions|9625,9631|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Discharge Instructions|9625,9631|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Discharge Instructions|9625,9631|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Discharge Instructions|9625,9631|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Event|Event|Discharge Instructions|9639,9644|false|false|false|||check
Anatomy|Body Location or Region|Discharge Instructions|9650,9658|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Discharge Instructions|9650,9658|false|false|false|C0332803|Surgical wound|incision
Event|Event|Discharge Instructions|9650,9658|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|9650,9658|false|false|false|C0184898|Surgical incisions|incision
Event|Event|Discharge Instructions|9670,9675|false|false|false|||signs
Finding|Finding|Discharge Instructions|9670,9675|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Discharge Instructions|9670,9675|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Disorder|Disease or Syndrome|Discharge Instructions|9679,9688|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|Discharge Instructions|9679,9688|false|false|false|||infection
Finding|Pathologic Function|Discharge Instructions|9679,9688|false|false|false|C3714514|Infection|infection
Event|Event|Discharge Instructions|9691,9695|false|false|false|||Take
Attribute|Clinical Attribute|Discharge Instructions|9701,9705|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|9701,9705|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|9701,9705|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|9701,9705|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Hazardous or Poisonous Substance|Discharge Instructions|9701,9714|false|false|false|C0002771|Analgesics|pain medicine
Drug|Organic Chemical|Discharge Instructions|9701,9714|false|false|false|C0002771|Analgesics|pain medicine
Drug|Pharmacologic Substance|Discharge Instructions|9701,9714|false|false|false|C0002771|Analgesics|pain medicine
Drug|Pharmacologic Substance|Discharge Instructions|9706,9714|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Event|Event|Discharge Instructions|9706,9714|false|false|false|||medicine
Event|Event|Discharge Instructions|9718,9728|false|false|false|||prescribed
Event|Event|Discharge Instructions|9731,9739|false|false|false|||Exercise
Finding|Daily or Recreational Activity|Discharge Instructions|9731,9739|false|false|false|C0015259|Exercise|Exercise
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|9731,9739|false|false|false|C1522704|Exercise Pain Management|Exercise
Event|Event|Discharge Instructions|9750,9757|false|false|false|||limited
Event|Event|Discharge Instructions|9761,9768|false|false|false|||walking
Finding|Daily or Recreational Activity|Discharge Instructions|9761,9768|false|true|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Finding|Finding|Discharge Instructions|9761,9768|false|true|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Finding|Sign or Symptom|Discharge Instructions|9761,9768|false|true|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Event|Activity|Discharge Instructions|9773,9780|true|false|false|C0206244|Lifting|lifting
Event|Event|Discharge Instructions|9773,9780|true|false|false|||lifting
Event|Event|Discharge Instructions|9782,9791|true|false|false|||straining
Finding|Physiologic Function|Discharge Instructions|9782,9791|true|false|false|C0442694|Straining (finding)|straining
Disorder|Disease or Syndrome|Discharge Instructions|9807,9814|false|false|false|C0011119|Decompression Sickness|bending
Event|Event|Discharge Instructions|9807,9814|false|false|false|||bending
Finding|Finding|Discharge Instructions|9807,9814|false|false|false|C0700231;C2584296|Bending - Changing basic body position;Does bend|bending
Finding|Physiologic Function|Discharge Instructions|9807,9814|false|false|false|C0700231;C2584296|Bending - Changing basic body position;Does bend|bending
Disorder|Injury or Poisoning|Discharge Instructions|9824,9829|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Event|Event|Discharge Instructions|9824,9829|false|false|false|||wound
Finding|Body Substance|Discharge Instructions|9824,9829|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|Discharge Instructions|9824,9829|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|Discharge Instructions|9824,9829|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Event|Event|Discharge Instructions|9834,9840|false|false|false|||closed
Anatomy|Body Space or Junction|Discharge Instructions|9846,9853|false|false|false|C0502420|Suture Joint|sutures
Event|Event|Discharge Instructions|9863,9867|false|false|false|||wash
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|9873,9877|false|false|false|C0018494|Hair|hair
Finding|Body Substance|Discharge Instructions|9873,9877|false|false|false|C0444095;C1546660|Hair Specimen;Hair Specimen Code|hair
Finding|Intellectual Product|Discharge Instructions|9873,9877|false|false|false|C0444095;C1546660|Hair Specimen;Hair Specimen Code|hair
Anatomy|Body Space or Junction|Discharge Instructions|9890,9897|false|false|false|C0502420|Suture Joint|sutures
Event|Event|Discharge Instructions|9905,9912|false|false|false|||staples
Event|Event|Discharge Instructions|9923,9930|false|false|false|||removed
Event|Event|Discharge Instructions|9942,9948|false|false|false|||shower
Finding|Finding|Discharge Instructions|9961,9965|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Discharge Instructions|9961,9965|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Discharge Instructions|9961,9965|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Disorder|Congenital Abnormality|Discharge Instructions|9981,9984|false|true|false|C1855179|CATARACT, ANTERIOR POLAR|cap
Drug|Biomedical or Dental Material|Discharge Instructions|9981,9984|false|true|false|C0006935|capsule (pharmacologic)|cap
Event|Event|Discharge Instructions|9981,9984|false|false|false|||cap
Finding|Gene or Genome|Discharge Instructions|9981,9984|false|true|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|cap
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|9981,9984|false|true|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|cap
Event|Event|Discharge Instructions|9988,9993|false|false|false|||cover
Finding|Functional Concept|Discharge Instructions|9988,9993|false|false|false|C1999244||cover
Anatomy|Body Location or Region|Discharge Instructions|10000,10004|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|10000,10004|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|Discharge Instructions|10000,10004|false|false|false|C0362076|Problems with head|head
Event|Event|Discharge Instructions|10000,10004|false|false|false|||head
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10000,10004|false|false|false|C0876917|Procedure on head|head
Event|Event|Discharge Instructions|10007,10015|false|false|false|||Increase
Event|Event|Discharge Instructions|10021,10027|false|false|false|||intake
Finding|Functional Concept|Discharge Instructions|10021,10027|false|false|false|C1512806|Intake|intake
Procedure|Health Care Activity|Discharge Instructions|10021,10027|false|false|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|intake
Drug|Substance|Discharge Instructions|10031,10037|false|false|false|C0302908|Liquid substance|fluids
Event|Event|Discharge Instructions|10031,10037|false|false|false|||fluids
Finding|Body Substance|Discharge Instructions|10031,10037|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10031,10037|false|false|false|C0016286|Fluid Therapy|fluids
Anatomy|Tissue|Discharge Instructions|10042,10047|false|false|false|C1304649|Tissue fiber|fiber
Drug|Organic Chemical|Discharge Instructions|10042,10047|false|false|false|C0225326;C1321801|Fiber brand of calcium polycarbophil;fiber|fiber
Drug|Pharmacologic Substance|Discharge Instructions|10042,10047|false|false|false|C0225326;C1321801|Fiber brand of calcium polycarbophil;fiber|fiber
Drug|Hazardous or Poisonous Substance|Discharge Instructions|10052,10060|false|false|false|C0027415|Narcotics|narcotic
Drug|Pharmacologic Substance|Discharge Instructions|10052,10060|false|false|false|C0027415|Narcotics|narcotic
Attribute|Clinical Attribute|Discharge Instructions|10061,10065|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|10061,10065|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|10061,10065|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|10061,10065|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Pharmacologic Substance|Discharge Instructions|10067,10075|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Event|Event|Discharge Instructions|10067,10075|false|false|false|||medicine
Event|Event|Discharge Instructions|10080,10085|false|false|false|||cause
Event|Event|Discharge Instructions|10086,10098|false|false|false|||constipation
Finding|Sign or Symptom|Discharge Instructions|10086,10098|false|false|false|C0009806|Constipation|constipation
Event|Event|Discharge Instructions|10113,10122|false|false|false|||recommend
Event|Event|Discharge Instructions|10123,10129|false|false|false|||taking
Drug|Pharmacologic Substance|Discharge Instructions|10134,10150|false|false|false|C0013231|Drugs, Non-Prescription|over the counter
Drug|Hazardous or Poisonous Substance|Discharge Instructions|10143,10150|false|false|false|C0702263|Counter brand of Terbufos|counter
Drug|Organic Chemical|Discharge Instructions|10143,10150|false|false|false|C0702263|Counter brand of Terbufos|counter
Finding|Body Substance|Discharge Instructions|10151,10156|false|false|false|C0015733|Feces|stool
Drug|Organic Chemical|Discharge Instructions|10151,10165|false|false|false|C0301470;C1154263|Stool Softener;Stool Softener brand of docusate sodium|stool softener
Drug|Pharmacologic Substance|Discharge Instructions|10151,10165|false|false|false|C0301470;C1154263|Stool Softener;Stool Softener brand of docusate sodium|stool softener
Event|Event|Discharge Instructions|10157,10165|false|false|false|||softener
Drug|Organic Chemical|Discharge Instructions|10175,10183|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Discharge Instructions|10175,10183|false|false|false|C1692318|docusate|Docusate
Drug|Organic Chemical|Discharge Instructions|10185,10191|false|false|false|C0282139|Colace|Colace
Drug|Pharmacologic Substance|Discharge Instructions|10185,10191|false|false|false|C0282139|Colace|Colace
Drug|Hazardous or Poisonous Substance|Discharge Instructions|10207,10215|false|false|false|C0027415|Narcotics|narcotic
Drug|Pharmacologic Substance|Discharge Instructions|10207,10215|false|false|false|C0027415|Narcotics|narcotic
Attribute|Clinical Attribute|Discharge Instructions|10216,10220|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|10216,10220|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|10216,10220|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|10216,10220|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Pharmacologic Substance|Discharge Instructions|10221,10231|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Discharge Instructions|10221,10231|false|false|false|||medication
Finding|Intellectual Product|Discharge Instructions|10221,10231|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Discharge Instructions|10241,10249|true|false|false|||directed
Event|Event|Discharge Instructions|10258,10264|true|false|false|||doctor
Finding|Intellectual Product|Discharge Instructions|10258,10264|true|false|false|C2348314|Doctor - Title|doctor
Event|Event|Discharge Instructions|10273,10277|true|false|false|||take
Drug|Pharmacologic Substance|Discharge Instructions|10283,10300|true|false|false|C0003209|Anti-Inflammatory Agents|anti-inflammatory
Drug|Pharmacologic Substance|Discharge Instructions|10301,10310|true|false|false|C0013227|Pharmaceutical Preparations|medicines
Event|Event|Discharge Instructions|10301,10310|true|false|false|||medicines
Drug|Organic Chemical|Discharge Instructions|10319,10325|true|false|false|C0699203|Motrin|Motrin
Drug|Pharmacologic Substance|Discharge Instructions|10319,10325|true|false|false|C0699203|Motrin|Motrin
Drug|Organic Chemical|Discharge Instructions|10327,10334|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Discharge Instructions|10327,10334|false|false|false|C0004057|aspirin|Aspirin
Event|Event|Discharge Instructions|10327,10334|false|false|false|||Aspirin
Drug|Organic Chemical|Discharge Instructions|10336,10341|false|false|false|C0593507|Advil|Advil
Drug|Pharmacologic Substance|Discharge Instructions|10336,10341|false|false|false|C0593507|Advil|Advil
Event|Event|Discharge Instructions|10336,10341|false|false|false|||Advil
Finding|Gene or Genome|Discharge Instructions|10336,10341|false|false|false|C1422473|AVIL gene|Advil
Drug|Organic Chemical|Discharge Instructions|10348,10357|false|false|false|C0020740|ibuprofen|Ibuprofen
Drug|Pharmacologic Substance|Discharge Instructions|10348,10357|false|false|false|C0020740|ibuprofen|Ibuprofen
Finding|Idea or Concept|Discharge Instructions|10358,10361|false|false|false|C1548556|Etc.|etc
Event|Event|Discharge Instructions|10379,10389|false|false|false|||discharged
Drug|Organic Chemical|Discharge Instructions|10393,10399|false|false|false|C0876060|Keppra|Keppra
Drug|Pharmacologic Substance|Discharge Instructions|10393,10399|false|false|false|C0876060|Keppra|Keppra
Drug|Organic Chemical|Discharge Instructions|10401,10414|false|false|false|C0377265|levetiracetam|Levetiracetam
Drug|Pharmacologic Substance|Discharge Instructions|10401,10414|false|false|false|C0377265|levetiracetam|Levetiracetam
Event|Event|Discharge Instructions|10401,10414|false|false|false|||Levetiracetam
Procedure|Laboratory Procedure|Discharge Instructions|10401,10414|false|false|false|C3693636|Measurement of levetiracetam|Levetiracetam
Event|Event|Discharge Instructions|10431,10438|true|false|false|||require
Disorder|Disease or Syndrome|Discharge Instructions|10439,10444|true|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Discharge Instructions|10439,10444|true|false|false|||blood
Finding|Body Substance|Discharge Instructions|10439,10444|true|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Occupational Activity|Discharge Instructions|10445,10449|true|false|false|C0043227|Work|work
Event|Activity|Discharge Instructions|10450,10460|true|false|false|C1283169||monitoring
Event|Event|Discharge Instructions|10450,10460|true|false|false|||monitoring
Procedure|Health Care Activity|Discharge Instructions|10450,10460|true|false|false|C0150369|Preventive monitoring|monitoring
Event|Event|Discharge Instructions|10462,10463|false|false|false|||
Attribute|Clinical Attribute|Discharge Instructions|10463,10472|false|false|false|C1382187|Clearance of substance|Clearance
Event|Event|Discharge Instructions|10463,10472|false|false|false|||Clearance
Phenomenon|Natural Phenomenon or Process|Discharge Instructions|10463,10472|false|false|false|C2825073|Clearance [PK]|Clearance
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10463,10472|false|false|false|C4554548|Clearance procedure|Clearance
Event|Event|Discharge Instructions|10476,10481|false|false|false|||drive
Event|Event|Discharge Instructions|10486,10492|false|false|false|||return
Event|Occupational Activity|Discharge Instructions|10496,10500|false|false|false|C0043227|Work|work
Event|Event|Discharge Instructions|10509,10518|false|false|false|||addressed
Finding|Idea or Concept|Discharge Instructions|10543,10549|false|false|false|C1549636|Address type - Office|office
Procedure|Health Care Activity|Discharge Instructions|10543,10555|false|false|false|C0028900|Office Visits|office visit
Event|Event|Discharge Instructions|10550,10555|false|false|false|||visit
Finding|Social Behavior|Discharge Instructions|10550,10555|false|false|false|C0545082|Visit|visit
Event|Event|Discharge Instructions|10558,10562|false|false|false|||Make
Finding|Functional Concept|Discharge Instructions|10558,10562|false|false|false|C0947322;C1881534|Make - Instruction Imperative;Manufacturer Name|Make
Finding|Intellectual Product|Discharge Instructions|10558,10562|false|false|false|C0947322;C1881534|Make - Instruction Imperative;Manufacturer Name|Make
Event|Event|Discharge Instructions|10563,10567|false|false|false|||sure
Finding|Intellectual Product|Discharge Instructions|10563,10567|false|false|false|C4724437|SURE Test|sure
Event|Event|Discharge Instructions|10571,10579|false|false|false|||continue
Finding|Idea or Concept|Discharge Instructions|10571,10579|false|false|false|C0549178|Continuous|continue
Event|Event|Discharge Instructions|10583,10586|false|false|false|||use
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10592,10612|false|false|false|C0454512|Incentive spirometry|incentive spirometer
Finding|Finding|Discharge Instructions|10620,10627|true|false|false|C4534363|At home|at home
Finding|Idea or Concept|Discharge Instructions|10623,10627|true|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Discharge Instructions|10623,10627|true|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Discharge Instructions|10623,10627|true|false|false|C1553498|home health encounter|home
Event|Event|Discharge Instructions|10650,10660|true|false|false|||instructed
Procedure|Health Care Activity|Discharge Instructions|10673,10681|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|10682,10694|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|10682,10694|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|10682,10694|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

