 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|31,35
No|36,38
:|38,39
_|42,43
_|43,44
_|44,45
<EOL>|45,46
<EOL>|47,48
Admission|48,57
Date|58,62
:|62,63
_|65,66
_|66,67
_|67,68
Discharge|82,91
Date|92,96
:|96,97
_|100,101
_|101,102
_|102,103
<EOL>|103,104
<EOL>|105,106
Date|106,110
of|111,113
Birth|114,119
:|119,120
_|122,123
_|123,124
_|124,125
Sex|138,141
:|141,142
F|145,146
<EOL>|146,147
<EOL>|148,149
Service|149,156
:|156,157
MEDICINE|158,166
<EOL>|166,167
<EOL>|168,169
Sulfa|181,186
(|187,188
Sulfonamide|188,199
Antibiotics|200,211
)|211,212
/|213,214
Codeine|215,222
/|223,224
Bactrim|225,232
<EOL>|232,233
<EOL>|234,235
Attending|235,244
:|244,245
_|246,247
_|247,248
_|248,249
.|249,250
<EOL>|250,251
<EOL>|252,253
Weakness|271,279
,|279,280
nausea|281,287
/|287,288
vomiting|288,296
<EOL>|298,299
<EOL>|299,300
<EOL>|301,302
Major|302,307
Surgical|308,316
or|317,319
Invasive|320,328
Procedure|329,338
:|338,339
<EOL>|339,340
none|340,344
<EOL>|344,345
<EOL>|345,346
<EOL>|347,348
This|376,380
is|381,383
a|384,385
_|386,387
_|387,388
_|388,389
yo|390,392
f|393,394
with|395,399
h|400,401
/|401,402
o|402,403
recently|404,412
diagnosed|413,422
metastatic|423,433
cancer|434,440
<EOL>|441,442
of|442,444
unknown|445,452
prior|453,458
presenting|459,469
with|470,474
nausea|475,481
,|481,482
vomiting|483,491
,|491,492
and|493,496
fever|497,502
to|503,505
<EOL>|506,507
101|507,510
today|511,516
.|516,517
Patient|518,525
has|526,529
been|530,534
vomiting|535,543
over|544,548
the|549,552
past|553,557
6|558,559
-|560,561
8|562,563
weeks|564,569
,|569,570
<EOL>|571,572
since|572,577
before|578,584
she|585,588
was|589,592
diagnosed|593,602
with|603,607
metastatic|608,618
cancer|619,625
.|625,626
She|627,630
also|631,635
<EOL>|636,637
reports|637,644
pain|645,649
over|650,654
her|655,658
upper|659,664
abdomen|665,672
and|673,676
has|677,680
very|681,685
poor|686,690
PO|691,693
intake|694,700
.|700,701
<EOL>|702,703
She|703,706
has|707,710
been|711,715
feeling|716,723
progressively|724,737
weak|738,742
over|743,747
this|748,752
time|753,757
period|758,764
.|764,765
<EOL>|766,767
Her|767,770
vomiting|771,779
and|780,783
abdominal|784,793
pain|794,798
has|799,802
not|803,806
increased|807,816
from|817,821
the|822,825
past|826,830
<EOL>|831,832
weeks|832,837
,|837,838
but|839,842
she|843,846
just|847,851
feels|852,857
more|858,862
fatigued|863,871
.|871,872
She|873,876
has|877,880
a|881,882
chronic|883,890
<EOL>|891,892
non-productive|892,906
cough|907,912
as|913,915
well|916,920
.|920,921
No|922,924
URI|925,928
symptoms|929,937
,|937,938
no|939,941
urinary|942,949
<EOL>|950,951
complaints|951,961
.|961,962
She|963,966
has|967,970
been|971,975
constipated|976,987
,|987,988
which|989,994
improves|995,1003
when|1004,1008
she|1009,1012
<EOL>|1013,1014
stops|1014,1019
her|1020,1023
anti-emetics|1024,1036
.|1036,1037
Last|1038,1042
bowel|1043,1048
movement|1049,1057
was|1058,1061
yesterday|1062,1071
.|1071,1072
She|1073,1076
<EOL>|1077,1078
is|1078,1080
passing|1081,1088
gas|1089,1092
.|1092,1093
She|1094,1097
has|1098,1101
lower|1102,1107
extremity|1108,1117
edema|1118,1123
,|1123,1124
which|1125,1130
has|1131,1134
been|1135,1139
<EOL>|1140,1141
present|1141,1148
for|1149,1152
the|1153,1156
past|1157,1161
several|1162,1169
weeks|1170,1175
.|1175,1176
<EOL>|1178,1179
Of|1179,1181
note|1182,1186
,|1186,1187
she|1188,1191
was|1192,1195
supposed|1196,1204
to|1205,1207
have|1208,1212
one|1213,1216
of|1217,1219
her|1220,1223
liver|1224,1229
mets|1230,1234
biopsied|1235,1243
<EOL>|1244,1245
in|1245,1247
the|1248,1251
past|1252,1256
several|1257,1264
weeks|1265,1270
,|1270,1271
but|1272,1275
she|1276,1279
was|1280,1283
taking|1284,1290
ibuprofen|1291,1300
so|1301,1303
the|1304,1307
<EOL>|1308,1309
biopsy|1309,1315
had|1316,1319
to|1320,1322
be|1323,1325
postponed|1326,1335
.|1335,1336
<EOL>|1338,1339
<EOL>|1340,1341
In|1341,1343
the|1344,1347
ED|1348,1350
,|1350,1351
initial|1352,1359
VS|1360,1362
were|1363,1367
:|1367,1368
97.6|1369,1373
117|1374,1377
128|1378,1381
/|1381,1382
74|1382,1384
18|1385,1387
95|1388,1390
%|1390,1391
RA|1392,1394
.|1394,1395
Labs|1396,1400
were|1401,1405
<EOL>|1406,1407
significant|1407,1418
for|1419,1422
WBC|1423,1426
of|1427,1429
18.7|1430,1434
,|1434,1435
with|1436,1440
77|1441,1443
%|1443,1444
polys|1445,1450
.|1450,1451
UA|1452,1454
was|1455,1458
significant|1459,1470
<EOL>|1471,1472
for|1472,1475
ketones|1476,1483
.|1483,1484
Patient|1485,1492
received|1493,1501
zofran|1502,1508
,|1508,1509
NS|1510,1512
.|1512,1513
She|1514,1517
had|1518,1521
a|1522,1523
CXR|1524,1527
that|1528,1532
<EOL>|1533,1534
showed|1534,1540
new|1541,1544
left|1545,1549
sided|1550,1555
opacity|1556,1563
that|1564,1568
may|1569,1572
reflect|1573,1580
PNA|1581,1584
superimposed|1585,1597
<EOL>|1598,1599
on|1599,1601
metastatic|1602,1612
diseae|1613,1619
vs|1620,1622
.|1622,1623
lymphangiitic|1624,1637
spread|1638,1644
of|1645,1647
cancer|1648,1654
.|1654,1655
She|1656,1659
<EOL>|1660,1661
received|1661,1669
vanc|1670,1674
and|1675,1678
cefepime|1679,1687
for|1688,1691
pneumonia|1692,1701
.|1701,1702
Vitals|1703,1709
on|1710,1712
transfer|1713,1721
<EOL>|1722,1723
are|1723,1726
:|1726,1727
99.6|1728,1732
110|1733,1736
118|1737,1740
/|1740,1741
78|1741,1743
20|1744,1746
99|1747,1749
%|1749,1750
.|1750,1751
<EOL>|1753,1754
Currently|1754,1763
,|1763,1764
she|1765,1768
continues|1769,1778
to|1779,1781
feel|1782,1786
weak|1787,1791
and|1792,1795
nauseous|1796,1804
.|1804,1805
She|1806,1809
is|1810,1812
<EOL>|1813,1814
trying|1814,1820
to|1821,1823
take|1824,1828
her|1829,1832
pants|1833,1838
off|1839,1842
,|1842,1843
but|1844,1847
feels|1848,1853
too|1854,1857
weak|1858,1862
and|1863,1866
tired|1867,1872
to|1873,1875
do|1876,1878
<EOL>|1879,1880
so|1880,1882
.|1882,1883
<EOL>|1885,1886
REVIEW|1886,1892
OF|1893,1895
SYSTEMS|1896,1903
:|1903,1904
<EOL>|1906,1907
(|1907,1908
+|1908,1909
)|1909,1910
per|1911,1914
HPI|1915,1918
<EOL>|1920,1921
(|1921,1922
-|1922,1923
)|1923,1924
night|1925,1930
sweats|1931,1937
,|1937,1938
headache|1939,1947
,|1947,1948
vision|1949,1955
changes|1956,1963
,|1963,1964
rhinorrhea|1965,1975
,|1975,1976
<EOL>|1977,1978
congestion|1978,1988
,|1988,1989
sore|1990,1994
throat|1995,2001
,|2001,2002
BRBPR|2003,2008
,|2008,2009
melena|2010,2016
,|2016,2017
hematochezia|2018,2030
,|2030,2031
dysuria|2032,2039
,|2039,2040
<EOL>|2041,2042
hematuria|2042,2051
.|2051,2052
<EOL>|2054,2055
<EOL>|2056,2057
<EOL>|2057,2058
<EOL>|2059,2060
<EOL>|2081,2082
#|2088,2089
high|2090,2094
grade|2095,2100
SBO|2101,2104
_|2105,2106
_|2106,2107
_|2107,2108
s|2109,2110
/|2110,2111
p|2111,2112
exploratory|2113,2124
laparotomy|2125,2135
,|2135,2136
lysis|2137,2142
of|2143,2145
<EOL>|2146,2147
adhesions|2147,2156
,|2156,2157
and|2158,2161
small|2162,2167
bowel|2168,2173
resection|2174,2183
with|2184,2188
enteroenterostomy|2189,2206
<EOL>|2207,2208
#|2208,2209
carcinoid|2210,2219
<EOL>|2219,2220
#|2220,2221
hyperlipidemia|2222,2236
<EOL>|2236,2237
#|2237,2238
vitamin|2239,2246
B12|2247,2250
deficiency|2251,2261
<EOL>|2261,2262
#|2262,2263
cervical|2264,2272
DJD|2273,2276
<EOL>|2276,2277
#|2277,2278
osteoarthritis|2279,2293
<EOL>|2294,2295
<EOL>|2295,2296
PSH|2296,2299
:|2299,2300
<EOL>|2301,2302
s|2302,2303
/|2303,2304
p|2304,2305
R|2306,2307
lung|2308,2312
resection|2313,2322
in|2323,2325
_|2326,2327
_|2327,2328
_|2328,2329
at|2330,2332
_|2333,2334
_|2334,2335
_|2335,2336
<EOL>|2336,2337
s|2337,2338
/|2338,2339
p|2339,2340
hysterectomy|2341,2353
in|2354,2356
_|2357,2358
_|2358,2359
_|2359,2360
<EOL>|2360,2361
s|2361,2362
/|2362,2363
p|2363,2364
R|2365,2366
arm|2367,2370
surgery|2371,2378
<EOL>|2378,2379
<EOL>|2379,2380
<EOL>|2381,2382
:|2396,2397
<EOL>|2397,2398
_|2398,2399
_|2399,2400
_|2400,2401
<EOL>|2401,2402
:|2416,2417
<EOL>|2417,2418
Mother|2418,2424
-|2425,2426
_|2427,2428
_|2428,2429
_|2429,2430
cancer|2431,2437
d.|2438,2440
at|2441,2443
_|2444,2445
_|2445,2446
_|2446,2447
<EOL>|2449,2450
Youngest|2450,2458
of|2459,2461
_|2462,2463
_|2463,2464
_|2464,2465
-|2466,2467
not|2468,2471
in|2472,2474
touch|2475,2480
with|2481,2485
siblings|2486,2494
<EOL>|2496,2497
Father|2497,2503
-|2504,2505
_|2506,2507
_|2507,2508
_|2508,2509
d.|2510,2512
at|2513,2515
_|2516,2517
_|2517,2518
_|2518,2519
<EOL>|2521,2522
<EOL>|2522,2523
<EOL>|2524,2525
Admission|2540,2549
Physical|2550,2558
Exam|2559,2563
:|2563,2564
<EOL>|2565,2566
VS|2566,2568
:|2568,2569
98.6|2570,2574
,|2574,2575
130|2576,2579
/|2579,2580
80|2580,2582
,|2582,2583
111|2584,2587
,|2587,2588
24|2589,2591
,|2591,2592
98|2593,2595
%|2595,2596
on|2597,2599
RA|2600,2602
<EOL>|2604,2605
GENERAL|2605,2612
:|2612,2613
Obese|2614,2619
woman|2620,2625
,|2625,2626
appears|2627,2634
comfortable|2635,2646
,|2646,2647
in|2648,2650
no|2651,2653
acute|2654,2659
distress|2660,2668
<EOL>|2670,2671
<EOL>|2671,2672
HEENT|2672,2677
:|2677,2678
PERRLA|2679,2685
,|2685,2686
EOMI|2687,2691
,|2691,2692
sclerae|2693,2700
anicteric|2701,2710
,|2710,2711
slightly|2712,2720
dry|2721,2724
mucus|2725,2730
<EOL>|2731,2732
membranes|2732,2741
<EOL>|2743,2744
NECK|2744,2748
:|2748,2749
supple|2750,2756
,|2756,2757
obese|2758,2763
<EOL>|2765,2766
LUNGS|2766,2771
:|2771,2772
Distant|2773,2780
breath|2781,2787
sounds|2788,2794
,|2794,2795
decreased|2796,2805
on|2806,2808
the|2809,2812
right|2813,2818
,|2818,2819
few|2820,2823
<EOL>|2824,2825
crackles|2825,2833
b|2834,2835
/|2835,2836
l|2836,2837
<EOL>|2839,2840
HEART|2840,2845
:|2845,2846
RRR|2847,2850
,|2850,2851
no|2852,2854
MRG|2855,2858
,|2858,2859
nl|2860,2862
S1|2863,2865
-|2865,2866
S2|2866,2868
<EOL>|2870,2871
ABDOMEN|2871,2878
:|2878,2879
+|2880,2881
bowel|2882,2887
sounds|2888,2894
,|2894,2895
soft|2896,2900
,|2900,2901
epigastric|2902,2912
and|2913,2916
RUQ|2917,2920
tenderness|2921,2931
to|2932,2934
<EOL>|2935,2936
palpation|2936,2945
,|2945,2946
markedly|2947,2955
enlarged|2956,2964
liver|2965,2970
,|2970,2971
with|2972,2976
liver|2977,2982
edge|2983,2987
palpable|2988,2996
5|2997,2998
<EOL>|2999,3000
cm|3000,3002
below|3003,3008
rib|3009,3012
cage|3013,3017
.|3017,3018
No|3019,3021
rebound|3022,3029
/|3029,3030
guarding|3030,3038
.|3038,3039
<EOL>|3041,3042
EXTREMITIES|3042,3053
:|3053,3054
2|3055,3056
+|3056,3057
lower|3058,3063
extremity|3064,3073
edema|3074,3079
,|3079,3080
2|3081,3082
+|3082,3083
pulses|3084,3090
radial|3091,3097
and|3098,3101
dp|3102,3104
<EOL>|3106,3107
NEURO|3107,3112
:|3112,3113
awake|3114,3119
,|3119,3120
A|3121,3122
&|3122,3123
Ox3|3123,3126
,|3126,3127
CNs|3128,3131
II|3132,3134
-|3134,3135
XII|3135,3138
grossly|3139,3146
intact|3147,3153
,|3153,3154
muscle|3155,3161
strength|3162,3170
<EOL>|3171,3172
_|3172,3173
_|3173,3174
_|3174,3175
throughout|3176,3186
<EOL>|3188,3189
<EOL>|3189,3190
Discharge|3190,3199
Physical|3200,3208
Exam|3209,3213
:|3213,3214
<EOL>|3214,3215
Vitals|3215,3221
-|3221,3222
Tm|3224,3226
99.8|3227,3231
BP|3232,3234
125|3235,3238
/|3238,3239
76|3239,3241
HR|3242,3244
105|3245,3248
RR|3249,3251
20|3252,3254
99RA|3255,3259
<EOL>|3259,3260
General|3260,3267
-|3267,3268
Alert|3269,3274
,|3274,3275
oriented|3276,3284
,|3284,3285
no|3286,3288
acute|3289,3294
distress|3295,3303
,|3303,3304
obese|3305,3310
appearing|3311,3320
<EOL>|3321,3322
woman|3322,3327
<EOL>|3329,3330
HEENT|3330,3335
-|3335,3336
Sclera|3337,3343
anicteric|3344,3353
,|3353,3354
MMM|3355,3358
,|3358,3359
oropharynx|3360,3370
clear|3371,3376
<EOL>|3378,3379
Neck|3379,3383
-|3383,3384
supple|3385,3391
,|3391,3392
JVP|3393,3396
not|3397,3400
elevated|3401,3409
,|3409,3410
no|3411,3413
LAD|3414,3417
<EOL>|3419,3420
Lungs|3420,3425
-|3425,3426
Clear|3427,3432
to|3433,3435
auscultation|3436,3448
bilaterally|3449,3460
with|3461,3465
decreased|3466,3475
breath|3476,3482
<EOL>|3483,3484
sound|3484,3489
on|3490,3492
left|3493,3497
posterior|3498,3507
basilar|3508,3515
lung|3516,3520
field|3521,3526
,|3526,3527
no|3528,3530
wheezes|3531,3538
,|3538,3539
rales|3540,3545
,|3545,3546
<EOL>|3547,3548
ronchi|3548,3554
<EOL>|3556,3557
CV|3557,3559
-|3559,3560
Regular|3561,3568
rate|3569,3573
and|3574,3577
rhythm|3578,3584
,|3584,3585
normal|3586,3592
S1|3593,3595
+|3596,3597
S2|3598,3600
,|3600,3601
no|3602,3604
murmurs|3605,3612
,|3612,3613
rubs|3614,3618
,|3618,3619
<EOL>|3620,3621
gallops|3621,3628
<EOL>|3630,3631
Abdomen|3631,3638
-|3638,3639
soft|3640,3644
,|3644,3645
obese|3646,3651
,|3651,3652
diffusely|3653,3662
tender|3663,3669
,|3669,3670
non-distended|3671,3684
,|3684,3685
bowel|3686,3691
<EOL>|3692,3693
sounds|3693,3699
present|3700,3707
,|3707,3708
no|3709,3711
rebound|3712,3719
tenderness|3720,3730
or|3731,3733
guarding|3734,3742
,|3742,3743
no|3744,3746
<EOL>|3747,3748
organomegaly|3748,3760
<EOL>|3762,3763
GU|3763,3765
-|3765,3766
no|3767,3769
foley|3770,3775
<EOL>|3777,3778
Ext|3778,3781
-|3781,3782
warm|3783,3787
,|3787,3788
well|3789,3793
perfused|3794,3802
,|3802,3803
2|3804,3805
+|3805,3806
pulses|3807,3813
,|3813,3814
no|3815,3817
clubbing|3818,3826
,|3826,3827
cyanosis|3828,3836
,|3836,3837
2|3838,3839
+|3839,3840
<EOL>|3841,3842
pitting|3842,3849
edema|3850,3855
<EOL>|3857,3858
Neuro|3858,3863
-|3863,3864
CNs2|3865,3869
-|3869,3870
12|3870,3872
intact|3873,3879
,|3879,3880
motor|3881,3886
function|3887,3895
grossly|3896,3903
normal|3904,3910
<EOL>|3912,3913
Labs|3913,3917
:|3917,3918
Reviewed|3919,3927
,|3927,3928
please|3929,3935
see|3936,3939
below|3940,3945
.|3945,3946
<EOL>|3948,3949
<EOL>|3949,3950
<EOL>|3951,3952
Pertinent|3952,3961
Results|3962,3969
:|3969,3970
<EOL>|3970,3971
ADMIT|3971,3976
LABS|3977,3981
:|3981,3982
<EOL>|3982,3983
<EOL>|3983,3984
_|3984,3985
_|3985,3986
_|3986,3987
04|3988,3990
:|3990,3991
35PM|3991,3995
BLOOD|3996,4001
WBC|4002,4005
-|4005,4006
18|4006,4008
.|4008,4009
7|4009,4010
*|4010,4011
#|4011,4012
RBC|4013,4016
-|4016,4017
3|4017,4018
.|4018,4019
49|4019,4021
*|4021,4022
Hgb|4023,4026
-|4026,4027
9|4027,4028
.|4028,4029
2|4029,4030
*|4030,4031
Hct|4032,4035
-|4035,4036
31|4036,4038
.|4038,4039
2|4039,4040
*|4040,4041
<EOL>|4042,4043
MCV|4043,4046
-|4046,4047
90|4047,4049
MCH|4050,4053
-|4053,4054
26|4054,4056
.|4056,4057
5|4057,4058
*|4058,4059
MCHC|4060,4064
-|4064,4065
29|4065,4067
.|4067,4068
6|4068,4069
*|4069,4070
RDW|4071,4074
-|4074,4075
18|4075,4077
.|4077,4078
6|4078,4079
*|4079,4080
Plt|4081,4084
_|4085,4086
_|4086,4087
_|4087,4088
<EOL>|4088,4089
_|4089,4090
_|4090,4091
_|4091,4092
04|4093,4095
:|4095,4096
35PM|4096,4100
BLOOD|4101,4106
Neuts|4107,4112
-|4112,4113
77|4113,4115
.|4115,4116
4|4116,4117
*|4117,4118
Lymphs|4119,4125
-|4125,4126
14|4126,4128
.|4128,4129
9|4129,4130
*|4130,4131
Monos|4132,4137
-|4137,4138
6.8|4138,4141
<EOL>|4142,4143
Eos|4143,4146
-|4146,4147
0.5|4147,4150
Baso|4151,4155
-|4155,4156
0.4|4156,4159
<EOL>|4159,4160
_|4160,4161
_|4161,4162
_|4162,4163
04|4164,4166
:|4166,4167
35PM|4167,4171
BLOOD|4172,4177
Plt|4178,4181
_|4182,4183
_|4183,4184
_|4184,4185
<EOL>|4185,4186
_|4186,4187
_|4187,4188
_|4188,4189
04|4190,4192
:|4192,4193
35PM|4193,4197
BLOOD|4198,4203
Glucose|4204,4211
-|4211,4212
90|4212,4214
UreaN|4215,4220
-|4220,4221
8|4221,4222
Creat|4223,4228
-|4228,4229
0.5|4229,4232
Na|4233,4235
-|4235,4236
139|4236,4239
K|4240,4241
-|4241,4242
3.5|4242,4245
<EOL>|4246,4247
Cl|4247,4249
-|4249,4250
99|4250,4252
HCO3|4253,4257
-|4257,4258
29|4258,4260
AnGap|4261,4266
-|4266,4267
15|4267,4269
<EOL>|4269,4270
_|4270,4271
_|4271,4272
_|4272,4273
04|4274,4276
:|4276,4277
35PM|4277,4281
BLOOD|4282,4287
ALT|4288,4291
-|4291,4292
12|4292,4294
AST|4295,4298
-|4298,4299
48|4299,4301
*|4301,4302
AlkPhos|4303,4310
-|4310,4311
328|4311,4314
*|4314,4315
TotBili|4316,4323
-|4323,4324
0.9|4324,4327
<EOL>|4327,4328
_|4328,4329
_|4329,4330
_|4330,4331
07|4332,4334
:|4334,4335
45AM|4335,4339
BLOOD|4340,4345
Calcium|4346,4353
-|4353,4354
8.4|4354,4357
Phos|4358,4362
-|4362,4363
2|4363,4364
.|4364,4365
5|4365,4366
*|4366,4367
#|4367,4368
Mg|4369,4371
-|4371,4372
2.0|4372,4375
<EOL>|4375,4376
_|4376,4377
_|4377,4378
_|4378,4379
04|4380,4382
:|4382,4383
35PM|4383,4387
BLOOD|4388,4393
Albumin|4394,4401
-|4401,4402
2|4402,4403
.|4403,4404
8|4404,4405
*|4405,4406
<EOL>|4406,4407
_|4407,4408
_|4408,4409
_|4409,4410
06|4411,4413
:|4413,4414
42PM|4414,4418
BLOOD|4419,4424
Lactate|4425,4432
-|4432,4433
2.0|4433,4436
<EOL>|4436,4437
<EOL>|4437,4438
DISCHARGE|4438,4447
LABS|4449,4453
:|4453,4454
<EOL>|4454,4455
<EOL>|4455,4456
_|4456,4457
_|4457,4458
_|4458,4459
06|4460,4462
:|4462,4463
05AM|4463,4467
BLOOD|4468,4473
WBC|4474,4477
-|4477,4478
16|4478,4480
.|4480,4481
8|4481,4482
*|4482,4483
RBC|4484,4487
-|4487,4488
3|4488,4489
.|4489,4490
20|4490,4492
*|4492,4493
Hgb|4494,4497
-|4497,4498
8|4498,4499
.|4499,4500
3|4500,4501
*|4501,4502
Hct|4503,4506
-|4506,4507
28|4507,4509
.|4509,4510
7|4510,4511
*|4511,4512
<EOL>|4513,4514
MCV|4514,4517
-|4517,4518
90|4518,4520
MCH|4521,4524
-|4524,4525
25|4525,4527
.|4527,4528
9|4528,4529
*|4529,4530
MCHC|4531,4535
-|4535,4536
28|4536,4538
.|4538,4539
9|4539,4540
*|4540,4541
RDW|4542,4545
-|4545,4546
18|4546,4548
.|4548,4549
1|4549,4550
*|4550,4551
Plt|4552,4555
_|4556,4557
_|4557,4558
_|4558,4559
<EOL>|4559,4560
_|4560,4561
_|4561,4562
_|4562,4563
06|4564,4566
:|4566,4567
05AM|4567,4571
BLOOD|4572,4577
Glucose|4578,4585
-|4585,4586
87|4586,4588
UreaN|4589,4594
-|4594,4595
10|4595,4597
Creat|4598,4603
-|4603,4604
0.4|4604,4607
Na|4608,4610
-|4610,4611
136|4611,4614
<EOL>|4615,4616
K|4616,4617
-|4617,4618
3.7|4618,4621
Cl|4622,4624
-|4624,4625
99|4625,4627
HCO3|4628,4632
-|4632,4633
27|4633,4635
AnGap|4636,4641
-|4641,4642
14|4642,4644
<EOL>|4644,4645
_|4645,4646
_|4646,4647
_|4647,4648
06|4649,4651
:|4651,4652
05AM|4652,4656
BLOOD|4657,4662
ALT|4663,4666
-|4666,4667
11|4667,4669
AST|4670,4673
-|4673,4674
45|4674,4676
*|4676,4677
LD|4678,4680
(|4680,4681
LDH|4681,4684
)|4684,4685
-|4685,4686
517|4686,4689
*|4689,4690
AlkPhos|4691,4698
-|4698,4699
282|4699,4702
*|4702,4703
<EOL>|4704,4705
TotBili|4705,4712
-|4712,4713
0.8|4713,4716
<EOL>|4716,4717
_|4717,4718
_|4718,4719
_|4719,4720
06|4721,4723
:|4723,4724
05AM|4724,4728
BLOOD|4729,4734
Calcium|4735,4742
-|4742,4743
8.4|4743,4746
Phos|4747,4751
-|4751,4752
2.7|4752,4755
Mg|4756,4758
-|4758,4759
2.2|4759,4762
<EOL>|4762,4763
<EOL>|4763,4764
IMAGING|4764,4771
:|4771,4772
_|4773,4774
_|4774,4775
_|4775,4776
<EOL>|4776,4777
Final|4777,4782
Report|4783,4789
<EOL>|4790,4791
HISTORY|4791,4798
:|4798,4799
New|4801,4804
diagnosis|4805,4814
of|4815,4817
metastatic|4818,4828
cancer|4829,4835
with|4836,4840
unknown|4841,4848
<EOL>|4849,4850
primary|4850,4857
.|4857,4858
Assess|4860,4866
for|4867,4870
extent|4871,4877
of|4878,4880
lesions|4881,4888
.|4888,4889
<EOL>|4892,4893
COMPARISON|4893,4903
:|4903,4904
CT|4906,4908
abdomen|4909,4916
and|4917,4920
pelvis|4921,4927
dated|4928,4933
_|4934,4935
_|4935,4936
_|4936,4937
.|4937,4938
<EOL>|4940,4941
TECHNIQUE|4941,4950
:|4950,4951
Multidetector|4953,4966
CT|4967,4969
of|4970,4972
the|4973,4976
torso|4977,4982
was|4983,4986
performed|4987,4996
with|4997,5001
<EOL>|5002,5003
intravenous|5003,5014
and|5015,5018
oral|5019,5023
contrast|5024,5032
.|5032,5033
Coronal|5035,5042
and|5043,5046
sagittal|5047,5055
<EOL>|5056,5057
reformations|5057,5069
were|5070,5074
provided|5075,5083
.|5083,5084
Images|5086,5092
are|5093,5096
substantially|5097,5110
degraded|5111,5119
<EOL>|5120,5121
due|5121,5124
to|5125,5127
the|5128,5131
patient|5132,5139
's|5139,5141
body|5142,5146
habitus|5147,5154
.|5154,5155
<EOL>|5158,5159
:|5167,5168
<EOL>|5169,5170
CHEST|5170,5175
:|5175,5176
<EOL>|5178,5179
There|5179,5184
are|5185,5188
innumerable|5189,5200
pulmonary|5201,5210
nodules|5211,5218
,|5218,5219
which|5220,5225
have|5226,5230
an|5231,5233
upper|5234,5239
<EOL>|5240,5241
lobe|5241,5245
<EOL>|5246,5247
predilection|5247,5259
,|5259,5260
particularly|5261,5273
in|5274,5276
the|5277,5280
left|5281,5285
upper|5286,5291
lobe|5292,5296
.|5296,5297
The|5299,5302
largest|5303,5310
<EOL>|5311,5312
nodule|5312,5318
<EOL>|5319,5320
measures|5320,5328
6|5329,5330
mm|5331,5333
in|5334,5336
diameter|5337,5345
(|5346,5347
sequence|5347,5355
3|5356,5357
image|5358,5363
8|5364,5365
)|5365,5366
.|5366,5367
Calcification|5369,5382
<EOL>|5383,5384
is|5384,5386
noted|5387,5392
within|5393,5399
the|5401,5404
right|5405,5410
pleural|5411,5418
cavity|5419,5425
(|5426,5427
sequence|5427,5435
3|5436,5437
image|5438,5443
24|5444,5446
)|5446,5447
,|5447,5448
<EOL>|5449,5450
which|5450,5455
is|5456,5458
likely|5459,5465
related|5466,5473
to|5474,5476
the|5477,5480
patient|5481,5488
's|5488,5490
history|5491,5498
of|5499,5501
previous|5502,5510
<EOL>|5511,5512
right|5512,5517
lung|5518,5522
surgery|5523,5530
.|5530,5531
No|5533,5535
pleural|5536,5543
effusion|5544,5552
.|5552,5553
No|5555,5557
pneumothorax|5558,5570
.|5570,5571
<EOL>|5573,5574
No|5574,5576
significant|5577,5588
mediastinal|5589,5600
,|5600,5601
axillary|5602,5610
or|5611,5613
hilar|5614,5619
adenopathy|5620,5630
.|5630,5631
<EOL>|5633,5634
Cardiac|5634,5641
size|5642,5646
is|5647,5649
<EOL>|5650,5651
normal|5651,5657
.|5657,5658
No|5660,5662
pericardial|5663,5674
effusion|5675,5683
.|5683,5684
<EOL>|5686,5687
ABDOMEN|5687,5694
:|5694,5695
<EOL>|5697,5698
The|5698,5701
liver|5702,5707
is|5708,5710
enlarged|5711,5719
and|5720,5723
there|5724,5729
are|5730,5733
innumerable|5734,5745
_|5746,5747
_|5747,5748
_|5748,5749
density|5750,5757
<EOL>|5758,5759
lesions|5759,5766
throughout|5767,5777
both|5778,5782
lobes|5783,5788
of|5789,5791
the|5792,5795
liver|5796,5801
which|5802,5807
are|5808,5811
replacing|5812,5821
<EOL>|5822,5823
the|5823,5826
vast|5827,5831
majority|5832,5840
of|5841,5843
the|5844,5847
hepatic|5848,5855
parenchyma|5856,5866
.|5866,5867
The|5869,5872
portal|5873,5879
vein|5880,5884
is|5885,5887
<EOL>|5888,5889
patent|5889,5895
.|5895,5896
No|5898,5900
intra|5901,5906
or|5907,5909
extrahepatic|5910,5922
duct|5923,5927
dilatation|5928,5938
.|5938,5939
The|5941,5944
<EOL>|5945,5946
gallbladder|5946,5957
is|5958,5960
unremarkable|5961,5973
.|5973,5974
There|5976,5981
is|5982,5984
a|5985,5986
small|5987,5992
amount|5993,5999
of|6000,6002
ascites|6003,6010
<EOL>|6011,6012
adjacent|6012,6020
to|6021,6023
the|6024,6027
right|6028,6033
lobe|6034,6038
of|6039,6041
the|6042,6045
liver|6046,6051
.|6051,6052
<EOL>|6055,6056
<EOL>|6058,6059
The|6059,6062
right|6063,6068
kidney|6069,6075
is|6076,6078
mildly|6079,6085
compressed|6086,6096
anteriorly|6097,6107
due|6108,6111
to|6112,6114
the|6115,6118
<EOL>|6119,6120
enlarged|6120,6128
liver|6129,6134
.|6134,6135
There|6136,6141
is|6142,6144
a|6145,6146
subcentimeter|6147,6160
_|6161,6162
_|6162,6163
_|6163,6164
density|6165,6172
lesion|6173,6179
in|6180,6182
<EOL>|6183,6184
the|6184,6187
upper|6188,6193
pole|6194,6198
of|6199,6201
the|6202,6205
right|6206,6211
kidney|6212,6218
,|6218,6219
likely|6220,6226
representing|6227,6239
a|6240,6241
<EOL>|6242,6243
subcentimeter|6243,6256
cyst|6257,6261
(|6262,6263
sequence|6263,6271
5|6272,6273
image|6274,6279
31|6280,6282
)|6282,6283
.|6283,6284
The|6286,6289
right|6290,6295
kidney|6296,6302
is|6303,6305
<EOL>|6306,6307
otherwise|6307,6316
unremarkable|6317,6329
.|6329,6330
The|6332,6335
left|6336,6340
kidney|6341,6347
is|6348,6350
within|6351,6357
normal|6358,6364
<EOL>|6365,6366
limits|6366,6372
.|6372,6373
The|6375,6378
adrenals|6379,6387
and|6388,6391
spleen|6392,6398
are|6399,6402
unremarkable|6403,6415
.|6415,6416
The|6418,6421
pancreas|6422,6430
<EOL>|6431,6432
is|6432,6434
within|6435,6441
normal|6442,6448
limits|6449,6455
.|6455,6456
The|6458,6461
small|6462,6467
and|6468,6471
large|6472,6477
bowel|6478,6483
are|6484,6487
<EOL>|6488,6489
unremarkable|6489,6501
.|6501,6502
No|6504,6506
retroperitoneal|6507,6522
or|6523,6525
mesenteric|6526,6536
adenopathy|6537,6547
.|6547,6548
<EOL>|6550,6551
<EOL>|6553,6554
PELVIS|6554,6560
:|6560,6561
<EOL>|6563,6564
The|6564,6567
images|6568,6574
of|6575,6577
the|6578,6581
pelvis|6582,6588
are|6589,6592
substantially|6593,6606
degraded|6607,6615
secondary|6616,6625
to|6626,6628
<EOL>|6629,6630
the|6630,6633
patient|6634,6641
's|6641,6643
body|6644,6648
habitus|6649,6656
.|6656,6657
No|6659,6661
pelvic|6662,6668
masses|6669,6675
are|6676,6679
identified|6680,6690
.|6690,6691
<EOL>|6693,6694
The|6694,6697
bladder|6698,6705
is|6706,6708
unremarkable|6709,6721
.|6721,6722
The|6724,6727
patient|6728,6735
is|6736,6738
status|6739,6745
post|6746,6750
<EOL>|6751,6752
supracervical|6752,6765
hysterectomy|6766,6778
.|6778,6779
No|6781,6783
pelvic|6784,6790
adenopathy|6791,6801
.|6801,6802
No|6803,6805
free|6806,6810
fluid|6811,6816
<EOL>|6817,6818
within|6818,6824
the|6825,6828
pelvis|6829,6835
.|6835,6836
<EOL>|6838,6839
<EOL>|6841,6842
OSSEOUS|6842,6849
STRUCTURES|6850,6860
:|6860,6861
<EOL>|6863,6864
Bilateral|6864,6873
symmetrical|6874,6885
sclerosis|6886,6895
is|6896,6898
identified|6899,6909
on|6910,6912
the|6913,6916
iliac|6917,6922
side|6923,6927
<EOL>|6928,6929
of|6929,6931
the|6932,6935
<EOL>|6936,6937
sacroiliac|6937,6947
joints|6948,6954
,|6954,6955
consistent|6956,6966
with|6967,6971
osteitis|6972,6980
condensans|6981,6991
ilii|6992,6996
.|6996,6997
<EOL>|6999,7000
There|7000,7005
is|7006,7008
severe|7009,7015
degenerative|7016,7028
change|7029,7035
within|7036,7042
the|7043,7046
right|7047,7052
hip|7053,7056
joint|7057,7062
<EOL>|7063,7064
with|7064,7068
joint|7069,7074
space|7075,7080
loss|7081,7085
and|7086,7089
osteophyte|7090,7100
formation|7101,7110
.|7110,7111
No|7113,7115
destructive|7116,7127
<EOL>|7128,7129
osseous|7129,7136
lesions|7137,7144
.|7144,7145
<EOL>|7148,7149
<EOL>|7151,7152
Multiple|7165,7173
pulmonary|7174,7183
and|7184,7187
hepatic|7188,7195
metastases|7196,7206
.|7206,7207
No|7209,7211
separate|7212,7220
primary|7221,7228
<EOL>|7229,7230
lesion|7230,7236
<EOL>|7237,7238
identified|7238,7248
.|7248,7249
<EOL>|7252,7253
<EOL>|7253,7254
<EOL>|7255,7256
_|7279,7280
_|7280,7281
_|7281,7282
yo|7283,7285
f|7286,7287
with|7288,7292
h|7293,7294
/|7294,7295
o|7295,7296
recently|7297,7305
diagnosed|7306,7315
metastatic|7316,7326
cancer|7327,7333
of|7334,7336
unknown|7337,7344
<EOL>|7345,7346
primary|7346,7353
presenting|7354,7364
with|7365,7369
nausea|7370,7376
,|7376,7377
vomiting|7378,7386
,|7386,7387
and|7388,7391
fever|7392,7397
to|7398,7400
101|7401,7404
on|7405,7407
<EOL>|7408,7409
day|7409,7412
of|7413,7415
admission|7416,7425
.|7425,7426
<EOL>|7428,7429
.|7429,7430
<EOL>|7430,7431
#|7431,7432
Fever|7433,7438
/|7438,7439
leukocytosis|7439,7451
:|7451,7452
Patient|7453,7460
presented|7461,7470
with|7471,7475
fever|7476,7481
and|7482,7485
<EOL>|7486,7487
leukocytosis|7487,7499
,|7499,7500
which|7501,7506
was|7507,7510
initially|7511,7520
concerning|7521,7531
for|7532,7535
post|7536,7540
<EOL>|7541,7542
obstructive|7542,7553
PNA|7554,7557
.|7557,7558
Patient|7559,7566
was|7567,7570
treated|7571,7578
with|7579,7583
vanc|7584,7588
-|7588,7589
cefepime|7589,7597
-|7597,7598
azithro|7598,7605
<EOL>|7606,7607
for|7607,7610
a|7611,7612
day|7613,7616
and|7617,7620
a|7621,7622
half|7623,7627
,|7627,7628
however|7629,7636
CT|7637,7639
torso|7640,7645
was|7646,7649
concerning|7650,7660
for|7661,7664
<EOL>|7665,7666
ongoing|7666,7673
malignancy|7674,7684
without|7685,7692
evidence|7693,7701
of|7702,7704
primary|7705,7712
tumor|7713,7718
.|7718,7719
There|7720,7725
was|7726,7729
<EOL>|7730,7731
no|7731,7733
concern|7734,7741
for|7742,7745
a|7746,7747
pneumonia|7748,7757
.|7757,7758
Consequently|7759,7771
,|7771,7772
abx|7773,7776
were|7777,7781
stopped|7782,7789
on|7790,7792
<EOL>|7793,7794
_|7794,7795
_|7795,7796
_|7796,7797
.|7797,7798
Patient|7799,7806
felt|7807,7811
weak|7812,7816
and|7817,7820
unable|7821,7827
to|7828,7830
go|7831,7833
home|7834,7838
,|7838,7839
as|7840,7842
she|7843,7846
lives|7847,7852
<EOL>|7853,7854
alone|7854,7859
and|7860,7863
so|7864,7866
was|7867,7870
screened|7871,7879
by|7880,7882
physical|7883,7891
therapy|7892,7899
and|7900,7903
discharged|7904,7914
to|7915,7917
<EOL>|7918,7919
rehab|7919,7924
facility|7925,7933
.|7933,7934
<EOL>|7935,7936
.|7936,7937
<EOL>|7937,7938
#|7938,7939
Failure|7940,7947
to|7948,7950
thrive|7951,7957
:|7957,7958
Patient|7959,7966
presents|7967,7975
with|7976,7980
6|7981,7982
weeks|7983,7988
of|7989,7991
nausea|7992,7998
,|7998,7999
<EOL>|8000,8001
vomiting|8001,8009
and|8010,8013
poor|8014,8018
PO|8019,8021
intake|8022,8028
likely|8029,8035
from|8036,8040
her|8041,8044
enlarged|8045,8053
liver|8054,8059
.|8059,8060
She|8061,8064
<EOL>|8065,8066
continues|8066,8075
to|8076,8078
have|8079,8083
bowel|8084,8089
movements|8090,8099
and|8100,8103
pass|8104,8108
gas|8109,8112
.|8112,8113
Patient|8114,8121
now|8122,8125
with|8126,8130
<EOL>|8131,8132
albumin|8132,8139
of|8140,8142
2.8|8143,8146
,|8146,8147
ketones|8148,8155
in|8156,8158
her|8159,8162
urine|8163,8168
,|8168,8169
weight|8170,8176
loss|8177,8181
and|8182,8185
new|8186,8189
<EOL>|8190,8191
peripheral|8191,8201
edema|8202,8207
,|8207,8208
concerning|8209,8219
for|8220,8223
poor|8224,8228
nutrition|8229,8238
/|8238,8239
starvation|8239,8249
<EOL>|8250,8251
ketosis|8251,8258
.|8258,8259
Nutrition|8260,8269
consult|8270,8277
followed|8278,8286
the|8287,8290
patient|8291,8298
throughout|8299,8309
her|8310,8313
<EOL>|8314,8315
hospital|8315,8323
stay|8324,8328
and|8329,8332
recommended|8333,8344
_|8345,8346
_|8346,8347
_|8347,8348
fat|8349,8352
Carnation|8353,8362
Instant|8363,8370
<EOL>|8371,8372
Breakfast|8372,8381
with|8382,8386
Beneprotein|8387,8398
.|8398,8399
<EOL>|8399,8400
.|8400,8401
<EOL>|8401,8402
#|8402,8403
Chronic|8404,8411
back|8412,8416
pain|8417,8421
:|8421,8422
Patient|8424,8431
was|8432,8435
continued|8436,8445
on|8446,8448
her|8449,8452
home|8453,8457
<EOL>|8458,8459
gabapentin|8459,8469
.|8469,8470
<EOL>|8471,8472
.|8472,8473
<EOL>|8473,8474
#|8474,8475
Depression|8476,8486
:|8486,8487
Patient|8489,8496
was|8497,8500
continued|8501,8510
on|8511,8513
home|8514,8518
bupropion|8519,8528
,|8528,8529
<EOL>|8530,8531
sertraline|8531,8541
<EOL>|8543,8544
.|8544,8545
<EOL>|8545,8546
#|8546,8547
HCTZ|8548,8552
:|8552,8553
Patient|8554,8561
's|8561,8563
hctz|8564,8568
was|8569,8572
discontinued|8573,8585
during|8586,8592
her|8593,8596
<EOL>|8597,8598
hospitalization|8598,8613
due|8614,8617
to|8618,8620
poor|8621,8625
PO|8626,8628
intake|8629,8635
and|8636,8639
concern|8640,8647
for|8648,8651
<EOL>|8652,8653
dehydration|8653,8664
.|8664,8665
Blood|8666,8671
pressures|8672,8681
were|8682,8686
well|8687,8691
-|8691,8692
controlled|8692,8702
such|8703,8707
that|8708,8712
HCTZ|8713,8717
<EOL>|8718,8719
was|8719,8722
not|8723,8726
deemed|8727,8733
necessary|8734,8743
.|8743,8744
This|8745,8749
issue|8750,8755
should|8756,8762
be|8763,8765
readdressed|8766,8777
by|8778,8780
<EOL>|8781,8782
PCP|8782,8785
.|8785,8786
<EOL>|8786,8787
.|8787,8788
<EOL>|8788,8789
#|8789,8790
Hyperlipidemia|8791,8805
:|8805,8806
Given|8807,8812
patient|8813,8820
's|8820,8822
metastatic|8823,8833
process|8834,8841
,|8841,8842
statin|8843,8849
was|8850,8853
<EOL>|8854,8855
discontinued|8855,8867
during|8868,8874
hospitalization|8875,8890
to|8891,8893
simplify|8894,8902
her|8903,8906
medical|8907,8914
<EOL>|8915,8916
regimen|8916,8923
.|8923,8924
<EOL>|8926,8927
.|8927,8928
<EOL>|8928,8929
#|8929,8930
Insomnia|8931,8939
:|8939,8940
Continued|8941,8950
home|8951,8955
trazodone|8956,8965
<EOL>|8967,8968
.|8968,8969
<EOL>|8969,8970
TRANSITION|8970,8980
ISSUES|8981,8987
<EOL>|8987,8988
#|8988,8989
CODE|8990,8994
:|8994,8995
FULL|8996,9000
(|9001,9002
Confirmed|9002,9011
)|9011,9012
<EOL>|9014,9015
#|9015,9016
CONTACT|9017,9024
:|9024,9025
_|9026,9027
_|9027,9028
_|9028,9029
(|9030,9031
friend|9031,9037
)|9037,9038
_|9039,9040
_|9040,9041
_|9041,9042
<EOL>|9044,9045
#|9045,9046
HCTZ|9047,9051
discontinued|9052,9064
on|9065,9067
admission|9068,9077
-|9077,9078
consider|9079,9087
restarting|9088,9098
if|9099,9101
<EOL>|9102,9103
considered|9103,9113
medically|9114,9123
necessary|9124,9133
by|9134,9136
PCP|9137,9140
<EOL>|9141,9142
#|9142,9143
_|9144,9145
_|9145,9146
_|9146,9147
fat|9148,9151
Carnation|9152,9161
Instant|9162,9169
Breakfast|9170,9179
with|9180,9184
Beneprotein|9185,9196
with|9197,9201
<EOL>|9202,9203
meals|9203,9208
<EOL>|9208,9209
#|9209,9210
Follow|9211,9217
up|9218,9220
with|9221,9225
oncology|9226,9234
for|9235,9238
further|9239,9246
diagnosis|9247,9256
and|9257,9260
management|9261,9271
<EOL>|9272,9273
of|9273,9275
malignancy|9276,9286
<EOL>|9286,9287
<EOL>|9288,9289
Medications|9289,9300
on|9301,9303
Admission|9304,9313
:|9313,9314
<EOL>|9314,9315
The|9315,9318
Preadmission|9319,9331
Medication|9332,9342
list|9343,9347
is|9348,9350
accurate|9351,9359
and|9360,9363
complete|9364,9372
.|9372,9373
<EOL>|9373,9374
1.|9374,9376
Albuterol|9377,9386
Inhaler|9387,9394
_|9395,9396
_|9396,9397
_|9397,9398
PUFF|9399,9403
IH|9404,9406
Q6H|9407,9410
:|9410,9411
PRN|9411,9414
SOB|9415,9418
<EOL>|9419,9420
2.|9420,9422
BuPROPion|9423,9432
150|9433,9436
mg|9437,9439
PO|9440,9442
DAILY|9443,9448
<EOL>|9449,9450
3.|9450,9452
Gabapentin|9453,9463
300|9464,9467
mg|9468,9470
PO|9471,9473
HS|9474,9476
<EOL>|9477,9478
4.|9478,9480
Sertraline|9481,9491
200|9492,9495
mg|9496,9498
PO|9499,9501
DAILY|9502,9507
<EOL>|9508,9509
5.|9509,9511
Simvastatin|9512,9523
40|9524,9526
mg|9527,9529
PO|9530,9532
DAILY|9533,9538
<EOL>|9539,9540
6.|9540,9542
traZODONE|9543,9552
100|9553,9556
mg|9557,9559
PO|9560,9562
HS|9563,9565
:|9565,9566
PRN|9566,9569
sleep|9570,9575
<EOL>|9576,9577
7.|9577,9579
Ibuprofen|9580,9589
800|9590,9593
mg|9594,9596
PO|9597,9599
Q12H|9600,9604
:|9604,9605
PRN|9605,9608
pain|9609,9613
<EOL>|9614,9615
8.|9615,9617
Hydrochlorothiazide|9618,9637
12.5|9638,9642
mg|9643,9645
PO|9646,9648
DAILY|9649,9654
<EOL>|9655,9656
9.|9656,9658
Ondansetron|9659,9670
4|9671,9672
mg|9673,9675
PO|9676,9678
Q8H|9679,9682
:|9682,9683
PRN|9683,9686
nausea|9687,9693
<EOL>|9694,9695
<EOL>|9695,9696
<EOL>|9697,9698
Discharge|9698,9707
Medications|9708,9719
:|9719,9720
<EOL>|9720,9721
1.|9721,9723
Albuterol|9724,9733
Inhaler|9734,9741
_|9742,9743
_|9743,9744
_|9744,9745
PUFF|9746,9750
IH|9751,9753
Q6H|9754,9757
:|9757,9758
PRN|9758,9761
SOB|9762,9765
<EOL>|9766,9767
2.|9767,9769
BuPROPion|9770,9779
150|9780,9783
mg|9784,9786
PO|9787,9789
DAILY|9790,9795
<EOL>|9796,9797
3.|9797,9799
Gabapentin|9800,9810
300|9811,9814
mg|9815,9817
PO|9818,9820
HS|9821,9823
<EOL>|9824,9825
4.|9825,9827
Sertraline|9828,9838
200|9839,9842
mg|9843,9845
PO|9846,9848
DAILY|9849,9854
<EOL>|9855,9856
5.|9856,9858
traZODONE|9859,9868
100|9869,9872
mg|9873,9875
PO|9876,9878
HS|9879,9881
:|9881,9882
PRN|9882,9885
sleep|9886,9891
<EOL>|9892,9893
6.|9893,9895
Ondansetron|9896,9907
4|9908,9909
mg|9910,9912
PO|9913,9915
Q8H|9916,9919
:|9919,9920
PRN|9920,9923
nausea|9924,9930
<EOL>|9931,9932
7.|9932,9934
Bisacodyl|9935,9944
10|9945,9947
mg|9948,9950
PO|9951,9953
/|9953,9954
PR|9954,9956
DAILY|9957,9962
:|9962,9963
PRN|9963,9966
constipation|9967,9979
<EOL>|9980,9981
8.|9981,9983
OxycoDONE|9984,9993
(|9994,9995
Immediate|9995,10004
Release|10005,10012
)|10012,10013
5|10015,10016
mg|10017,10019
PO|10020,10022
Q6H|10023,10026
:|10026,10027
PRN|10027,10030
pain|10031,10035
<EOL>|10036,10037
please|10037,10043
hold|10044,10048
for|10049,10052
sedation|10053,10061
,|10061,10062
RR|10063,10065
<|10065,10066
10|10066,10068
<EOL>|10069,10070
RX|10070,10072
*|10073,10074
oxycodone|10074,10083
5|10084,10085
mg|10086,10088
1|10089,10090
tablet|10091,10097
(|10097,10098
s|10098,10099
)|10099,10100
by|10101,10103
mouth|10104,10109
every|10110,10115
6|10116,10117
hours|10118,10123
Disp|10124,10128
#|10129,10130
*|10130,10131
30|10131,10133
<EOL>|10134,10135
Tablet|10135,10141
Refills|10142,10149
:|10149,10150
*|10150,10151
0|10151,10152
<EOL>|10152,10153
9.|10153,10155
Enoxaparin|10156,10166
Sodium|10167,10173
40|10174,10176
mg|10177,10179
SC|10180,10182
DAILY|10183,10188
<EOL>|10189,10190
<EOL>|10190,10191
<EOL>|10192,10193
Discharge|10193,10202
Disposition|10203,10214
:|10214,10215
<EOL>|10215,10216
Extended|10216,10224
Care|10225,10229
<EOL>|10229,10230
<EOL>|10231,10232
Facility|10232,10240
:|10240,10241
<EOL>|10241,10242
_|10242,10243
_|10243,10244
_|10244,10245
<EOL>|10245,10246
<EOL>|10247,10248
Discharge|10248,10257
Diagnosis|10258,10267
:|10267,10268
<EOL>|10268,10269
Metastatic|10269,10279
disease|10280,10287
of|10288,10290
unknown|10291,10298
primary|10299,10306
:|10306,10307
Weakness|10308,10316
and|10317,10320
nausea|10321,10327
<EOL>|10328,10329
likely|10329,10335
from|10336,10340
tumor|10341,10346
burden|10347,10353
<EOL>|10353,10354
<EOL>|10354,10355
<EOL>|10356,10357
Mental|10378,10384
Status|10385,10391
:|10391,10392
Clear|10393,10398
and|10399,10402
coherent|10403,10411
.|10411,10412
<EOL>|10412,10413
Level|10413,10418
of|10419,10421
Consciousness|10422,10435
:|10435,10436
Alert|10437,10442
and|10443,10446
interactive|10447,10458
.|10458,10459
<EOL>|10459,10460
Activity|10460,10468
Status|10469,10475
:|10475,10476
Ambulatory|10477,10487
-|10488,10489
Independent|10490,10501
.|10501,10502
<EOL>|10502,10503
<EOL>|10503,10504
<EOL>|10505,10506
Dear|10530,10534
Ms.|10535,10538
_|10539,10540
_|10540,10541
_|10541,10542
,|10542,10543
<EOL>|10543,10544
<EOL>|10544,10545
You|10545,10548
were|10549,10553
admitted|10554,10562
to|10563,10565
_|10566,10567
_|10567,10568
_|10568,10569
for|10570,10573
evaluation|10574,10584
of|10585,10587
several|10588,10595
weeks|10596,10601
of|10602,10604
<EOL>|10605,10606
weakness|10606,10614
and|10615,10618
nausea|10619,10625
.|10625,10626
You|10627,10630
had|10631,10634
some|10635,10639
markers|10640,10647
of|10648,10650
infection|10651,10660
,|10660,10661
so|10662,10664
you|10665,10668
<EOL>|10669,10670
were|10670,10674
initially|10675,10684
given|10685,10690
antibiotics|10691,10702
.|10702,10703
However|10704,10711
,|10711,10712
a|10713,10714
scan|10715,10719
of|10720,10722
your|10723,10727
torso|10728,10733
<EOL>|10734,10735
showed|10735,10741
metastatic|10742,10752
disease|10753,10760
from|10761,10765
a|10766,10767
cancer|10768,10774
of|10775,10777
unknown|10778,10785
origin|10786,10792
in|10793,10795
<EOL>|10796,10797
your|10797,10801
liver|10802,10807
and|10808,10811
lungs|10812,10817
.|10817,10818
Your|10819,10823
weakness|10824,10832
and|10833,10836
nausea|10837,10843
are|10844,10847
most|10848,10852
likely|10853,10859
<EOL>|10860,10861
due|10861,10864
to|10865,10867
your|10868,10872
enlarged|10873,10881
liver|10882,10887
.|10887,10888
<EOL>|10889,10890
<EOL>|10890,10891
You|10891,10894
are|10895,10898
scheduled|10899,10908
to|10909,10911
see|10912,10915
your|10916,10920
oncologist|10921,10931
this|10932,10936
week|10937,10941
,|10941,10942
so|10943,10945
please|10946,10952
<EOL>|10953,10954
follow|10954,10960
-|10960,10961
up|10961,10963
with|10964,10968
them|10969,10973
so|10974,10976
that|10977,10981
they|10982,10986
may|10987,10990
proceed|10991,10998
with|10999,11003
the|11004,11007
further|11008,11015
<EOL>|11016,11017
diagnosis|11017,11026
and|11027,11030
treatment|11031,11040
of|11041,11043
your|11044,11048
malignancy|11049,11059
.|11059,11060
<EOL>|11060,11061
<EOL>|11061,11062
You|11062,11065
are|11066,11069
being|11070,11075
discharged|11076,11086
to|11087,11089
a|11090,11091
rehabilitation|11092,11106
facility|11107,11115
to|11116,11118
help|11119,11123
<EOL>|11124,11125
you|11125,11128
regain|11129,11135
some|11136,11140
strength|11141,11149
before|11150,11156
going|11157,11162
home|11163,11167
.|11167,11168
Your|11169,11173
anticipated|11174,11185
<EOL>|11186,11187
length|11187,11193
of|11194,11196
stay|11197,11201
is|11202,11204
LESS|11205,11209
THAN|11210,11214
30|11215,11217
DAYS|11218,11222
.|11222,11223
<EOL>|11224,11225
<EOL>|11225,11226
Please|11226,11232
see|11233,11236
the|11237,11240
attached|11241,11249
sheet|11250,11255
for|11256,11259
your|11260,11264
updated|11265,11272
medication|11273,11283
list|11284,11288
.|11288,11289
<EOL>|11290,11291
<EOL>|11291,11292
It|11292,11294
was|11295,11298
a|11299,11300
pleasure|11301,11309
taking|11310,11316
care|11317,11321
of|11322,11324
you|11325,11328
in|11329,11331
the|11332,11335
hospital|11336,11344
.|11344,11345
We|11346,11348
wish|11349,11353
<EOL>|11354,11355
you|11355,11358
all|11359,11362
the|11363,11366
best|11367,11371
.|11371,11372
<EOL>|11372,11373
<EOL>|11374,11375
Followup|11375,11383
Instructions|11384,11396
:|11396,11397
<EOL>|11397,11398
_|11398,11399
_|11399,11400
_|11400,11401
<EOL>|11401,11402

