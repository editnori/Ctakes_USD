CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Orthopedics|Title|false|false||ORTHOPAEDICSnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|sulfa|Drug|false|false||Sulfanull|Sulfonamide Anti-Infective Agents|Drug|false|false||Sulfonamide
null|Sulfonamide Anti-Infective Agents|Drug|false|false||Sulfonamide
null|Sulfonamides|Drug|false|false||Sulfonamide
null|Sulfonamides|Drug|false|false||Sulfonamide
null|Sulfonamide [EPC]|Drug|false|false||Sulfonamidenull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||Antibiotics
null|Antibiotics|Drug|false|false||Antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||Antibiotics
null|Antibiotics, Gynecological|Drug|false|false||Antibiotics
null|antibiotics, intestinal|Drug|false|false||Antibiotics
null|Antibiotic throat preparations|Drug|false|false||Antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||Antibiotics
null|Antibiotics for systemic use|Drug|false|false||Antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||Antibioticsnull|penicillins|Drug|false|false||Penicillins
null|penicillins|Drug|false|false||Penicillinsnull|Poisoning by, adverse effect of and underdosing of penicillins|Disorder|false|false||Penicillins
null|Poisoning by penicillin|Disorder|false|false||Penicillinsnull|Adverse reaction to penicillins|Finding|false|false||Penicillinsnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Chief complaint (finding)|Finding|false|false||Chief Complaintnull|Complaint (finding)|Finding|false|false||Complaintnull|null|Attribute|false|false||Complaintnull|Neck Pain|Finding|false|false|C0027530;C3159206|neck painnull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|neck
null|Neck problem|Finding|false|false|C0027530;C3159206|necknull|dendritic spine neck|Anatomy|false|false|C0007859;C1549543;C0030193;C0812434;C0684335|neck
null|Neck|Anatomy|false|false|C0007859;C1549543;C0030193;C0812434;C0684335|necknull|Administration Method - Pain|Finding|false|false|C0027530;C3159206|pain
null|Pain|Finding|false|false|C0027530;C3159206|painnull|null|Attribute|false|false||painnull|Falls|Finding|false|false||fallnull|Autumn|Time|false|false||fallnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|History of present illness (finding)|Finding|false|false||History of Present Illnessnull|null|Attribute|false|false||History of Present Illnessnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Present illness|Finding|false|false||Present Illnessnull|Present|Finding|false|false||Present
null|Presentation|Finding|false|false||Presentnull|Illness (finding)|Finding|false|false||Illnessnull|Male Gender|Finding|false|false||malenull|Male, Self-Reported|Subject|false|false||male
null|Males|Subject|false|false||malenull|Male Phenotype|Modifier|false|false||malenull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Processing type - Evaluation|Finding|false|false|C0027530|evaluationnull|Evaluation procedure|Procedure|false|false|C0027530|evaluation
null|Evaluation|Procedure|false|false|C0027530|evaluationnull|Neck|Anatomy|false|false|C1261322;C0220825;C1550157|cervicalnull|Cervical|Modifier|false|false||cervicalnull|Fracture|Disorder|false|false||fracturenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Bathroom|Device|false|false||bathroom
null|Toilet Facilities|Device|false|false||bathroomnull|Bent|Modifier|false|false||bentnull|Does hit (finding)|Finding|false|false||hittingnull|Struck by|Modifier|false|false||hittingnull|Problems with head|Disorder|false|false|C0018670;C0152336|headnull|Procedure on head|Procedure|false|false|C0018670;C0152336|headnull|Structure of head of caudate nucleus|Anatomy|false|false|C0362076;C0876917|head
null|Head|Anatomy|false|false|C0362076;C0876917|headnull|Head Device|Device|false|false||headnull|Unconscious State|Finding|true|false||loss of consciousnessnull|Loss (adaptation)|Finding|true|false||lossnull|Loss (quantitative)|LabModifier|false|false||lossnull|Consciousness related finding|Finding|false|false||consciousness
null|Conscious|Finding|false|false||consciousness
null|null|Finding|false|false||consciousnessnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Headache|Finding|false|false||headachenull|Neck Pain|Finding|false|false|C0027530;C3159206|neck painnull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|neck
null|Neck problem|Finding|false|false|C0027530;C3159206|necknull|dendritic spine neck|Anatomy|false|false|C0007859;C1549543;C0030193;C0812434;C0684335;C2598155|neck
null|Neck|Anatomy|false|false|C0007859;C1549543;C0030193;C0812434;C0684335;C2598155|necknull|Administration Method - Pain|Finding|false|false|C0027530;C3159206|pain
null|Pain|Finding|false|false|C0027530;C3159206|painnull|null|Attribute|false|false|C0027530;C3159206|painnull|Organization unit type - Hospital|Finding|false|false|C0018670;C0152336|hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Laceration of head|Disorder|false|false|C0018670;C0152336|head lacerationnull|Problems with head|Disorder|false|false|C0018670;C0152336|headnull|Procedure on head|Procedure|false|false|C0018670;C0152336|headnull|Structure of head of caudate nucleus|Anatomy|false|false|C0362076;C0043246;C1547192;C0876917;C0856548|head
null|Head|Anatomy|false|false|C0362076;C0043246;C1547192;C0876917;C0856548|headnull|Head Device|Device|false|false||headnull|Laceration|Disorder|false|false|C0018670;C0152336|lacerationnull|X-Ray Computed Tomography|Procedure|false|false||CT scannull|Radionuclide Imaging|Procedure|false|false||scan
null|Scanning|Procedure|false|false||scannull|Fracture|Disorder|false|false||fracturenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Numbness|Finding|true|false||numbness
null|Hypesthesia|Finding|true|false||numbnessnull|Paresthesia|Disorder|false|false|C0446516;C1140621|tinglingnull|Has tingling sensation|Finding|false|false|C1140621;C0446516|tinglingnull|Alveolar rhabdomyosarcoma|Disorder|false|false|C1140621;C0446516|armsnull|Adherence to Refills and Medications Scale|Finding|false|false|C0446516|arms
null|KIDINS220 gene|Finding|false|false|C0446516|armsnull|Upper arm|Anatomy|false|false|C0030554;C5575339;C2681631;C5782111;C2242996;C0206655|armsnull|null|Attribute|false|false|C0446516|armsnull|Leg|Anatomy|false|false|C0206655;C5781420;C2242996;C0030554|legsnull|null|Attribute|false|false|C1140621|legsnull|Weakness|Finding|true|false|C1140621;C0446516|weakness
null|Asthenia|Finding|true|false|C1140621;C0446516|weaknessnull|Alveolar rhabdomyosarcoma|Disorder|true|false|C1140621;C0446516|armsnull|Adherence to Refills and Medications Scale|Finding|true|false|C0446516|arms
null|KIDINS220 gene|Finding|true|false|C0446516|armsnull|Upper arm|Anatomy|false|false|C3714552;C0004093;C0206655;C5575339;C2681631;C5782111|armsnull|null|Attribute|true|false|C0446516|armsnull|Leg|Anatomy|false|false|C0206655;C3714552;C0004093;C5781420|legsnull|null|Attribute|false|false|C1140621|legsnull|Fecal Incontinence|Disorder|true|false|C0021853|bowel incontinencenull|Intestines|Anatomy|false|false|C0015732|bowelnull|Incontinence|Disorder|true|false||incontinencenull|Urinary Retention|Finding|true|false|C0005682|bladder retentionnull|Neoplasm of uncertain or unknown behavior of bladder|Disorder|true|false|C0005682|bladder
null|Benign neoplasm of bladder|Disorder|true|false|C0005682|bladder
null|Carcinoma in situ of bladder|Disorder|true|false|C0005682|bladdernull|Procedures on bladder|Procedure|true|false|C0005682|bladdernull|Urinary Bladder|Anatomy|false|false|C0496930;C0154017;C0154091;C0872388;C0080274|bladdernull|cellular entity retention|Finding|false|false||retention
null|Retention (Psychology)|Finding|false|false||retention
null|Urinary Retention|Finding|false|false||retention
null|Retention of content|Finding|false|false||retentionnull|Retention - dental|Attribute|false|false||retentionnull|Anesthesia substance|Drug|false|false||anesthesianull|null|Finding|false|false||anesthesia
null|Absence of sensation|Finding|false|false||anesthesianull|Anesthesia procedures|Procedure|false|false||anesthesia
null|Dental anesthesia|Procedure|false|false||anesthesianull|null|Attribute|false|false||anesthesianull|Chest Pain|Finding|true|false|C1527391;C0817096|chest painnull|null|Attribute|true|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0741025;C2926613;C0008031|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025;C2926613;C0008031|chestnull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Dyspnea|Finding|true|false||shortness of breathnull|null|Attribute|true|false||shortness of breathnull|Breath|Finding|false|false||breathnull|Abdominal Pain|Finding|false|false|C0000726|abdominal painnull|Abdomen|Anatomy|false|false|C1549543;C0030193;C0000737|abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Administration Method - Pain|Finding|false|false|C0000726|pain
null|Pain|Finding|false|false|C0000726|painnull|null|Attribute|false|false||painnull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|PMH - past medical history|Finding|false|false||PMH
null|Medical History|Finding|false|false||PMHnull|FBL gene|Finding|false|false||fibnull|Malignant tumor of colon|Disorder|false|false|C0009368;C4071907|colon canull|Neoplasm of uncertain or unknown behavior of colon|Disorder|false|false|C0009368;C4071907|colon
null|Colonic Diseases|Disorder|false|false|C0009368;C4071907|colon
null|Carcinoma in situ of colon|Disorder|false|false|C0009368;C4071907|colonnull|COLON PROBLEM|Finding|false|false|C0009368;C4071907|colonnull|Colon structure (body structure)|Anatomy|false|false|C0750873;C0007102;C0009373;C0154061;C0496907|colon
null|Abdomen+Pelvis>Colon|Anatomy|false|false|C0750873;C0007102;C0009373;C0154061;C0496907|colonnull|TUBE,COLON,22FR,RADIOPAQUE RUBBER B#7370|Device|false|false||colonnull|Colon <Coloninae>|Entity|false|false||colonnull|Hypertensive disease|Disorder|false|false||htnnull|COPD pharmacologic substance|Drug|false|false||copdnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||copd
null|Chronic Obstructive Airway Disease|Disorder|false|false||copdnull|ARCN1 gene|Finding|false|false||copdnull|Multiple Epiphyseal Dysplasia|Disorder|false|false||MEDnull|Master of Education|Finding|false|false||MED
null|COMP wt Allele|Finding|false|false||MED
null|COL9A3 gene|Finding|false|false||MED
null|SCN8A wt Allele|Finding|false|false||MED
null|COL9A2 gene|Finding|false|false||MED
null|COMP gene|Finding|false|false||MED
null|SCN8A gene|Finding|false|false||MEDnull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|allopurinol|Drug|false|false||allopurinol
null|allopurinol|Drug|false|false||allopurinolnull|Asacol|Drug|false|false||asacol
null|Asacol|Drug|false|false||asacolnull|Pregnenolone Carbonitrile|Drug|false|false||pcn
null|Pregnenolone Carbonitrile|Drug|false|false||pcnnull|PLEC wt Allele|Finding|false|false||pcn
null|PCNT gene|Finding|false|false||pcn
null|PLEC gene|Finding|false|false||pcnnull|sulfa|Drug|false|false||sulfanull|Social and personal history|Finding|false|false||Social History
null|Social History|Finding|false|false||Social Historynull|Social|Finding|false|false||Socialnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Family Medical History|Finding|false|false||Family Historynull|Entity Name Part Type - family|Finding|false|false||Family
null|Last Name|Finding|false|false||Family
null|Living Arrangement - Family|Finding|false|false||Family
null|Family (taxonomic)|Finding|false|false||Family
null|Family Collection|Finding|false|false||Familynull|Family|Subject|false|false||Familynull|History of present illness (finding)|Finding|false|true||History
null|History of previous events|Finding|false|true||History
null|Historical aspects qualifier|Finding|false|true||History
null|Medical History|Finding|false|true||History
null|Concept History|Finding|false|true||Historynull|History|Subject|false|false||Historynull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|Ostomy Collar|Device|false|false||collar
null|null|Device|false|false||collarnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|LAT protein, human|Drug|false|false||lat
null|L-Type Amino Acid Transporter|Drug|false|false||lat
null|L-Type Amino Acid Transporter|Drug|false|false||lat
null|ORC3 protein, human|Drug|false|false||lat
null|ORC3 protein, human|Drug|false|false||lat
null|LAT protein, human|Drug|false|false||latnull|LAT gene|Finding|false|false|C0446516;C1140618;C1269078|lat
null|ORC3 wt Allele|Finding|false|false|C0446516;C1140618;C1269078|lat
null|ORC3 gene|Finding|false|false|C0446516;C1140618;C1269078|lat
null|SPNS1 gene|Finding|false|false|C0446516;C1140618;C1269078|latnull|Latin Language|Entity|false|false||latnull|Anorectal Malformations|Disorder|false|false|C0446516;C1140618;C1269078|armnull|AKR1A1 wt Allele|Finding|false|false|C0446516;C1140618;C1269078|arm
null|ARMC9 gene|Finding|false|false|C0446516;C1140618;C1269078|armnull|Protocol Treatment Arm|Procedure|false|false|C0446516;C1140618;C1269078|arm
null|Axillary Reverse Mapping|Procedure|false|false|C0446516;C1140618;C1269078|arm
null|Study Arm|Procedure|false|false|C0446516;C1140618;C1269078|armnull|Upper arm|Anatomy|false|false|C1705279;C1335085;C1425844;C2240043;C1824218;C3715044;C1522541;C5400986;C4761640;C3495676|arm
null|null|Anatomy|false|false|C1705279;C1335085;C1425844;C2240043;C1824218;C3715044;C1522541;C5400986;C4761640;C3495676|arm
null|Upper Extremity|Anatomy|false|false|C1705279;C1335085;C1425844;C2240043;C1824218;C3715044;C1522541;C5400986;C4761640;C3495676|armnull|Thumb structure|Anatomy|false|false||thumbnull|Middle|Modifier|false|false||midnull|Upper extremity>Finger|Anatomy|false|false||finger
null|Fingers|Anatomy|false|false||finger
null|Fingers not including thumb|Anatomy|false|false||fingernull|Multiple Epiphyseal Dysplasia|Disorder|false|false|C0446516;C1140618;C1269078|mednull|Master of Education|Finding|false|false|C0446516;C1140618;C1269078|med
null|COMP wt Allele|Finding|false|false|C0446516;C1140618;C1269078|med
null|COL9A3 gene|Finding|false|false|C0446516;C1140618;C1269078|med
null|SCN8A wt Allele|Finding|false|false|C0446516;C1140618;C1269078|med
null|COL9A2 gene|Finding|false|false|C0446516;C1140618;C1269078|med
null|COMP gene|Finding|false|false|C0446516;C1140618;C1269078|med
null|SCN8A gene|Finding|false|false|C0446516;C1140618;C1269078|mednull|Anorectal Malformations|Disorder|false|false|C0446516;C1140618;C1269078|armnull|AKR1A1 wt Allele|Finding|false|false|C0446516;C1140618;C1269078|arm
null|ARMC9 gene|Finding|false|false|C0446516;C1140618;C1269078|armnull|Protocol Treatment Arm|Procedure|false|false|C0446516;C1140618;C1269078|arm
null|Axillary Reverse Mapping|Procedure|false|false|C0446516;C1140618;C1269078|arm
null|Study Arm|Procedure|false|false|C0446516;C1140618;C1269078|armnull|Upper arm|Anatomy|false|false|C3495676;C0026760;C1824218;C3715044;C1522541;C5400986;C4761640;C4321267;C1419866;C1549978;C5781216;C1456376;C1413596;C1413597|arm
null|null|Anatomy|false|false|C3495676;C0026760;C1824218;C3715044;C1522541;C5400986;C4761640;C4321267;C1419866;C1549978;C5781216;C1456376;C1413596;C1413597|arm
null|Upper Extremity|Anatomy|false|false|C3495676;C0026760;C1824218;C3715044;C1522541;C5400986;C4761640;C4321267;C1419866;C1549978;C5781216;C1456376;C1413596;C1413597|armnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Trunk of elephant|Anatomy|false|false||Trunk
null|Trunk structure|Anatomy|false|false||Trunk
null|dendritic shaft|Anatomy|false|false||Trunknull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Pelvis>Groin|Anatomy|false|false|C0562271|Groin
null|Inguinal region|Anatomy|false|false|C0562271|Groin
null|Inguinal part of abdomen|Anatomy|false|false|C0562271|Groinnull|Examination of knee joint|Procedure|false|false|C0816951;C4266533;C0018246;C1963703;C0022742;C4299094;C0022745|Kneenull|Knee region structure|Anatomy|false|false|C0562271|Knee
null|Knee|Anatomy|false|false|C0562271|Knee
null|Lower extremity>Knee|Anatomy|false|false|C0562271|Knee
null|Knee joint|Anatomy|false|false|C0562271|Kneenull|Multiple Epiphyseal Dysplasia|Disorder|false|false|C0230445;C1305418|Mednull|Master of Education|Finding|false|false|C0230445;C1305418|Med
null|COMP wt Allele|Finding|false|false|C0230445;C1305418|Med
null|COL9A3 gene|Finding|false|false|C0230445;C1305418|Med
null|SCN8A wt Allele|Finding|false|false|C0230445;C1305418|Med
null|COL9A2 gene|Finding|false|false|C0230445;C1305418|Med
null|COMP gene|Finding|false|false|C0230445;C1305418|Med
null|SCN8A gene|Finding|false|false|C0230445;C1305418|Mednull|Structure of calf of leg|Anatomy|false|false|C4321267;C1419866;C1549978;C5781216;C1456376;C1413596;C1413597;C0026760|Calf
null|null|Anatomy|false|false|C4321267;C1419866;C1549978;C5781216;C1456376;C1413596;C1413597;C0026760|Calfnull|Cattle calf (organism)|Entity|false|false||Calfnull|Clava structure (body structure)|Anatomy|false|false||Grtnull|Lower extremity>Toes|Anatomy|false|false||Toe
null|Toes|Anatomy|false|false||Toenull|Lower extremity>Toes|Anatomy|false|false||Toe
null|Toes|Anatomy|false|false||Toenull|Lower extremity>Thigh|Anatomy|false|false||Thigh
null|Thigh structure|Anatomy|false|false||Thighnull|motor movement|Finding|false|false||Motornull|Motor Device|Device|false|false||Motornull|imidazole mustard|Drug|false|false|C3495985;C0175372|Bic
null|imidazole mustard|Drug|false|false|C3495985;C0175372|Bicnull|MIR155HG gene|Finding|false|false|C3495985;C0175372|Bic
null|MIR155 gene|Finding|false|false|C3495985;C0175372|Bicnull|BIC Regimen|Procedure|false|false|C3495985;C0175372|Bicnull|Structure of inferior brachium of corpora quadrigemina|Anatomy|false|false|C0063382;C1537811;C2681931;C5202575|Bic
null|nucleus of the brachium of the inferior colliculus|Anatomy|false|false|C0063382;C1537811;C2681931;C5202575|Bicnull|TRI-AAT9-1 gene|Finding|false|false||Tri
null|Temptation and Restraint Inventory|Finding|false|false||Trinull|Babinski Reflex|Finding|false|false||Babinskinull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Clonus|Finding|false|false||Clonusnull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|BRIEF Health Literacy Screening Tool|Finding|false|false||Brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||Briefnull|Brief|Time|false|false||Briefnull|Shortened|Modifier|false|false||Briefnull|Hospital course|Finding|false|false||Hospital Coursenull|null|Attribute|false|false||Hospital Coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||Coursenull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Level of Care - Surgery|Finding|false|false||Surgery
null|Surgical procedure finding|Finding|false|false||Surgery
null|Surgical aspects|Finding|false|false||Surgerynull|Operative Surgical Procedures|Procedure|false|false||Surgerynull|General surgery specialty|Title|false|false||Surgery
null|Surgery specialty|Title|false|false||Surgerynull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Examination and observation for unspecified reason|Finding|false|false||observation
null|null|Finding|false|false||observation
null|null|Finding|false|false||observation
null|Observation (finding)|Finding|false|false||observationnull|Observation - diagnostic procedure|Procedure|false|false||observation
null|Observation in research|Procedure|false|false||observation
null|Patient observation|Procedure|false|false||observationnull|Fracture|Disorder|false|false||fracturenull|Postoperative deep vein thrombosis|Disorder|false|false|C5239664|postoperative DVTnull|Postoperative Period|Time|false|false||postoperativenull|DVT prophylaxis|Procedure|false|false|C5239664|DVT prophylaxisnull|Deep thrombophlebitis|Disorder|false|false|C5239664|DVT
null|Deep Vein Thrombosis|Disorder|false|false|C5239664|DVTnull|area DVT|Anatomy|false|false|C0853245;C0589110;C2926618;C0199176;C0149871;C0151950|DVTnull|null|Attribute|false|false|C5239664|DVTnull|Prophylactic treatment|Procedure|false|false|C5239664|prophylaxisnull|prevention & control|Modifier|false|false||prophylaxisnull|Diet (animal life circumstance)|Drug|false|false||Diet
null|Diet|Drug|false|false||Dietnull|diet - supply|Finding|false|false||Dietnull|Diet therapy|Procedure|false|false||Dietnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Oral pain|Finding|false|false|C0226896|oral painnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C0221776;C1527415;C4521986;C3244316;C4284232;C1549543;C0030193;C1272919|oralnull|Oral|Modifier|false|false||oralnull|Administration Method - Pain|Finding|false|false|C0226896|pain
null|Pain|Finding|false|false|C0226896|painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false|C0226896|medication
null|Medications|Finding|false|false|C0226896|medicationnull|Diagnostic Service Section ID - Physical Therapy|Finding|false|false||Physical therapynull|Physical therapy|Procedure|false|false||Physical therapynull|Physical therapy (field)|Title|false|false||Physical therapynull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|physical therapy mobilization (treatment)|Procedure|false|false||mobilization
null|Mobilization (procedure)|Procedure|false|false||mobilizationnull|Ambulate|Finding|false|false||ambulatenull|Hypertensive (finding)|Finding|false|false||hypertensivenull|MEDICINE CONSULT|Procedure|false|false||Medicine consultnull|Pharmaceutical Preparations|Drug|false|false||Medicinenull|Medicine|Title|false|false||Medicinenull|Consultation|Procedure|false|false||consultnull|Long Variable|Modifier|false|false||long
null|Long|Modifier|false|false||longnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Antihypertensive Agents|Drug|false|false||antihypertensivesnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Too low|Finding|false|false||too lownull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Too quickly|Finding|false|false||too quicklynull|Hospital course|Finding|false|false||Hospital coursenull|null|Attribute|false|false||Hospital coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||coursenull|null|Modifier|false|false||unremarkablenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Apyrexial|Finding|false|false||afebrilenull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Taking vital signs|Procedure|false|false||vital signsnull|null|Attribute|false|false||vital signs
null|Vital signs|Attribute|false|false||vital signsnull|Vital High Nitrogen Enteral Nutrition|Drug|false|false||vitalnull|Vital (qualifier value)|Modifier|false|false||vitalnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Feeling comfortable|Finding|false|false||comfortablenull|Oral pain|Finding|false|false|C0226896|oral painnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C0221776;C1272919;C1527415;C4521986|oralnull|Oral|Modifier|false|false||oralnull|Demonstrates adequate pain control|Finding|false|false||pain controlnull|Pain control|Procedure|false|false||pain control
null|Pain management (procedure)|Procedure|false|false||pain controlnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Control brand of phenylpropanolamine|Drug|false|false||control
null|CONTROL veterinary product|Drug|false|false||control
null|control substance|Drug|false|false||control
null|Control brand of phenylpropanolamine|Drug|false|false||controlnull|Control - Relationship modifier|Finding|false|false||control
null|Control function|Finding|false|false||control
null|Scientific Control|Finding|false|false||controlnull|Control Groups|Subject|false|false||controlnull|True Control Status|Modifier|false|false||control
null|control aspects|Modifier|false|false||controlnull|null|Finding|false|false||regular dietnull|Regular|Modifier|false|false||regularnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every four hours|Time|false|false||Q4Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|C1orf210 gene|Finding|false|false||tempnull|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Procedure|false|false||tempnull|Temperature|LabModifier|false|false||tempnull|Headache|Finding|false|false||headachenull|allopurinol|Drug|false|false||Allopurinol
null|allopurinol|Drug|false|false||Allopurinolnull|Daily|Time|false|false||DAILYnull|mesalamine|Drug|false|false||Mesalamine
null|mesalamine|Drug|false|false||Mesalaminenull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|metoprolol tartrate|Drug|false|false||Metoprolol Tartrate
null|metoprolol tartrate|Drug|false|false||Metoprolol Tartratenull|metoprolol|Drug|false|false||Metoprolol
null|metoprolol|Drug|false|false||Metoprololnull|tartrate|Drug|false|false||Tartrate
null|Tartrates|Drug|false|false||Tartrate
null|tartrate|Drug|false|false||Tartratenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|omeprazole|Drug|false|false||Omeprazole
null|omeprazole|Drug|false|false||Omeprazolenull|Daily|Time|false|false||DAILYnull|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarinnull|Daily|Time|false|false||DAILYnull|oxycodone|Drug|false|false||OxycoDONE
null|oxycodone|Drug|false|false||OxycoDONEnull|Oxycodone measurement|Procedure|false|false||OxycoDONEnull|Immediate Release Dosage Form|Drug|false|false||Immediate Releasenull|Query Priority - Immediate|Finding|false|false||Immediate
null|immediate - ResponseCode|Finding|false|false||Immediatenull|Immediate|Time|false|false||Immediate
null|Stat (do immediately)|Time|false|false||Immediatenull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Every four hours|Time|false|false||Q4Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|diazepam|Drug|false|false||Diazepam
null|diazepam|Drug|false|false||Diazepamnull|Every twelve hours|Time|false|false||Q12Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Spasm|Finding|false|false||spasmsnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Fracture|Disorder|false|false||fracturenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Disease|Disorder|false|false||Conditionnull|Logical Condition|Finding|false|false||Conditionnull|null|Attribute|false|false||Conditionnull|Condition|Modifier|false|false||Conditionnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|Discharge instructions|Finding|false|false||Discharge Instructionsnull|hospital discharge instructions (treatment)|Procedure|false|false||Discharge Instructionsnull|null|Attribute|false|false||Discharge Instructionsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|Following|Time|false|false||following
null|Status post|Time|false|false||followingnull|Computer Operation|Procedure|false|false||operation
null|Operative Surgical Procedures|Procedure|false|false||operationnull|Operation Activity|Event|false|false||operationnull|Anterior cervical spine approach|Modifier|false|false||Anterior Cervicalnull|Adenohypophyseal Diseases|Disorder|false|false|C0027530|Anteriornull|Anterior|Modifier|false|false||Anteriornull|Neck|Anatomy|false|false|C0751437|Cervicalnull|Cervical|Modifier|false|false||Cervicalnull|Decompression - action (qualifier value)|Finding|false|false||Decompressionnull|Decompression|Procedure|false|false||Decompression
null|Decompressive incision|Procedure|false|false||Decompressionnull|external decompression|Phenomenon|false|false||Decompressionnull|Fused structure|Finding|false|false||Fusionnull|Fusion procedure|Procedure|false|false||Fusionnull|Stat (do immediately)|Time|false|false||Immediatelynull|Computer Operation|Procedure|false|false||operation
null|Operative Surgical Procedures|Procedure|false|false||operationnull|Operation Activity|Event|false|false||operationnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|Greater Than|LabModifier|false|false||greater thannull|Greater|LabModifier|false|false||greaternull|liquid-based cytology (procedure)|Procedure|false|false||lbsnull|Pounds|LabModifier|false|false||lbsnull|2 Weeks|Time|false|false||2 weeksnull|week|Time|false|false||weeksnull|More|LabModifier|false|false||morenull|Feeling comfortable|Finding|false|false||comfortablenull|Coxsackievirus and Adenovirus Receptor, human|Drug|false|false|C1166663|car
null|Coxsackievirus and Adenovirus Receptor, human|Drug|false|false|C1166663|car
null|Chimeric antigen receptor|Drug|false|false|C1166663|car
null|Chimeric antigen receptor|Drug|false|false|C1166663|car
null|Extracellular Calcium-Sensing Receptor, Human|Drug|false|false|C1166663|carnull|Carney Complex|Disorder|false|false|C1166663|carnull|Car - Mode of Arrival Code|Finding|false|false|C1166663|car
null|Chimeric antigen receptor|Finding|false|false|C1166663|car
null|CASR wt Allele|Finding|false|false|C1166663|car
null|Extracellular Calcium-Sensing Receptor, Human|Finding|false|false|C1166663|car
null|CXADR wt Allele|Finding|false|false|C1166663|car
null|CXADR gene|Finding|false|false|C1166663|car
null|PRKAR1A wt Allele|Finding|false|false|C1166663|car
null|CXADRP1 gene|Finding|false|false|C1166663|car
null|NR1I3 gene|Finding|false|false|C1166663|car
null|SPG7 gene|Finding|false|false|C1166663|car
null|TRIM13 wt Allele|Finding|false|false|C1166663|car
null|Caronte Gene|Finding|false|false|C1166663|car
null|SPG7 wt Allele|Finding|false|false|C1166663|car
null|NR1I3 wt Allele|Finding|false|false|C1166663|carnull|actomyosin contractile ring|Anatomy|false|false|C3539542;C4039583;C5890846;C3540475;C1547285;C3273602;C4039583;C1413828;C3811749;C2239319;C1858724;C1417827;C5890847;C1420354;C5960871;C1706434;C5890846;C0406810|carnull|Automobiles|Device|false|false||carnull|Car <Caridae>|Entity|false|false||car
null|Carib language|Entity|false|false||carnull|Chairs|Device|false|false||chairnull|Chairperson|Subject|false|false||chairnull|Greater Than|LabModifier|false|false||more thannull|More|LabModifier|false|false||morenull|45 Minutes|Time|false|false||45 minutesnull|Minute of time|Time|false|false||minutesnull|Minute Unit of Plane Angle|LabModifier|false|false||minutes
null|Minute (diminutive)|LabModifier|false|false||minutes
null|Small|LabModifier|false|false||minutesnull|Encounter due to care involving use of rehabilitation procedures|Finding|false|false||Rehabilitation
null|Rehabilitation aspects|Finding|false|false||Rehabilitationnull|Rehabilitation therapy|Procedure|false|false||Rehabilitationnull|null|Title|false|false||Rehabilitationnull|Diagnostic Service Section ID - Physical Therapy|Finding|false|false||Physical Therapynull|Physical therapy|Procedure|false|false||Physical Therapynull|Physical therapy (field)|Title|false|false||Physical Therapynull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Therapy Object (animal model)|Finding|false|false||Therapy
null|therapeutic aspects|Finding|false|false||Therapynull|Therapeutic procedure|Procedure|false|false||Therapynull|3 times|Finding|false|false||3 timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Walking (function)|Finding|false|false||walknull|Minute of time|Time|false|false||minutesnull|Minute Unit of Plane Angle|LabModifier|false|false||minutes
null|Minute (diminutive)|LabModifier|false|false||minutes
null|Small|LabModifier|false|false||minutesnull|part of|Modifier|false|false||part ofnull|Role Class - part|Finding|false|false||partnull|Part|Modifier|false|false||partnull|Part Dosing Unit|LabModifier|false|false||partnull|Recovery - healing process|Finding|false|false||recoverynull|null|Event|false|false||recoverynull|recovery - adjustment|LabModifier|false|false||recoverynull|Much|Finding|false|false||muchnull|Telephone Extension Number|Finding|false|false||Extension
null|Extension|Finding|false|false||Extensionnull|Exercise|Finding|false|false||Exercisenull|Exercise Pain Management|Procedure|false|false||Exercisenull|Ostomy Collar|Device|false|false||collar
null|null|Device|false|false||collarnull|per day|Time|false|false||/daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Swallowing G-code|Finding|false|false||Swallowing
null|Does swallow|Finding|false|false||Swallowing
null|Deglutition|Finding|false|false||Swallowingnull|outcomes otolaryngology swallowing (treatment)|Procedure|false|false||Swallowingnull|null|Attribute|false|false||Swallowingnull|Deglutition Disorders|Disorder|true|false||Difficulty swallowingnull|Has difficulty doing (qualifier value)|Finding|false|false||Difficultynull|Swallowing G-code|Finding|false|false||swallowing
null|Does swallow|Finding|false|false||swallowing
null|Deglutition|Finding|false|false||swallowingnull|outcomes otolaryngology swallowing (treatment)|Procedure|false|false||swallowingnull|null|Attribute|false|false||swallowingnull|Rare|Modifier|false|false||uncommonnull|Type - ParameterizedDataType|Finding|false|false||type
null|SGCG gene|Finding|false|false||typenull|null|Modifier|false|false||typenull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Small|LabModifier|false|false||smallnull|bite injury|Disorder|false|false||bitesnull|Slow|Modifier|false|false||slowlynull|Ostomy Collar|Device|false|false||collar
null|null|Device|false|false||collarnull|Helpful|Modifier|false|false||helpfulnull|Movement|Finding|false|false||movementnull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|neck
null|Neck problem|Finding|false|false|C0027530;C3159206|necknull|dendritic spine neck|Anatomy|false|false|C0812434;C0684335|neck
null|Neck|Anatomy|false|false|C0812434;C0684335|necknull|Ostomy Collar|Device|false|false||collar
null|null|Device|false|false||collarnull|null|Device|false|false||Cervical Collarnull|Neck|Anatomy|false|false|C1828220|Cervicalnull|Cervical|Modifier|false|false||Cervicalnull|Ostomy Collar|Device|false|false||Collar
null|null|Device|false|false||Collarnull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|Neck
null|Neck problem|Finding|false|false|C0027530;C3159206|Necknull|dendritic spine neck|Anatomy|false|false|C1828220;C0812434;C0684335|Neck
null|Neck|Anatomy|false|false|C1828220;C0812434;C0684335|Necknull|Application of brace (procedure)|Procedure|false|false|C0027530;C0027530;C3159206|Bracenull|Braces - Orthopedic appliances|Device|false|false||Brace
null|Braces - garment|Device|false|false||Bracenull|Application of brace (procedure)|Procedure|false|false||bracenull|Braces - Orthopedic appliances|Device|false|false||brace
null|Braces - garment|Device|false|false||bracenull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Follow-up status|Finding|false|false||follow-upnull|follow-up|Procedure|false|false||follow-upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|Appointments|Event|false|false||appointmentnull|week|Time|false|false||weeksnull|Ostomy Collar|Device|false|false||collar
null|null|Device|false|false||collarnull|take a shower|Finding|false|false||take a showernull|Shower (physical object)|Device|false|false||showernull|Motion|Phenomenon|false|false|C0027530;C3159206|motionnull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|neck
null|Neck problem|Finding|false|false|C0027530;C3159206|necknull|dendritic spine neck|Anatomy|false|false|C0812434;C0684335;C0026597|neck
null|Neck|Anatomy|false|false|C0812434;C0684335;C0026597|necknull|Ostomy Collar|Device|false|false||collar
null|null|Device|false|false||collarnull|Place - dosing instruction imperative|Finding|false|false||Placenull|null|Procedure|false|false||Placenull|put - instruction imperative|Event|false|false||Placenull|Place|Modifier|false|false||Placenull|Ostomy Collar|Device|false|false||collar
null|null|Device|false|false||collarnull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|neck
null|Neck problem|Finding|false|false|C0027530;C3159206|necknull|dendritic spine neck|Anatomy|false|false|C0812434;C0684335|neck
null|Neck|Anatomy|false|false|C0812434;C0684335|necknull|Stat (do immediately)|Time|false|false||immediatelynull|Shower (physical object)|Device|false|false||showernull|Wound care management|Procedure|false|false||Wound Care
null|wound care|Procedure|false|false||Wound Carenull|Wound Care kit|Device|false|false||Wound Carenull|Traumatic Wound|Disorder|false|false||Wound
null|Wounds and Injuries|Disorder|false|false||Wound
null|Traumatic injury|Disorder|false|false||Woundnull|Route of Administration - Wound|Finding|false|false||Wound
null|null|Finding|false|false||Wound
null|Specimen Type - Wound|Finding|false|false||Woundnull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|Laceration|Disorder|false|false|C0036270|lacerationnull|Scalp structure|Anatomy|false|false|C0041834;C0013103;C0043246|scalpnull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false|C0036270|drainagenull|Erythema|Disorder|false|false|C0036270|rednessnull|Redness|Finding|false|false||rednessnull|Red color|Modifier|false|false||rednessnull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Staple, Surgical|Device|false|false||staplesnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Additional|Finding|false|false||Additionalnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|Control brand of phenylpropanolamine|Drug|false|false||control
null|CONTROL veterinary product|Drug|false|false||control
null|control substance|Drug|false|false||control
null|Control brand of phenylpropanolamine|Drug|false|false||controlnull|Control - Relationship modifier|Finding|false|false||control
null|Control function|Finding|false|false||control
null|Scientific Control|Finding|false|false||controlnull|Control Groups|Subject|false|false||controlnull|True Control Status|Modifier|false|false||control
null|control aspects|Modifier|false|false||controlnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|72 Hours|Time|false|false||72 hoursnull|Hour|Time|false|false||hoursnull|refill|Finding|false|false||refillnull|Narcotics|Drug|false|false||narcotic
null|Narcotics|Drug|false|false||narcoticnull|Prescription (procedure)|Procedure|false|false||prescriptionsnull|null|Attribute|false|false||prescriptionsnull|Infantile Neuroaxonal Dystrophy|Disorder|false|false||plannull|Treatment Plan|Finding|false|false||plan
null|Planned|Finding|false|false||plan
null|null|Finding|false|false||plannull|Mail|Device|false|false||mailednull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Clinic|Device|false|false||clinic
null|Ambulatory Care Facilities|Device|false|false||clinicnull|Clinic|Entity|false|false||clinic
null|Ambulatory Care Facilities|Entity|false|false||clinicnull|Patient location type - Clinic|Modifier|false|false||clinic
null|Person location type - Clinic|Modifier|false|false||clinicnull|Narcotics|Drug|false|false||narcotic
null|Narcotics|Drug|false|false||narcoticnull|Oxycontin|Drug|false|false||oxycontin
null|Oxycontin|Drug|false|false||oxycontinnull|oxycodone|Drug|false|false||oxycodone
null|oxycodone|Drug|false|false||oxycodonenull|Oxycodone measurement|Procedure|false|false||oxycodonenull|Percocet|Drug|false|false||percocet
null|Percocet|Drug|false|false||percocetnull|Prescription (procedure)|Procedure|false|false||prescriptionsnull|null|Attribute|false|false||prescriptionsnull|Diagnostic Service Section ID - Pharmacy|Finding|false|false||pharmacy
null|Pharmacy domain|Finding|false|false||pharmacynull|Pharmaceutical Services|Procedure|false|false||pharmacynull|Pharmacy facility|Device|false|false||pharmacynull|Pharmacy (field)|Title|false|false||pharmacynull|Pharmacy facility|Entity|false|false||pharmacynull|In addition to|Finding|false|false||addition
null|Add - instruction imperative|Finding|false|false||additionnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|90 days|Time|false|false||90 daysnull|day|Time|false|false||daysnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Follow-up status|Finding|false|false||Follow upnull|follow-up|Procedure|false|false||Follow upnull|Follow - dosing instruction imperative|Finding|false|false||Follow
null|Follow|Finding|false|false||Follownull|Followed by|Time|false|false||Follownull|Address type - Office|Finding|false|false||officenull|Office|Device|false|false||officenull|Organization unit type - Office|Entity|false|false||officenull|Appointments|Event|false|false||appointmentnull|2 Weeks|Time|false|false||2 weeksnull|week|Time|false|false||weeksnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Computer Operation|Procedure|false|false||operation
null|Operative Surgical Procedures|Procedure|false|false||operationnull|Operation Activity|Event|false|false||operationnull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Visit|Finding|false|false||visitnull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0332803;C0184898|incisionnull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Plain x-ray|Procedure|false|false||x raysnull|Roentgen Rays|Phenomenon|false|false||x raysnull|Radiation|Phenomenon|false|false||raysnull|Rajiformes|Entity|false|false||raysnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|6 weeks|Time|false|false||6 weeksnull|week|Time|false|false||weeksnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Computer Operation|Procedure|false|false||operation
null|Operative Surgical Procedures|Procedure|false|false||operationnull|Operation Activity|Event|false|false||operationnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|most likely|Finding|false|false||most likelynull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Flexion/extension|Modifier|false|false||Flexion/Extensionnull|null|Finding|false|false||Flexionnull|W flexion|Attribute|false|false||Flexionnull|Telephone Extension Number|Finding|false|false||Extension
null|Extension|Finding|false|false||Extensionnull|X-rays, Homeopathic Preparations|Drug|false|false||X-raysnull|Plain x-ray|Procedure|false|false||X-rays
null|Diagnostic radiologic examination|Procedure|false|false||X-raysnull|Roentgen Rays|Phenomenon|false|false||X-raysnull|Often - answer to question|Finding|false|false||oftennull|Frequently|Time|false|false||oftennull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|Ostomy Collar|Device|false|false||collar
null|null|Device|false|false||collarnull|1 Week|Time|false|false||1 weeknull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Address type - Office|Finding|false|false||officenull|Office|Device|false|false||officenull|Organization unit type - Office|Entity|false|false||officenull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Academic degree|Finding|false|false||degreesnull|Degree or extent|LabModifier|false|false||degreesnull|Degrees fahrenheit|LabModifier|false|false||Fahrenheitnull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|Traumatic Wound|Disorder|false|false||wound
null|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|Diagnostic Service Section ID - Physical Therapy|Finding|false|false||Physical Therapynull|Physical therapy|Procedure|false|false||Physical Therapynull|Physical therapy (field)|Title|false|false||Physical Therapynull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Therapy Object (animal model)|Finding|false|false||Therapy
null|therapeutic aspects|Finding|false|false||Therapynull|Therapeutic procedure|Procedure|false|false||Therapynull|Activity (animal life circumstance)|Finding|false|false||activity
null|Physical activity|Finding|false|false||activitynull|Activities|Event|false|false||activitynull|null|Modifier|false|false||activitynull|Ostomy Collar|Device|false|false||collar
null|null|Device|false|false||collarnull|Full-time employment (finding)|Finding|false|false||full timenull|Full|Modifier|false|false||fullnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|week|Time|false|false||weeksnull|Referral category - Ambulatory|Finding|false|false||ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||ambulatory
null|Ambulatory|Finding|false|false||ambulatory
null|Level of Care - Ambulatory|Finding|false|false||ambulatorynull|ambulatory encounter|Procedure|false|false||ambulatorynull|Specialty Type - Ambulatory|Title|false|false||ambulatorynull|Self-Help Devices|Device|false|false||assistive devicesnull|Medical Devices|Device|false|false||devices
null|device aspects|Device|false|false||devices
null|Devices|Device|false|false||devicesnull|Safety|Phenomenon|false|false||safetynull|Decompression Sickness|Disorder|false|false||bendingnull|Bending - Changing basic body position|Finding|false|false||bending
null|Does bend|Finding|false|false||bendingnull|Bent|Modifier|false|false||bendingnull|Musculoskeletal torsion (function)|Finding|true|false||twisting
null|Torsion (malposition)|Finding|true|false||twistingnull|Biomaterial Treatment|Finding|false|false||Treatment
null|Treating|Finding|false|false||Treatment
null|therapeutic aspects|Finding|false|false||Treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||Treatment
null|Administration (procedure)|Procedure|false|false||Treatment
null|Therapeutic procedure|Procedure|false|false||Treatmentnull|Frequency|Finding|false|false||Frequency
null|How Often|Finding|false|false||Frequencynull|With frequency|Time|false|false||Frequency
null|Frequencies (time pattern)|Time|false|false||Frequencynull|Kind of quantity - Frequency|LabModifier|false|false||Frequency
null|Statistical Frequency|LabModifier|false|false||Frequency
null|Spatial Frequency|LabModifier|false|false||Frequencynull|Monitor brand of insecticide|Drug|false|false|C1123023;C4520765|monitor
null|Monitor brand of insecticide|Drug|false|false|C1123023;C4520765|monitornull|Monitor Device|Device|false|false||monitor
null|Monitoring Device|Device|false|false||monitornull|Monitor, occupation|Subject|false|false||monitornull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765;C0008114;C0018670;C0152336;C0230005|skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765;C0008114;C0018670;C0152336;C0230005|skinnull|Skin Specimen Source Code|Finding|false|false|C0018670;C0152336;C1123023;C4520765;C0230005;C0008114|skin
null|Skin Specimen|Finding|false|false|C0018670;C0152336;C1123023;C4520765;C0230005;C0008114|skinnull|Skin, Human|Anatomy|false|false|C0178298;C0496955;C1546781;C0444099;C0728873;C0362076|skin
null|Skin|Anatomy|false|false|C0178298;C0496955;C1546781;C0444099;C0728873;C0362076|skinnull|examination of chin|Procedure|false|false|C0008114;C0230005|chinnull|Chin|Anatomy|false|false|C2226982;C0178298;C0496955;C0362076;C1546781;C0444099|chinnull|Occipital region|Anatomy|false|false|C2226982;C0699900;C0362076;C1546781;C0444099;C1265875;C0178298;C0496955;C0876917|back of headnull|Problems with head|Disorder|false|false|C0018670;C0152336;C0230005;C0008114;C1123023;C4520765|headnull|Procedure on head|Procedure|false|false|C0018670;C0152336;C0230005|headnull|Structure of head of caudate nucleus|Anatomy|false|false|C1546781;C0444099;C0362076;C0876917;C1265875;C0178298;C0496955;C0699900|head
null|Head|Anatomy|false|false|C1546781;C0444099;C0362076;C0876917;C1265875;C0178298;C0496955;C0699900|headnull|Head Device|Device|false|false||headnull|Disintegration (morphologic abnormality)|Disorder|false|false|C0230005;C0018670;C0152336|breakdownnull|Catabolism|Finding|false|false|C0230005;C0018670;C0152336|breakdownnull|Ostomy Collar|Device|false|false||collar
null|null|Device|false|false||collarnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions