 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|32,36
No|37,39
:|39,40
_|43,44
_|44,45
_|45,46
<EOL>|46,47
<EOL>|48,49
Admission|49,58
Date|59,63
:|63,64
_|66,67
_|67,68
_|68,69
Discharge|83,92
Date|93,97
:|97,98
_|101,102
_|102,103
_|103,104
<EOL>|104,105
<EOL>|106,107
Date|107,111
of|112,114
Birth|115,120
:|120,121
_|123,124
_|124,125
_|125,126
Sex|139,142
:|142,143
M|146,147
<EOL>|147,148
<EOL>|149,150
Service|150,157
:|157,158
MEDICINE|159,167
<EOL>|167,168
<EOL>|169,170
Allergies|170,179
:|179,180
<EOL>|181,182
No|182,184
Known|185,190
Allergies|191,200
/|201,202
Adverse|203,210
Drug|211,215
Reactions|216,225
<EOL>|225,226
<EOL>|227,228
Attending|228,237
:|237,238
_|239,240
_|240,241
_|241,242
.|242,243
<EOL>|243,244
<EOL>|245,246
Chief|246,251
Complaint|252,261
:|261,262
<EOL>|262,263
Visual|263,269
hallucinations|270,284
<EOL>|284,285
<EOL>|286,287
Major|287,292
Surgical|293,301
or|302,304
Invasive|305,313
Procedure|314,323
:|323,324
<EOL>|324,325
N|325,326
/|326,327
A|327,328
<EOL>|328,329
<EOL>|329,330
<EOL>|331,332
History|332,339
of|340,342
Present|343,350
Illness|351,358
:|358,359
<EOL>|359,360
_|360,361
_|361,362
_|362,363
male|364,368
with|369,373
_|374,375
_|375,376
_|376,377
disease|378,385
,|385,386
dyslipidemia|387,399
,|399,400
and|401,404
a|405,406
<EOL>|406,407
history|407,414
of|415,417
prostate|418,426
cancer|427,433
(|434,435
s|435,436
/|436,437
p|437,438
prostatectomy|439,452
)|452,453
who|454,457
was|458,461
referred|462,470
<EOL>|470,471
to|471,473
the|474,477
ED|478,480
by|481,483
his|484,487
neurologist|488,499
for|500,503
worsening|504,513
gait|514,518
,|518,519
falls|520,525
,|525,526
and|527,530
<EOL>|530,531
visual|531,537
hallucinations|538,552
.|552,553
<EOL>|554,555
<EOL>|555,556
The|556,559
following|560,569
history|570,577
is|578,580
taken|581,586
from|587,591
chart|592,597
review|598,604
:|604,605
<EOL>|606,607
<EOL>|607,608
The|608,611
patient|612,619
was|620,623
seen|624,628
by|629,631
his|632,635
neurologist|636,647
on|648,650
_|651,652
_|652,653
_|653,654
at|655,657
which|658,663
time|664,668
he|669,671
<EOL>|671,672
was|672,675
noted|676,681
to|682,684
have|685,689
visual|690,696
hallucinations|697,711
and|712,715
worsening|716,725
gait|726,730
<EOL>|730,731
freezing|731,739
.|739,740
For|741,744
his|745,748
gait|749,753
freezing|754,762
,|762,763
his|764,767
mirapex|768,775
was|776,779
increased|780,789
by|790,792
<EOL>|792,793
0.125|793,798
mg|799,801
every|802,807
week|808,812
to|813,815
a|816,817
goal|818,822
dose|823,827
of|828,830
0.75|831,835
mg|836,838
t|839,840
.|840,841
i|841,842
.|842,843
d|843,844
.|844,845
He|846,848
<EOL>|848,849
successfully|849,861
up|862,864
-|864,865
titrated|865,873
the|874,877
medicine|878,886
to|887,889
0.75|890,894
/|894,895
0.625|895,900
/|900,901
0.625|901,906
but|907,910
<EOL>|910,911
began|911,916
to|917,919
have|920,924
visual|925,931
hallucinations|932,946
and|947,950
confusion|951,960
so|961,963
on|964,966
_|967,968
_|968,969
_|969,970
his|971,974
<EOL>|974,975
neurologist|975,986
recommended|987,998
decreasing|999,1009
the|1010,1013
dose|1014,1018
to|1019,1021
0.625|1022,1027
TID|1028,1031
.|1031,1032
<EOL>|1033,1034
Despite|1034,1041
<EOL>|1041,1042
the|1042,1045
changes|1046,1053
to|1054,1056
his|1057,1060
Mirapex|1061,1068
,|1068,1069
the|1070,1073
patient|1074,1081
's|1081,1083
daughter|1084,1092
has|1093,1096
noted|1097,1102
<EOL>|1102,1103
progressive|1103,1114
gait|1115,1119
stiffness|1120,1129
and|1130,1133
increased|1134,1143
difficulty|1144,1154
standing|1155,1163
.|1163,1164
<EOL>|1164,1165
This|1165,1169
has|1170,1173
resulted|1174,1182
in|1183,1185
difficulty|1186,1196
with|1197,1201
simply|1202,1208
getting|1209,1216
to|1217,1219
the|1220,1223
<EOL>|1223,1224
bathroom|1224,1232
leading|1233,1240
to|1241,1243
episodes|1244,1252
of|1253,1255
incontinence|1256,1268
.|1268,1269
A|1270,1271
UA|1272,1274
performed|1275,1284
on|1285,1287
<EOL>|1287,1288
_|1288,1289
_|1289,1290
_|1290,1291
was|1292,1295
reassuring|1296,1306
.|1306,1307
<EOL>|1308,1309
<EOL>|1309,1310
On|1310,1312
the|1313,1316
day|1317,1320
of|1321,1323
presentation|1324,1336
to|1337,1339
the|1340,1343
hospital|1344,1352
,|1352,1353
the|1354,1357
patient|1358,1365
began|1366,1371
to|1372,1374
<EOL>|1374,1375
experience|1375,1385
visual|1386,1392
hallucinations|1393,1407
of|1408,1410
a|1411,1412
motor|1413,1418
cross|1419,1424
race|1425,1429
in|1430,1432
his|1433,1436
<EOL>|1436,1437
backyard|1437,1445
.|1445,1446
He|1447,1449
subsequently|1450,1462
had|1463,1466
a|1467,1468
fall|1469,1473
while|1474,1479
transferring|1480,1492
from|1493,1497
the|1498,1501
<EOL>|1501,1502
couch|1502,1507
to|1508,1510
a|1511,1512
chair|1513,1518
.|1518,1519
His|1520,1523
wife|1524,1528
was|1529,1532
unable|1533,1539
to|1540,1542
get|1543,1546
him|1547,1550
off|1551,1554
the|1555,1558
floor|1559,1564
.|1564,1565
<EOL>|1565,1566
The|1566,1569
fall|1570,1574
was|1575,1578
witnessed|1579,1588
and|1589,1592
there|1593,1598
was|1599,1602
no|1603,1605
head|1606,1610
strike|1611,1617
.|1617,1618
Per|1619,1622
the|1623,1626
<EOL>|1626,1627
patient|1627,1634
's|1634,1636
wife|1637,1641
,|1641,1642
his|1643,1646
gait|1647,1651
has|1652,1655
acutely|1656,1663
worsened|1664,1672
over|1673,1677
the|1678,1681
past|1682,1686
24|1687,1689
<EOL>|1689,1690
hours|1690,1695
to|1696,1698
the|1699,1702
point|1703,1708
where|1709,1714
he|1715,1717
has|1718,1721
been|1722,1726
unable|1727,1733
to|1734,1736
ambulate|1737,1745
on|1746,1748
his|1749,1752
<EOL>|1752,1753
own|1753,1756
.|1756,1757
The|1758,1761
patient|1762,1769
's|1769,1771
daughter|1772,1780
called|1781,1787
his|1788,1791
neurologist|1792,1803
who|1804,1807
<EOL>|1807,1808
recommended|1808,1819
presentation|1820,1832
to|1833,1835
the|1836,1839
ED|1840,1842
.|1842,1843
<EOL>|1844,1845
<EOL>|1845,1846
In|1846,1848
the|1849,1852
ED|1853,1855
,|1855,1856
the|1857,1860
patient|1861,1868
was|1869,1872
afebrile|1873,1881
,|1881,1882
HRs|1883,1886
_|1887,1888
_|1888,1889
_|1889,1890
,|1890,1891
normotensive|1892,1904
,|1904,1905
and|1906,1909
<EOL>|1909,1910
SpO2|1910,1914
100|1915,1918
%|1918,1919
RA|1920,1922
.|1922,1923
On|1924,1926
exam|1927,1931
he|1932,1934
was|1935,1938
noted|1939,1944
to|1945,1947
have|1948,1952
cogwheeling|1953,1964
of|1965,1967
upper|1968,1973
<EOL>|1973,1974
extremities|1974,1985
and|1986,1989
decrease|1990,1998
_|1999,2000
_|2000,2001
_|2001,2002
strength|2003,2011
.|2011,2012
Labs|2013,2017
were|2018,2022
remarkable|2023,2033
for|2034,2037
a|2038,2039
<EOL>|2039,2040
negative|2040,2048
urine|2049,2054
and|2055,2058
serum|2059,2064
tox|2065,2068
,|2068,2069
Na|2070,2072
132|2073,2076
,|2076,2077
K|2078,2079
5.8|2080,2083
(|2084,2085
hemolyzed|2085,2094
and|2095,2098
no|2099,2101
<EOL>|2102,2103
EKG|2103,2106
<EOL>|2106,2107
changes|2107,2114
)|2114,2115
,|2115,2116
negative|2117,2125
troponin|2126,2134
,|2134,2135
normal|2136,2142
LFTs|2143,2147
,|2147,2148
unremarkable|2149,2161
CBC|2162,2165
.|2165,2166
<EOL>|2167,2168
Chest|2168,2173
<EOL>|2173,2174
Xray|2174,2178
showed|2179,2185
no|2186,2188
acute|2189,2194
process|2195,2202
and|2203,2206
CTH|2207,2210
was|2211,2214
reassuring|2215,2225
.|2225,2226
He|2227,2229
was|2230,2233
<EOL>|2233,2234
evaluated|2234,2243
by|2244,2246
neurology|2247,2256
who|2257,2260
recommended|2261,2272
admission|2273,2282
to|2283,2285
medicine|2286,2294
for|2295,2298
<EOL>|2298,2299
failure|2299,2306
to|2307,2309
thrive|2310,2316
,|2316,2317
to|2318,2320
continue|2321,2329
the|2330,2333
patient|2334,2341
's|2341,2343
home|2344,2348
medications|2349,2360
,|2360,2361
<EOL>|2361,2362
and|2362,2365
complete|2366,2374
a|2375,2376
toxo|2377,2381
-|2381,2382
metabolic|2382,2391
workup|2392,2398
.|2398,2399
The|2400,2403
patient|2404,2411
was|2412,2415
given|2416,2421
his|2422,2425
<EOL>|2425,2426
home|2426,2430
pramipexole|2431,2442
and|2443,2446
pravastatin|2447,2458
before|2459,2465
he|2466,2468
was|2469,2472
admitted|2473,2481
.|2481,2482
<EOL>|2484,2485
<EOL>|2485,2486
On|2486,2488
arrival|2489,2496
to|2497,2499
the|2500,2503
floor|2504,2509
,|2509,2510
the|2511,2514
patient|2515,2522
is|2523,2525
comfortable|2526,2537
in|2538,2540
bed|2541,2544
.|2544,2545
He|2546,2548
<EOL>|2549,2550
is|2550,2552
<EOL>|2552,2553
not|2553,2556
accompanied|2557,2568
by|2569,2571
family|2572,2578
on|2579,2581
my|2582,2584
interview|2585,2594
.|2594,2595
He|2596,2598
knows|2599,2604
that|2605,2609
he|2610,2612
is|2613,2615
<EOL>|2616,2617
in|2617,2619
<EOL>|2619,2620
the|2620,2623
hospital|2624,2632
and|2633,2636
that|2637,2641
it|2642,2644
is|2645,2647
_|2648,2649
_|2649,2650
_|2650,2651
.|2651,2652
He|2653,2655
is|2656,2658
not|2659,2662
sure|2663,2667
why|2668,2671
he|2672,2674
is|2675,2677
here|2678,2682
<EOL>|2682,2683
and|2683,2686
begins|2687,2693
to|2694,2696
tell|2697,2701
me|2702,2704
about|2705,2710
a|2711,2712
party|2713,2718
in|2719,2721
his|2722,2725
house|2726,2731
with|2732,2736
a|2737,2738
motor|2739,2744
<EOL>|2744,2745
cross|2745,2750
race|2751,2755
in|2756,2758
his|2759,2762
backyard|2763,2771
.|2771,2772
When|2773,2777
I|2778,2779
asked|2780,2785
him|2786,2789
about|2790,2795
his|2796,2799
fall|2800,2804
,|2804,2805
he|2806,2808
<EOL>|2808,2809
mentions|2809,2817
that|2818,2822
he|2823,2825
has|2826,2829
not|2830,2833
had|2834,2837
a|2838,2839
fall|2840,2844
for|2845,2848
_|2849,2850
_|2850,2851
_|2851,2852
years|2853,2858
.|2858,2859
He|2860,2862
denies|2863,2869
any|2870,2873
<EOL>|2873,2874
fevers|2874,2880
,|2880,2881
chills|2882,2888
,|2888,2889
cough|2890,2895
,|2895,2896
chest|2897,2902
pain|2903,2907
,|2907,2908
abdominal|2909,2918
pain|2919,2923
,|2923,2924
nausea|2925,2931
,|2931,2932
<EOL>|2932,2933
diarrhea|2933,2941
,|2941,2942
or|2943,2945
dysuria|2946,2953
.|2953,2954
<EOL>|2955,2956
<EOL>|2956,2957
REVIEW|2957,2963
OF|2964,2966
SYSTEMS|2967,2974
:|2974,2975
<EOL>|2975,2976
=|2976,2977
=|2977,2978
=|2978,2979
=|2979,2980
=|2980,2981
=|2981,2982
=|2982,2983
=|2983,2984
=|2984,2985
=|2985,2986
=|2986,2987
=|2987,2988
=|2988,2989
=|2989,2990
=|2990,2991
=|2991,2992
=|2992,2993
=|2993,2994
<EOL>|2994,2995
Per|2995,2998
HPI|2999,3002
,|3002,3003
otherwise|3004,3013
,|3013,3014
10|3015,3017
-|3017,3018
point|3018,3023
review|3024,3030
of|3031,3033
systems|3034,3041
was|3042,3045
within|3046,3052
normal|3053,3059
<EOL>|3059,3060
limits|3060,3066
.|3066,3067
<EOL>|3067,3068
<EOL>|3068,3069
<EOL>|3070,3071
Past|3071,3075
Medical|3076,3083
History|3084,3091
:|3091,3092
<EOL>|3092,3093
_|3093,3094
_|3094,3095
_|3095,3096
disease|3097,3104
<EOL>|3104,3105
_|3105,3106
_|3106,3107
_|3107,3108
Body|3109,3113
Dementia|3114,3122
<EOL>|3123,3124
dyslipidemia|3124,3136
<EOL>|3137,3138
prostate|3138,3146
cancer|3147,3153
(|3154,3155
s|3155,3156
/|3156,3157
p|3157,3158
prostatectomy|3159,3172
)|3172,3173
<EOL>|3173,3174
<EOL>|3175,3176
Social|3176,3182
History|3183,3190
:|3190,3191
<EOL>|3191,3192
_|3192,3193
_|3193,3194
_|3194,3195
<EOL>|3195,3196
Family|3196,3202
History|3203,3210
:|3210,3211
<EOL>|3211,3212
His|3212,3215
mother|3216,3222
died|3223,3227
at|3228,3230
age|3231,3234
_|3235,3236
_|3236,3237
_|3237,3238
of|3239,3241
"|3242,3243
old|3243,3246
age|3247,3250
.|3250,3251
"|3251,3252
<EOL>|3252,3253
His|3253,3256
father|3257,3263
died|3264,3268
of|3269,3271
prostate|3272,3280
cancer|3281,3287
at|3288,3290
_|3291,3292
_|3292,3293
_|3293,3294
.|3294,3295
He|3297,3299
has|3300,3303
an|3304,3306
older|3307,3312
<EOL>|3313,3314
sister|3314,3320
<EOL>|3320,3321
(|3321,3322
age|3322,3325
_|3326,3327
_|3327,3328
_|3328,3329
and|3330,3333
a|3334,3335
younger|3336,3343
sister|3344,3350
(|3351,3352
age|3352,3355
_|3356,3357
_|3357,3358
_|3358,3359
.|3359,3360
He|3362,3364
has|3365,3368
a|3369,3370
younger|3371,3378
<EOL>|3379,3380
brother|3380,3387
<EOL>|3387,3388
(|3388,3389
age|3389,3392
_|3393,3394
_|3394,3395
_|3395,3396
.|3396,3397
As|3399,3401
noted|3402,3407
,|3407,3408
he|3409,3411
has|3412,3415
2|3416,3417
daughters|3418,3427
.|3427,3428
There|3430,3435
is|3436,3438
no|3439,3441
family|3442,3448
<EOL>|3448,3449
history|3449,3456
of|3457,3459
neurologic|3460,3470
illness|3471,3478
or|3479,3481
dementia|3482,3490
.|3490,3491
There|3493,3498
is|3499,3501
no|3502,3504
family|3505,3511
<EOL>|3511,3512
history|3512,3519
of|3520,3522
neurodevelopmental|3523,3541
mental|3542,3548
disorders|3549,3558
such|3559,3563
as|3564,3566
learning|3567,3575
<EOL>|3575,3576
disability|3576,3586
or|3587,3589
ADHD|3590,3594
.|3594,3595
There|3597,3602
is|3603,3605
no|3606,3608
family|3609,3615
history|3616,3623
of|3624,3626
psychiatric|3627,3638
<EOL>|3638,3639
problems|3639,3647
.|3647,3648
<EOL>|3648,3649
<EOL>|3650,3651
Physical|3651,3659
Exam|3660,3664
:|3664,3665
<EOL>|3665,3666
ADMISSION|3666,3675
PHYSICAL|3676,3684
EXAM|3685,3689
:|3689,3690
<EOL>|3690,3691
=|3691,3692
=|3692,3693
=|3693,3694
=|3694,3695
=|3695,3696
=|3696,3697
=|3697,3698
=|3698,3699
=|3699,3700
=|3700,3701
=|3701,3702
=|3702,3703
=|3703,3704
=|3704,3705
=|3705,3706
=|3706,3707
=|3707,3708
=|3708,3709
=|3709,3710
=|3710,3711
=|3711,3712
=|3712,3713
=|3713,3714
=|3714,3715
<EOL>|3715,3716
VITALS|3716,3722
:|3722,3723
reviewed|3724,3732
in|3733,3735
OMR|3736,3739
<EOL>|3740,3741
GENERAL|3741,3748
:|3748,3749
Alert|3750,3755
and|3756,3759
interactive|3760,3771
.|3771,3772
In|3773,3775
no|3776,3778
acute|3779,3784
distress|3785,3793
.|3793,3794
<EOL>|3794,3795
HEENT|3795,3800
:|3800,3801
PERRL|3802,3807
,|3807,3808
EOMI|3809,3813
.|3813,3814
Sclera|3815,3821
anicteric|3822,3831
and|3832,3835
without|3836,3843
injection|3844,3853
.|3853,3854
MMM|3855,3858
.|3858,3859
<EOL>|3859,3860
NECK|3860,3864
:|3864,3865
No|3866,3868
cervical|3869,3877
lymphadenopathy|3878,3893
.|3893,3894
No|3895,3897
JVD|3898,3901
.|3901,3902
<EOL>|3902,3903
CARDIAC|3903,3910
:|3910,3911
Regular|3912,3919
rhythm|3920,3926
,|3926,3927
normal|3928,3934
rate|3935,3939
.|3939,3940
Audible|3941,3948
S1|3949,3951
and|3952,3955
S2|3956,3958
.|3958,3959
No|3960,3962
<EOL>|3962,3963
murmurs|3963,3970
/|3970,3971
rubs|3971,3975
/|3975,3976
gallops|3976,3983
.|3983,3984
<EOL>|3984,3985
LUNGS|3985,3990
:|3990,3991
Clear|3992,3997
to|3998,4000
auscultation|4001,4013
bilaterally|4014,4025
.|4025,4026
No|4027,4029
wheezes|4030,4037
,|4037,4038
rhonchi|4039,4046
or|4047,4049
<EOL>|4049,4050
rales|4050,4055
.|4055,4056
No|4057,4059
increased|4060,4069
work|4070,4074
of|4075,4077
breathing|4078,4087
.|4087,4088
<EOL>|4088,4089
BACK|4089,4093
:|4093,4094
No|4095,4097
CVA|4098,4101
tenderness|4102,4112
.|4112,4113
<EOL>|4113,4114
ABDOMEN|4114,4121
:|4121,4122
Normal|4123,4129
bowels|4130,4136
sounds|4137,4143
,|4143,4144
non|4145,4148
distended|4149,4158
,|4158,4159
non-tender|4160,4170
to|4171,4173
deep|4174,4178
<EOL>|4178,4179
palpation|4179,4188
in|4189,4191
all|4192,4195
four|4196,4200
quadrants|4201,4210
.|4210,4211
No|4212,4214
organomegaly|4215,4227
.|4227,4228
<EOL>|4228,4229
EXTREMITIES|4229,4240
:|4240,4241
No|4242,4244
clubbing|4245,4253
,|4253,4254
cyanosis|4255,4263
,|4263,4264
or|4265,4267
edema|4268,4273
.|4273,4274
Pulses|4275,4281
DP|4282,4284
/|4284,4285
Radial|4285,4291
<EOL>|4292,4293
2|4293,4294
+|4294,4295
<EOL>|4295,4296
bilaterally|4296,4307
.|4307,4308
<EOL>|4308,4309
SKIN|4309,4313
:|4313,4314
Warm|4315,4319
.|4319,4320
Cap|4321,4324
refill|4325,4331
<|4332,4333
2s|4333,4335
.|4335,4336
No|4337,4339
rashes|4340,4346
.|4346,4347
<EOL>|4347,4348
NEUROLOGIC|4348,4358
:|4358,4359
AOx3|4360,4364
.|4364,4365
CN2|4366,4369
-|4369,4370
12|4370,4372
intact|4373,4379
.|4379,4380
cogwheel|4381,4389
UE|4390,4392
b|4393,4394
/|4394,4395
l|4395,4396
.|4396,4397
Increased|4398,4407
tone|4408,4412
<EOL>|4412,4413
in|4413,4415
LEs|4416,4419
,|4419,4420
_|4421,4422
_|4422,4423
_|4423,4424
strength|4425,4433
b|4434,4435
/|4435,4436
l|4436,4437
_|4438,4439
_|4439,4440
_|4440,4441
.|4441,4442
Normal|4443,4449
sensation|4450,4459
.|4459,4460
<EOL>|4460,4461
<EOL>|4461,4462
DISCHARGE|4462,4471
PHYSICAL|4472,4480
EXAM|4481,4485
<EOL>|4485,4486
=|4486,4487
=|4487,4488
=|4488,4489
=|4489,4490
=|4490,4491
=|4491,4492
=|4492,4493
=|4493,4494
=|4494,4495
=|4495,4496
=|4496,4497
=|4497,4498
=|4498,4499
=|4499,4500
=|4500,4501
=|4501,4502
=|4502,4503
=|4503,4504
=|4504,4505
=|4505,4506
=|4506,4507
=|4507,4508
<EOL>|4508,4509
24|4509,4511
HR|4512,4514
Data|4515,4519
(|4520,4521
last|4521,4525
updated|4526,4533
_|4534,4535
_|4535,4536
_|4536,4537
@|4538,4539
2340|4540,4544
)|4544,4545
<EOL>|4545,4546
Temp|4550,4554
:|4554,4555
97.7|4556,4560
(|4561,4562
Tm|4562,4564
98.4|4565,4569
)|4569,4570
,|4570,4571
BP|4572,4574
:|4574,4575
130|4576,4579
/|4579,4580
80|4580,4582
(|4583,4584
130|4584,4587
-|4587,4588
153|4588,4591
/|4591,4592
80|4592,4594
-|4594,4595
90|4595,4597
)|4597,4598
,|4598,4599
HR|4600,4602
:|4602,4603
80|4604,4606
<EOL>|4606,4607
(|4607,4608
80|4608,4610
-|4610,4611
104|4611,4614
)|4614,4615
,|4615,4616
RR|4617,4619
:|4619,4620
18|4621,4623
(|4624,4625
_|4625,4626
_|4626,4627
_|4627,4628
)|4628,4629
,|4629,4630
O2|4631,4633
sat|4634,4637
:|4637,4638
100|4639,4642
%|4642,4643
(|4644,4645
95|4645,4647
-|4647,4648
100|4648,4651
)|4651,4652
,|4652,4653
O2|4654,4656
delivery|4657,4665
:|4665,4666
Ra|4667,4669
<EOL>|4670,4671
<EOL>|4671,4672
<EOL>|4672,4673
GENERAL|4673,4680
:|4680,4681
In|4682,4684
no|4685,4687
acute|4688,4693
distress|4694,4702
.|4702,4703
Talking|4704,4711
very|4712,4716
quietly|4717,4724
.|4724,4725
<EOL>|4725,4726
CARDIAC|4726,4733
:|4733,4734
Regular|4735,4742
rhythm|4743,4749
,|4749,4750
normal|4751,4757
rate|4758,4762
.|4762,4763
Audible|4764,4771
S1|4772,4774
and|4775,4778
S2|4779,4781
.|4781,4782
No|4783,4785
<EOL>|4785,4786
murmurs|4786,4793
/|4793,4794
rubs|4794,4798
/|4798,4799
gallops|4799,4806
.|4806,4807
<EOL>|4807,4808
LUNGS|4808,4813
:|4813,4814
Clear|4815,4820
to|4821,4823
auscultation|4824,4836
bilaterally|4837,4848
.|4848,4849
No|4850,4852
wheezes|4853,4860
,|4860,4861
rhonchi|4862,4869
or|4870,4872
<EOL>|4872,4873
rales|4873,4878
.|4878,4879
No|4880,4882
increased|4883,4892
work|4893,4897
of|4898,4900
breathing|4901,4910
.|4910,4911
<EOL>|4911,4912
ABDOMEN|4912,4919
:|4919,4920
Normal|4921,4927
bowels|4928,4934
sounds|4935,4941
,|4941,4942
non|4943,4946
distended|4947,4956
,|4956,4957
non-tender|4958,4968
to|4969,4971
deep|4972,4976
<EOL>|4976,4977
palpation|4977,4986
in|4987,4989
all|4990,4993
four|4994,4998
quadrants|4999,5008
.|5008,5009
<EOL>|5009,5010
EXTREMITIES|5010,5021
:|5021,5022
No|5023,5025
clubbing|5026,5034
,|5034,5035
cyanosis|5036,5044
,|5044,5045
or|5046,5048
edema|5049,5054
.|5054,5055
Pulses|5056,5062
DP|5063,5065
/|5065,5066
Radial|5066,5072
<EOL>|5073,5074
2|5074,5075
+|5075,5076
<EOL>|5076,5077
bilaterally|5077,5088
.|5088,5089
<EOL>|5089,5090
SKIN|5090,5094
:|5094,5095
Warm|5096,5100
.|5100,5101
<EOL>|5101,5102
NEUROLOGIC|5102,5112
:|5112,5113
AOx3|5114,5118
.|5118,5119
CN2|5120,5123
-|5123,5124
12|5124,5126
intact|5127,5133
.|5133,5134
cogwheel|5135,5143
UE|5144,5146
b|5147,5148
/|5148,5149
l|5149,5150
.|5150,5151
Increased|5152,5161
tone|5162,5166
<EOL>|5166,5167
in|5167,5169
LEs|5170,5173
,|5173,5174
_|5175,5176
_|5176,5177
_|5177,5178
strength|5179,5187
b|5188,5189
/|5189,5190
l|5190,5191
_|5192,5193
_|5193,5194
_|5194,5195
.|5195,5196
Normal|5197,5203
sensation|5204,5213
.|5213,5214
<EOL>|5214,5215
<EOL>|5215,5216
<EOL>|5217,5218
Pertinent|5218,5227
Results|5228,5235
:|5235,5236
<EOL>|5236,5237
ADMISSION|5237,5246
LABS|5247,5251
:|5251,5252
<EOL>|5252,5253
=|5253,5254
=|5254,5255
=|5255,5256
=|5256,5257
=|5257,5258
=|5258,5259
=|5259,5260
=|5260,5261
=|5261,5262
=|5262,5263
=|5263,5264
=|5264,5265
=|5265,5266
=|5266,5267
=|5267,5268
<EOL>|5268,5269
_|5269,5270
_|5270,5271
_|5271,5272
10|5273,5275
:|5275,5276
30PM|5276,5280
BLOOD|5281,5286
WBC|5287,5290
-|5290,5291
8.6|5291,5294
RBC|5295,5298
-|5298,5299
4|5299,5300
.|5300,5301
03|5301,5303
*|5303,5304
Hgb|5305,5308
-|5308,5309
12|5309,5311
.|5311,5312
8|5312,5313
*|5313,5314
Hct|5315,5318
-|5318,5319
38|5319,5321
.|5321,5322
2|5322,5323
*|5323,5324
<EOL>|5325,5326
MCV|5326,5329
-|5329,5330
95|5330,5332
MCH|5333,5336
-|5336,5337
31.8|5337,5341
MCHC|5342,5346
-|5346,5347
33.5|5347,5351
RDW|5352,5355
-|5355,5356
13.0|5356,5360
RDWSD|5361,5366
-|5366,5367
45.2|5367,5371
Plt|5372,5375
_|5376,5377
_|5377,5378
_|5378,5379
<EOL>|5379,5380
_|5380,5381
_|5381,5382
_|5382,5383
10|5384,5386
:|5386,5387
30PM|5387,5391
BLOOD|5392,5397
Neuts|5398,5403
-|5403,5404
48.1|5404,5408
_|5409,5410
_|5410,5411
_|5411,5412
Monos|5413,5418
-|5418,5419
15|5419,5421
.|5421,5422
9|5422,5423
*|5423,5424
<EOL>|5425,5426
Eos|5426,5429
-|5429,5430
2.0|5430,5433
Baso|5434,5438
-|5438,5439
0.6|5439,5442
Im|5443,5445
_|5446,5447
_|5447,5448
_|5448,5449
AbsNeut|5450,5457
-|5457,5458
4|5458,5459
.|5459,5460
13|5460,5462
AbsLymp|5463,5470
-|5470,5471
2|5471,5472
.|5472,5473
86|5473,5475
<EOL>|5476,5477
AbsMono|5477,5484
-|5484,5485
1|5485,5486
.|5486,5487
36|5487,5489
*|5489,5490
AbsEos|5491,5497
-|5497,5498
0|5498,5499
.|5499,5500
17|5500,5502
AbsBaso|5503,5510
-|5510,5511
0|5511,5512
.|5512,5513
05|5513,5515
<EOL>|5515,5516
_|5516,5517
_|5517,5518
_|5518,5519
10|5520,5522
:|5522,5523
30PM|5523,5527
BLOOD|5528,5533
_|5534,5535
_|5535,5536
_|5536,5537
PTT|5538,5541
-|5541,5542
23|5542,5544
.|5544,5545
4|5545,5546
*|5546,5547
_|5548,5549
_|5549,5550
_|5550,5551
<EOL>|5551,5552
_|5552,5553
_|5553,5554
_|5554,5555
10|5556,5558
:|5558,5559
30PM|5559,5563
BLOOD|5564,5569
Glucose|5570,5577
-|5577,5578
100|5578,5581
UreaN|5582,5587
-|5587,5588
17|5588,5590
Creat|5591,5596
-|5596,5597
0.8|5597,5600
Na|5601,5603
-|5603,5604
132|5604,5607
*|5607,5608
<EOL>|5609,5610
K|5610,5611
-|5611,5612
5|5612,5613
.|5613,5614
8|5614,5615
*|5615,5616
Cl|5617,5619
-|5619,5620
98|5620,5622
HCO3|5623,5627
-|5627,5628
19|5628,5630
*|5630,5631
AnGap|5632,5637
-|5637,5638
15|5638,5640
<EOL>|5640,5641
_|5641,5642
_|5642,5643
_|5643,5644
10|5645,5647
:|5647,5648
30PM|5648,5652
BLOOD|5653,5658
ALT|5659,5662
-|5662,5663
18|5663,5665
AST|5666,5669
-|5669,5670
38|5670,5672
AlkPhos|5673,5680
-|5680,5681
39|5681,5683
*|5683,5684
TotBili|5685,5692
-|5692,5693
0.4|5693,5696
<EOL>|5696,5697
_|5697,5698
_|5698,5699
_|5699,5700
10|5701,5703
:|5703,5704
30PM|5704,5708
BLOOD|5709,5714
Lipase|5715,5721
-|5721,5722
47|5722,5724
<EOL>|5724,5725
_|5725,5726
_|5726,5727
_|5727,5728
10|5729,5731
:|5731,5732
30PM|5732,5736
BLOOD|5737,5742
cTropnT|5743,5750
-|5750,5751
<|5751,5752
0|5752,5753
.|5753,5754
01|5754,5756
<EOL>|5756,5757
_|5757,5758
_|5758,5759
_|5759,5760
10|5761,5763
:|5763,5764
30PM|5764,5768
BLOOD|5769,5774
Albumin|5775,5782
-|5782,5783
4.0|5783,5786
Calcium|5787,5794
-|5794,5795
9.9|5795,5798
Phos|5799,5803
-|5803,5804
3.7|5804,5807
Mg|5808,5810
-|5810,5811
2.0|5811,5814
<EOL>|5814,5815
_|5815,5816
_|5816,5817
_|5817,5818
10|5819,5821
:|5821,5822
30PM|5822,5826
BLOOD|5827,5832
VitB12|5833,5839
-|5839,5840
570|5840,5843
<EOL>|5843,5844
_|5844,5845
_|5845,5846
_|5846,5847
10|5848,5850
:|5850,5851
30PM|5851,5855
BLOOD|5856,5861
TSH|5862,5865
-|5865,5866
1.4|5866,5869
<EOL>|5869,5870
_|5870,5871
_|5871,5872
_|5872,5873
07|5874,5876
:|5876,5877
00AM|5877,5881
BLOOD|5882,5887
Trep|5888,5892
Ab|5893,5895
-|5895,5896
NEG|5896,5899
<EOL>|5899,5900
_|5900,5901
_|5901,5902
_|5902,5903
10|5904,5906
:|5906,5907
30PM|5907,5911
BLOOD|5912,5917
ASA|5918,5921
-|5921,5922
NEG|5922,5925
Ethanol|5926,5933
-|5933,5934
NEG|5934,5937
Acetmnp|5938,5945
-|5945,5946
NEG|5946,5949
<EOL>|5950,5951
Tricycl|5951,5958
-|5958,5959
NEG|5959,5962
<EOL>|5962,5963
<EOL>|5963,5964
IMAGING|5964,5971
:|5971,5972
<EOL>|5972,5973
=|5973,5974
=|5974,5975
=|5975,5976
=|5976,5977
=|5977,5978
=|5978,5979
=|5979,5980
=|5980,5981
<EOL>|5981,5982
_|5982,5983
_|5983,5984
_|5984,5985
Imaging|5986,5993
CT|5994,5996
HEAD|5997,6001
W|6002,6003
/|6003,6004
O|6004,6005
CONTRAST|6006,6014
<EOL>|6016,6017
FINDINGS|6017,6025
:|6025,6026
<EOL>|6028,6029
There|6029,6034
is|6035,6037
no|6038,6040
evidence|6041,6049
of|6050,6052
infarction|6053,6063
,|6063,6064
hemorrhage|6065,6075
,|6075,6076
edema|6077,6082
,|6082,6083
or|6084,6086
mass|6087,6091
.|6091,6092
<EOL>|6094,6095
There|6095,6100
is|6101,6103
<EOL>|6104,6105
prominence|6105,6115
of|6116,6118
the|6119,6122
ventricles|6123,6133
and|6134,6137
sulci|6138,6143
suggestive|6144,6154
of|6155,6157
<EOL>|6158,6159
involutional|6159,6171
changes|6172,6179
.|6179,6180
<EOL>|6181,6182
There|6182,6187
is|6188,6190
no|6191,6193
evidence|6194,6202
of|6203,6205
fracture|6206,6214
.|6214,6215
The|6217,6220
visualized|6221,6231
portion|6232,6239
of|6240,6242
the|6243,6246
<EOL>|6247,6248
remaining|6248,6257
<EOL>|6258,6259
paranasal|6259,6268
sinuses|6269,6276
and|6277,6280
middle|6281,6287
ear|6288,6291
cavities|6292,6300
are|6301,6304
clear|6305,6310
.|6310,6311
The|6313,6316
<EOL>|6317,6318
visualized|6318,6328
portion|6329,6336
of|6337,6339
the|6340,6343
orbits|6344,6350
are|6351,6354
unremarkable|6355,6367
apart|6368,6373
from|6374,6378
<EOL>|6379,6380
bilateral|6380,6389
lens|6390,6394
replacements|6395,6407
.|6407,6408
<EOL>|6409,6410
IMPRESSION|6410,6420
:|6420,6421
<EOL>|6422,6423
1|6423,6424
.|6424,6425
No|6426,6428
acute|6429,6434
intracranial|6435,6447
abnormality|6448,6459
.|6459,6460
No|6462,6464
hydrocephalus|6465,6478
.|6478,6479
<EOL>|6480,6481
<EOL>|6481,6482
_|6482,6483
_|6483,6484
_|6484,6485
Imaging|6486,6493
CHEST|6494,6499
(|6500,6501
PA|6501,6503
&|6504,6505
LAT|6506,6509
)|6509,6510
<EOL>|6511,6512
IMPRESSION|6512,6522
:|6522,6523
<EOL>|6525,6526
Mild|6526,6530
atelectasis|6531,6542
in|6543,6545
the|6546,6549
lung|6550,6554
bases|6555,6560
without|6561,6568
focal|6569,6574
consolidation|6575,6588
.|6588,6589
<EOL>|6591,6592
<EOL>|6592,6593
Age|6593,6596
-|6596,6597
indeterminate|6597,6610
moderate|6611,6619
to|6620,6622
severe|6623,6629
compression|6630,6641
deformity|6642,6651
of|6652,6654
a|6655,6656
<EOL>|6657,6658
low|6658,6661
thoracic|6662,6670
vertebral|6671,6680
body|6681,6685
.|6685,6686
<EOL>|6687,6688
<EOL>|6688,6689
DISCHARGE|6689,6698
LABS|6699,6703
:|6703,6704
<EOL>|6704,6705
=|6705,6706
=|6706,6707
=|6707,6708
=|6708,6709
=|6709,6710
=|6710,6711
=|6711,6712
=|6712,6713
=|6713,6714
=|6714,6715
=|6715,6716
=|6716,6717
=|6717,6718
=|6718,6719
=|6719,6720
<EOL>|6720,6721
_|6721,6722
_|6722,6723
_|6723,6724
06|6725,6727
:|6727,6728
21AM|6728,6732
BLOOD|6733,6738
WBC|6739,6742
-|6742,6743
7.0|6743,6746
RBC|6747,6750
-|6750,6751
4|6751,6752
.|6752,6753
02|6753,6755
*|6755,6756
Hgb|6757,6760
-|6760,6761
12|6761,6763
.|6763,6764
9|6764,6765
*|6765,6766
Hct|6767,6770
-|6770,6771
38|6771,6773
.|6773,6774
1|6774,6775
*|6775,6776
<EOL>|6777,6778
MCV|6778,6781
-|6781,6782
95|6782,6784
MCH|6785,6788
-|6788,6789
32|6789,6791
.|6791,6792
1|6792,6793
*|6793,6794
MCHC|6795,6799
-|6799,6800
33.9|6800,6804
RDW|6805,6808
-|6808,6809
12.8|6809,6813
RDWSD|6814,6819
-|6819,6820
44.4|6820,6824
Plt|6825,6828
_|6829,6830
_|6830,6831
_|6831,6832
<EOL>|6832,6833
_|6833,6834
_|6834,6835
_|6835,6836
06|6837,6839
:|6839,6840
21AM|6840,6844
BLOOD|6845,6850
Glucose|6851,6858
-|6858,6859
88|6859,6861
UreaN|6862,6867
-|6867,6868
10|6868,6870
Creat|6871,6876
-|6876,6877
0.7|6877,6880
Na|6881,6883
-|6883,6884
140|6884,6887
<EOL>|6888,6889
K|6889,6890
-|6890,6891
4.0|6891,6894
Cl|6895,6897
-|6897,6898
104|6898,6901
HCO3|6902,6906
-|6906,6907
24|6907,6909
AnGap|6910,6915
-|6915,6916
12|6916,6918
<EOL>|6918,6919
_|6919,6920
_|6920,6921
_|6921,6922
06|6923,6925
:|6925,6926
21AM|6926,6930
BLOOD|6931,6936
Calcium|6937,6944
-|6944,6945
9.5|6945,6948
Phos|6949,6953
-|6953,6954
3.2|6954,6957
Mg|6958,6960
-|6960,6961
1.|6961,6963
_|6963,6964
_|6964,6965
_|6965,6966
male|6967,6971
with|6972,6976
_|6977,6978
_|6978,6979
_|6979,6980
disease|6981,6988
,|6988,6989
dyslipidemia|6990,7002
,|7002,7003
and|7004,7007
a|7008,7009
<EOL>|7009,7010
history|7010,7017
of|7018,7020
prostate|7021,7029
cancer|7030,7036
(|7037,7038
s|7038,7039
/|7039,7040
p|7040,7041
prostatectomy|7042,7055
)|7055,7056
who|7057,7060
was|7061,7064
referred|7065,7073
<EOL>|7073,7074
to|7074,7076
the|7077,7080
ED|7081,7083
by|7084,7086
his|7087,7090
neurologist|7091,7102
for|7103,7106
worsening|7107,7116
gait|7117,7121
,|7121,7122
falls|7123,7128
,|7128,7129
and|7130,7133
<EOL>|7133,7134
visual|7134,7140
hallucinations|7141,7155
concerning|7156,7166
for|7167,7170
progression|7171,7182
of|7183,7185
his|7186,7189
<EOL>|7189,7190
neurologic|7190,7200
disorder|7201,7209
.|7209,7210
<EOL>|7211,7212
<EOL>|7212,7213
ACUTE|7213,7218
/|7218,7219
ACTIVE|7219,7225
ISSUES|7226,7232
:|7232,7233
<EOL>|7233,7234
=|7234,7235
=|7235,7236
=|7236,7237
=|7237,7238
=|7238,7239
=|7239,7240
=|7240,7241
=|7241,7242
=|7242,7243
=|7243,7244
=|7244,7245
=|7245,7246
=|7246,7247
=|7247,7248
=|7248,7249
=|7249,7250
=|7250,7251
=|7251,7252
=|7252,7253
=|7253,7254
<EOL>|7254,7255
_|7255,7256
_|7256,7257
_|7257,7258
disease|7259,7266
<EOL>|7266,7267
_|7267,7268
_|7268,7269
_|7269,7270
Body|7271,7275
Dementia|7276,7284
<EOL>|7285,7286
#|7286,7287
Visual|7287,7293
Hallucinations|7294,7308
<EOL>|7309,7310
The|7310,7313
patient|7314,7321
appears|7322,7329
to|7330,7332
have|7333,7337
acute|7338,7343
on|7344,7346
chronic|7347,7354
progression|7355,7366
of|7367,7369
his|7370,7373
<EOL>|7373,7374
_|7374,7375
_|7375,7376
_|7376,7377
disease|7378,7385
.|7385,7386
Unclear|7387,7394
if|7395,7397
this|7398,7402
is|7403,7405
disease|7406,7413
progression|7414,7425
or|7426,7428
<EOL>|7428,7429
underlying|7429,7439
medical|7440,7447
cause|7448,7453
.|7453,7454
Continued|7455,7464
mirapex|7465,7472
,|7472,7473
rasagiline|7474,7484
,|7484,7485
and|7486,7489
<EOL>|7490,7491
rivastigmine|7491,7503
.|7503,7504
Neurology|7505,7514
recommended|7515,7526
started|7527,7534
Seroquel|7535,7543
for|7544,7547
his|7548,7551
<EOL>|7552,7553
hallucinations|7553,7567
.|7567,7568
<EOL>|7568,7569
<EOL>|7569,7570
He|7570,7572
was|7573,7576
evaluated|7577,7586
by|7587,7589
physical|7590,7598
therapy|7599,7606
who|7607,7610
recommended|7611,7622
rehab|7623,7628
.|7628,7629
This|7630,7634
<EOL>|7635,7636
recommendation|7636,7650
was|7651,7654
discussed|7655,7664
with|7665,7669
the|7670,7673
family|7674,7680
who|7681,7684
opted|7685,7690
for|7691,7694
<EOL>|7695,7696
discharge|7696,7705
to|7706,7708
home|7709,7713
with|7714,7718
home|7719,7723
physical|7724,7732
therapy|7733,7740
as|7741,7743
this|7744,7748
was|7749,7752
in|7753,7755
line|7756,7760
<EOL>|7761,7762
with|7762,7766
the|7767,7770
patient|7771,7778
's|7778,7780
goals|7781,7786
of|7787,7789
care|7790,7794
.|7794,7795
<EOL>|7795,7796
<EOL>|7796,7797
TRANSITIONAL|7797,7809
ISSUES|7810,7816
:|7816,7817
<EOL>|7817,7818
[|7818,7819
]|7819,7820
f|7821,7822
/|7822,7823
u|7823,7824
visual|7825,7831
hallucination|7832,7845
symptoms|7846,7854
on|7855,7857
Seroquel|7858,7866
<EOL>|7866,7867
[|7867,7868
]|7868,7869
f|7870,7871
/|7871,7872
u|7872,7873
physical|7874,7882
therapy|7883,7890
at|7891,7893
home|7894,7898
<EOL>|7898,7899
<EOL>|7900,7901
Medications|7901,7912
on|7913,7915
Admission|7916,7925
:|7925,7926
<EOL>|7926,7927
The|7927,7930
Preadmission|7931,7943
Medication|7944,7954
list|7955,7959
may|7960,7963
be|7964,7966
inaccurate|7967,7977
and|7978,7981
requires|7982,7990
<EOL>|7991,7992
futher|7992,7998
investigation|7999,8012
.|8012,8013
<EOL>|8013,8014
1.|8014,8016
Rasagiline|8017,8027
1|8028,8029
mg|8030,8032
PO|8033,8035
DAILY|8036,8041
<EOL>|8042,8043
2.|8043,8045
Pramipexole|8046,8057
0.625|8058,8063
mg|8064,8066
PO|8067,8069
TID|8070,8073
<EOL>|8074,8075
3.|8075,8077
rivastigmine|8078,8090
9.5|8091,8094
mg|8095,8097
/|8097,8098
24|8098,8100
hr|8101,8103
transdermal|8104,8115
DAILY|8116,8121
<EOL>|8122,8123
4.|8123,8125
Pravastatin|8126,8137
40|8138,8140
mg|8141,8143
PO|8144,8146
QPM|8147,8150
<EOL>|8151,8152
5.|8152,8154
Cyanocobalamin|8155,8169
Dose|8170,8174
is|8175,8177
Unknown|8178,8185
PO|8187,8189
DAILY|8190,8195
<EOL>|8196,8197
6.|8197,8199
Loratadine|8200,8210
10|8211,8213
mg|8214,8216
PO|8217,8219
DAILY|8220,8225
<EOL>|8226,8227
<EOL>|8227,8228
<EOL>|8229,8230
Discharge|8230,8239
Medications|8240,8251
:|8251,8252
<EOL>|8252,8253
1.|8253,8255
QUEtiapine|8257,8267
Fumarate|8268,8276
25|8277,8279
mg|8280,8282
PO|8283,8285
QHS|8286,8289
<EOL>|8290,8291
RX|8291,8293
*|8294,8295
quetiapine|8295,8305
25|8306,8308
mg|8309,8311
1|8312,8313
tablet|8314,8320
(|8320,8321
s|8321,8322
)|8322,8323
by|8324,8326
mouth|8327,8332
AT|8333,8335
NIGHT|8336,8341
Disp|8342,8346
#|8347,8348
*|8348,8349
30|8349,8351
<EOL>|8352,8353
Tablet|8353,8359
Refills|8360,8367
:|8367,8368
*|8368,8369
0|8369,8370
<EOL>|8371,8372
2.|8372,8374
Loratadine|8376,8386
10|8387,8389
mg|8390,8392
PO|8393,8395
DAILY|8396,8401
<EOL>|8403,8404
3.|8404,8406
Pramipexole|8408,8419
0.625|8420,8425
mg|8426,8428
PO|8429,8431
TID|8432,8435
<EOL>|8437,8438
4.|8438,8440
Pravastatin|8442,8453
40|8454,8456
mg|8457,8459
PO|8460,8462
QPM|8463,8466
<EOL>|8468,8469
5.|8469,8471
Rasagiline|8473,8483
1|8484,8485
mg|8486,8488
PO|8489,8491
DAILY|8492,8497
<EOL>|8499,8500
6.|8500,8502
rivastigmine|8504,8516
9.5|8517,8520
mg|8521,8523
/|8523,8524
24|8524,8526
hr|8527,8529
transdermal|8530,8541
DAILY|8542,8547
<EOL>|8549,8550
<EOL>|8550,8551
<EOL>|8552,8553
Discharge|8553,8562
Disposition|8563,8574
:|8574,8575
<EOL>|8575,8576
Home|8576,8580
With|8581,8585
Service|8586,8593
<EOL>|8593,8594
<EOL>|8595,8596
Facility|8596,8604
:|8604,8605
<EOL>|8605,8606
_|8606,8607
_|8607,8608
_|8608,8609
<EOL>|8609,8610
<EOL>|8611,8612
Discharge|8612,8621
Diagnosis|8622,8631
:|8631,8632
<EOL>|8632,8633
_|8633,8634
_|8634,8635
_|8635,8636
Dementia|8637,8645
<EOL>|8645,8646
<EOL>|8647,8648
Discharge|8648,8657
Condition|8658,8667
:|8667,8668
<EOL>|8668,8669
Mental|8669,8675
Status|8676,8682
:|8682,8683
Confused|8684,8692
-|8693,8694
sometimes|8695,8704
.|8704,8705
<EOL>|8705,8706
Level|8706,8711
of|8712,8714
Consciousness|8715,8728
:|8728,8729
Alert|8730,8735
and|8736,8739
interactive|8740,8751
.|8751,8752
<EOL>|8752,8753
<EOL>|8753,8754
<EOL>|8755,8756
Discharge|8756,8765
Instructions|8766,8778
:|8778,8779
<EOL>|8779,8780
Dear|8780,8784
Mr.|8785,8788
_|8789,8790
_|8790,8791
_|8791,8792
,|8792,8793
<EOL>|8794,8795
<EOL>|8795,8796
It|8796,8798
was|8799,8802
a|8803,8804
privilege|8805,8814
caring|8815,8821
for|8822,8825
you|8826,8829
at|8830,8832
_|8833,8834
_|8834,8835
_|8835,8836
.|8836,8837
<EOL>|8838,8839
<EOL>|8839,8840
WHY|8840,8843
WAS|8844,8847
I|8848,8849
IN|8850,8852
THE|8853,8856
HOSPITAL|8857,8865
?|8865,8866
<EOL>|8867,8868
-|8868,8869
You|8870,8873
were|8874,8878
sent|8879,8883
to|8884,8886
the|8887,8890
emergency|8891,8900
room|8901,8905
by|8906,8908
your|8909,8913
neurologist|8914,8925
who|8926,8929
<EOL>|8930,8931
was|8931,8934
concerned|8935,8944
that|8945,8949
you|8950,8953
were|8954,8958
having|8959,8965
visual|8966,8972
hallucinations|8973,8987
.|8987,8988
<EOL>|8988,8989
<EOL>|8989,8990
WHAT|8990,8994
HAPPENED|8995,9003
TO|9004,9006
ME|9007,9009
IN|9010,9012
THE|9013,9016
HOSPITAL|9017,9025
?|9025,9026
<EOL>|9027,9028
-|9028,9029
You|9030,9033
were|9034,9038
started|9039,9046
on|9047,9049
a|9050,9051
new|9052,9055
medication|9056,9066
to|9067,9069
help|9070,9074
treat|9075,9080
your|9081,9085
<EOL>|9086,9087
symptoms|9087,9095
.|9095,9096
<EOL>|9096,9097
<EOL>|9097,9098
WHAT|9098,9102
SHOULD|9103,9109
I|9110,9111
DO|9112,9114
AFTER|9115,9120
I|9121,9122
LEAVE|9123,9128
THE|9129,9132
HOSPITAL|9133,9141
?|9141,9142
<EOL>|9143,9144
-|9144,9145
Continue|9146,9154
to|9155,9157
take|9158,9162
all|9163,9166
your|9167,9171
medicines|9172,9181
and|9182,9185
keep|9186,9190
your|9191,9195
<EOL>|9196,9197
appointments|9197,9209
.|9209,9210
<EOL>|9211,9212
<EOL>|9212,9213
We|9213,9215
wish|9216,9220
you|9221,9224
the|9225,9228
best|9229,9233
!|9233,9234
<EOL>|9235,9236
<EOL>|9236,9237
Sincerely|9237,9246
,|9246,9247
<EOL>|9248,9249
Your|9249,9253
_|9254,9255
_|9255,9256
_|9256,9257
Team|9258,9262
<EOL>|9263,9264
<EOL>|9265,9266
Followup|9266,9274
Instructions|9275,9287
:|9287,9288
<EOL>|9288,9289
_|9289,9290
_|9290,9291
_|9291,9292
<EOL>|9292,9293

