CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|true|false||Unit
null|Unit device|Device|true|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|true|false||Unit
null|Unit of Measure|LabModifier|true|false||Unit
null|Unit|LabModifier|true|false||Unit
null|Enzyme Unit|LabModifier|true|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Level of Care - Surgery|Finding|false|false||SURGERY
null|Surgical procedure finding|Finding|false|false||SURGERY
null|Surgical aspects|Finding|false|false||SURGERYnull|Operative Surgical Procedures|Procedure|false|false||SURGERYnull|General surgery specialty|Title|false|false||SURGERY
null|Surgery specialty|Title|false|false||SURGERYnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|codeine|Drug|false|false||Codeine
null|codeine|Drug|false|false||Codeinenull|Augmentin|Drug|false|false||Augmentin
null|Augmentin|Drug|false|false||Augmentinnull|Topamax|Drug|false|false||Topamax
null|Topamax|Drug|false|false||Topamaxnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Complaint (finding)|Finding|false|false||Complaintnull|null|Attribute|false|false||Complaintnull|localized swelling in left breast|Finding|false|false||left breast swellingnull|Left breast|Anatomy|false|false||left breastnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Swelling of breast|Finding|false|false||breast swellingnull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||breastnull|Breast problem|Finding|false|false||breastnull|Procedures on breast|Procedure|false|false||breastnull|Breast|Anatomy|false|false||breastnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Evacuation of hematoma|Procedure|false|false||Evacuation of hematomanull|Evacuation procedure|Procedure|false|false||Evacuationnull|Hematoma|Finding|false|false||hematomanull|History of present illness (finding)|Finding|false|false||History of Present Illnessnull|null|Attribute|false|false||History of Present Illnessnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Present illness|Finding|false|false||Present Illnessnull|Present|Finding|false|false||Present
null|Presentation|Finding|false|false||Presentnull|Illness (finding)|Finding|false|false||Illnessnull|Woman|Subject|false|false||woman
null|Human, Female adult|Subject|false|false||womannull|ANTICOAGULATION (finding)|Finding|false|false||anticoagulation
null|Anticoagulation function|Finding|false|false||anticoagulation
null|Decreased Coagulation Activity [PE]|Finding|false|false||anticoagulationnull|Anticoagulation Therapy|Procedure|false|false||anticoagulationnull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||breastnull|Breast problem|Finding|false|false||breastnull|Procedures on breast|Procedure|false|false||breastnull|Breast|Anatomy|false|false||breastnull|Cardiomyopathy, Familial Idiopathic|Disorder|false|false||IDCnull|LMNA wt Allele|Finding|false|false||IDCnull|grade 3 education level|Finding|false|false||Grade 3
null|Tumor grade G3|Finding|false|false||Grade 3
null|Grade three rank|Finding|false|false||Grade 3
null|Simpson Grade 3|Finding|false|false||Grade 3null|Histopathologic Grade|Finding|false|false||Grade
null|Grade|Finding|false|false||Grade
null|School Grade|Finding|false|false||Gradenull|Lumpectomy of breast|Procedure|false|false||breast lumpectomynull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||breastnull|Breast problem|Finding|false|false||breastnull|Procedures on breast|Procedure|false|false||breastnull|Breast|Anatomy|false|false||breastnull|Lumpectomy of breast|Procedure|false|false||lumpectomy
null|Excision of mass (procedure)|Procedure|false|false||lumpectomynull|Sentinel Lymph Node Biopsy|Procedure|false|false||SLNBnull|localized swelling in left breast|Finding|false|false||left breast swellingnull|Left breast|Anatomy|false|false||left breastnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Swelling of breast|Finding|false|false||breast swellingnull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||breastnull|Breast problem|Finding|false|false||breastnull|Procedures on breast|Procedure|false|false||breastnull|Breast|Anatomy|false|false||breastnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Hematoma|Finding|false|false||hematomanull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Dyslipidemias|Disorder|false|false||Dyslipidemianull|Varicosity|Disorder|false|false||varicose veinsnull|Varicose|Modifier|false|false||varicosenull|Procedure on vein|Procedure|false|false||veinsnull|Veins|Anatomy|false|false||veinsnull|Ligation|Procedure|false|false||ligationnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|OSA protein, Drosophila|Drug|false|false||OSA
null|OSA protein, Drosophila|Drug|false|false||OSAnull|Sleep Apnea, Obstructive|Disorder|false|false||OSAnull|Osa <eudicots>|Entity|false|false||OSA
null|Osage language|Entity|false|false||OSA
null|Osa|Entity|false|false||OSAnull|CENPJ gene|Finding|false|false||CPapnull|Continuous Positive Airway Pressure|Procedure|false|false||CPapnull|recent upper respiratory infection|Finding|false|false||recent URInull|Recent|Time|false|false||recentnull|Upper Respiratory Infections|Disorder|false|false||URInull|Uniform Resource Identifier|Finding|false|false||URI
null|URI1 gene|Finding|false|false||URI
null|URI1 wt Allele|Finding|false|false||URInull|Course|Time|false|false||coursenull|Zithromax|Drug|false|false||Zithromax
null|Zithromax|Drug|false|false||Zithromaxnull|Bilateral|Modifier|false|false||bilateralnull|Personal Experience Scales|Finding|false|false||PEs
null|PES1 gene|Finding|false|false||PEsnull|Structure of ankle and/or foot (body structure)|Anatomy|false|false||PEs
null|Hindfoot of quadruped|Anatomy|false|false||PEs
null|Paw|Anatomy|false|false||PEs
null|Foot|Anatomy|false|false||PEsnull|Iranian Persian language|Entity|false|false||PEsnull|Antiphospholipid Syndrome|Disorder|false|false||antiphospholipid antibody syndromenull|Antiphospholipid Antibodies|Drug|false|false||antiphospholipid antibody
null|Antiphospholipid Antibodies|Drug|false|false||antiphospholipid antibodynull|Antiphospholipid antibody positivity|Finding|false|false||antiphospholipid antibodynull|Immunoglobulins|Drug|false|false||antibody
null|Immunoglobulins|Drug|false|false||antibody
null|Antibodies|Drug|false|false||antibody
null|Antibodies|Drug|false|false||antibody
null|Antibodies|Drug|false|false||antibodynull|Antibody (immunoassay)|Procedure|false|false||antibodynull|Immunoglobulin complex location, circulating|Anatomy|false|false||antibody
null|immunoglobulin complex location|Anatomy|false|false||antibodynull|Syndrome|Disorder|false|false||syndromenull|ANTICOAGULATION (finding)|Finding|false|false||anticoagulation
null|Anticoagulation function|Finding|false|false||anticoagulation
null|Decreased Coagulation Activity [PE]|Finding|false|false||anticoagulationnull|Anticoagulation Therapy|Procedure|false|false||anticoagulationnull|Last|Modifier|false|false||lastnull|United States Military enlisted E3 (qualifier value)|Finding|false|false||A1Cnull|Hemoglobin A1c measurement|Procedure|false|false||A1Cnull|Cerebral hemisphere structure (body structure)|Anatomy|false|false||cerebral
null|Brain|Anatomy|false|false||cerebralnull|Aneurysm|Finding|false|false||aneurysmnull|null|Finding|false|false||unchangednull|About The Same|Modifier|false|false||unchangednull|Gastroesophageal reflux disease|Disorder|false|false||GERDnull|Diverticulosis|Disorder|false|false||diverticulosisnull|Colonic Polyps|Disorder|true|false||colon polypsnull|Neoplasm of uncertain or unknown behavior of colon|Disorder|true|false||colon
null|Colonic Diseases|Disorder|true|false||colon
null|Carcinoma in situ of colon|Disorder|true|false||colonnull|COLON PROBLEM|Finding|true|false||colonnull|Colon structure (body structure)|Anatomy|false|false||colon
null|Abdomen+Pelvis>Colon|Anatomy|false|false||colonnull|TUBE,COLON,22FR,RADIOPAQUE RUBBER B#7370|Device|true|false||colonnull|Colon <Coloninae>|Entity|true|false||colonnull|polyps|Disorder|false|false||polypsnull|null|Finding|false|false||polypsnull|Cancer patients and suicide and depression|Disorder|false|false||depression
null|Mental Depression|Disorder|false|false||depression
null|Depressive disorder|Disorder|false|false||depression
null|Depressed mood|Disorder|false|false||depressionnull|Depression - motion|Finding|false|false||depression
null|null|Finding|false|false||depressionnull|Depression - recess|Modifier|false|false||depressionnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Candidiasis, Chronic Mucocutaneous|Disorder|false|false||CMC
null|Capillary malformation (disorder)|Disorder|false|false||CMCnull|MCC protocol|Procedure|false|false||CMCnull|Circulating Melanoma Cell|Anatomy|false|false||CMCnull|Cleveland Multiport Catheter|Device|false|false||CMCnull|Chamic Languages|Entity|false|false||CMCnull|Arthroplasty|Procedure|false|false||joint arthroplastynull|Joint problem|Finding|false|false||jointnull|null|Anatomy|false|false||joint
null|Joints|Anatomy|false|false||joint
null|Articular system|Anatomy|false|false||jointnull|Joint Device|Device|false|false||jointnull|Temporomandibular joint arthroplasty by dentist|Procedure|false|false||arthroplasty
null|Arthroplasty|Procedure|false|false||arthroplasty
null|Reconstruction of joint|Procedure|false|false||arthroplastynull|Repair of musculotendinous cuff of shoulder|Procedure|false|false||rotator cuff repairnull|Rotator Cuff|Anatomy|false|false||rotator cuffnull|null|Device|false|false||rotatornull|Cuffing (morphologic abnormality)|Finding|false|false||cuffnull|Cuff - body part|Anatomy|false|false||cuffnull|Cuff Device|Device|false|false||cuffnull|Repair|Finding|false|false||repair
null|Wound Healing|Finding|false|false||repairnull|Repair - Remedial Action|Procedure|false|false||repair
null|Surgical repair|Procedure|false|false||repairnull|Excision|Procedure|false|false||excision
null|removal technique|Procedure|false|false||excisionnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|GSC-DT gene|Finding|false|false||digitnull|Digit structure|Anatomy|false|false||digitnull|Digit - number character|LabModifier|false|false||digitnull|Mass of body structure|Finding|false|false||mass
null|Morphology, Attenuation, Size, and Structure Criteria|Finding|false|false||mass
null|null|Finding|false|false||mass
null|FBN1 wt Allele|Finding|false|false||mass
null|FBN1 gene|Finding|false|false||mass
null|Mass of body region|Finding|false|false||massnull|Mass, a measure of quantity of matter|LabModifier|false|false||mass
null|Molecular Mass|LabModifier|false|false||massnull|Calculi|Finding|false|false||stonenull|Malignant neoplasm of pancreatic duct|Disorder|false|false||pancreatic ductnull|Abdomen>Pancreatic duct|Anatomy|false|false||pancreatic duct
null|Pancreatic duct|Anatomy|false|false||pancreatic ductnull|Pancreatic Hormones|Drug|false|false||pancreatic
null|Pancreatic Hormones|Drug|false|false||pancreatic
null|Pancreatic Hormones|Drug|false|false||pancreaticnull|Pancreas|Anatomy|false|false||pancreaticnull|Duct (organ) structure|Anatomy|false|false||duct
null|canal [body parts]|Anatomy|false|false||ductnull|Duct Device|Device|false|false||ductnull|Exploration procedure|Procedure|false|false||explorationnull|Consent Type - Hysterectomy|Finding|false|false||hysterectomynull|Hysterectomy|Procedure|false|false||hysterectomynull|Tonsillectomy|Procedure|false|false||tonsillectomynull|Social and personal history|Finding|false|false||Social History
null|Social History|Finding|false|false||Social Historynull|Social|Finding|false|false||Socialnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Family Medical History|Finding|false|false||Family Historynull|Entity Name Part Type - family|Finding|false|false||Family
null|Last Name|Finding|false|false||Family
null|Living Arrangement - Family|Finding|false|false||Family
null|Family (taxonomic)|Finding|false|false||Family
null|Family Collection|Finding|false|false||Familynull|Family|Subject|false|false||Familynull|History of present illness (finding)|Finding|false|true||History
null|History of previous events|Finding|false|true||History
null|Historical aspects qualifier|Finding|false|true||History
null|Medical History|Finding|false|true||History
null|Concept History|Finding|false|true||Historynull|History|Subject|false|false||Historynull|Entity Name Part Type - family|Finding|true|false||family
null|Last Name|Finding|true|false||family
null|Living Arrangement - Family|Finding|true|false||family
null|Family (taxonomic)|Finding|true|false||family
null|Family Collection|Finding|true|false||familynull|Family|Subject|true|false||familynull|Deep thrombophlebitis|Disorder|true|false||DVT
null|Deep Vein Thrombosis|Disorder|true|false||DVTnull|area DVT|Anatomy|true|false||DVTnull|null|Attribute|true|false||DVTnull|Sister|Subject|false|false||sistersnull|Atrial Fibrillation|Disorder|false|false||atrial fibrillationnull|null|Attribute|false|false||atrial fibrillationnull|Atrial Fibrillation by ECG Finding|Lab|false|false||atrial fibrillationnull|Heart Atrium|Anatomy|false|false||atrialnull|Fibrillation|Disorder|false|false||fibrillationnull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|C1orf210 gene|Finding|false|false||Tempnull|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Procedure|false|false||Tempnull|Temperature|LabModifier|false|false||Tempnull|delivery (history)|Finding|false|false||delivery
null|Transfer Technique|Finding|false|false||delivery
null|null|Finding|false|false||deliverynull|Obstetric Delivery|Procedure|false|false||deliverynull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GEN
null|GEN1 wt Allele|Finding|false|false||GEN
null|GEN1 gene|Finding|false|false||GENnull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|Pleasant|Finding|false|false||pleasantnull|HEENT|Anatomy|false|false||HEENTnull|Scleral Diseases|Disorder|false|false||scleranull|examination of sclera|Procedure|false|false||scleranull|Sclera|Anatomy|false|false||scleranull|Anicteric|Finding|false|false||anictericnull|Pulmonary ventilator management|Procedure|false|false||PULMnull|Increased work of breathing|Finding|true|false||increased work of breathingnull|Increased (finding)|Finding|true|false||increased
null|Increase|Finding|true|false||increasednull|Increased|LabModifier|true|false||increasednull|Work of Breathing|Finding|true|false||work of breathingnull|Work|Event|true|false||worknull|outcomes otolaryngology breathing|Finding|true|false||breathing
null|Inspiration (function)|Finding|true|false||breathing
null|Respiration|Finding|true|false||breathingnull|null|Attribute|true|false||breathingnull|respiratory system process|Phenomenon|true|false||breathingnull|Feeling comfortable|Finding|true|false||comfortablenull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||BREASTnull|Breast problem|Finding|false|false||BREASTnull|Procedures on breast|Procedure|false|false||BREASTnull|Breast|Anatomy|false|false||BREASTnull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||breastnull|Breast problem|Finding|false|false||breastnull|Procedures on breast|Procedure|false|false||breastnull|Breast|Anatomy|false|false||breastnull|dependent|Finding|false|false||dependentnull|Dependent - ability|Modifier|false|false||dependent
null|Conditional|Modifier|false|false||dependentnull|Ecchymosis|Finding|false|false||ecchymosis
null|Skin Bruise|Finding|false|false||ecchymosisnull|MILDLY|Modifier|false|false||mildly
null|Mild (qualifier value)|Modifier|false|false||mildlynull|inferiority|Finding|false|false||inferiornull|Inferior|Modifier|false|false||inferiornull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||breastnull|Breast problem|Finding|false|false||breastnull|Procedures on breast|Procedure|false|false||breastnull|Breast|Anatomy|false|false||breastnull|Surgical wound|Disorder|false|false||incisionnull|Surgical incisions|Procedure|false|false||incisionnull|Cranial incision point|Anatomy|false|false||incisionnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Serosanguineous|Modifier|false|false||serosanguineousnull|system output|Finding|false|false||outputnull|Measurement of fluid output|Procedure|false|false||outputnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false||ABDnull|ABD (body structure)|Anatomy|false|false||ABD
null|Abdomen|Anatomy|false|false||ABDnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|true|false||softnull|Soft|Modifier|true|false||softnull|Hernia|Disorder|true|false||hernianull|Hereditary Multiple Exostoses|Disorder|true|false||EXTnull|EXT1 wt Allele|Finding|true|false||EXT
null|EXT1 gene|Finding|true|false||EXTnull|Feels warm|Finding|true|false||Warmnull|warming process|Phenomenon|true|false||Warmnull|Well (answer to question)|Finding|true|false||wellnull|Well (container)|Device|true|false||wellnull|Microplate Well|Modifier|true|false||well
null|Good|Modifier|true|false||well
null|Healthy|Modifier|true|false||wellnull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|Emotional tenderness|Finding|true|false||tenderness
null|Sore to touch|Finding|true|false||tendernessnull|Neurology speciality|Title|true|false||NEUROnull|Neurologic (qualifier value)|Modifier|true|false||NEUROnull|Focal Neurologic Deficits|Finding|true|false||focal neurologic deficitsnull|Focal|Modifier|true|false||focalnull|Neurologic Deficits|Finding|true|false||neurologic deficitsnull|Neurologic (qualifier value)|Modifier|true|false||neurologicnull|Deficit|Modifier|true|false||deficitsnull|Psychiatric problem|Disorder|true|false||PSYCH
null|Mental disorders|Disorder|true|false||PSYCHnull|Judgment|Finding|false|false||judgmentnull|Insight|Finding|false|false||insightnull|Memory observations|Finding|false|false||memory
null|Memory G-code|Finding|false|false||memory
null|Memory|Finding|false|false||memorynull|Memory Device|Device|false|false||memorynull|Mood (psychological function)|Finding|false|false||mood
null|mood (physical finding)|Finding|false|false||mood
null|Mood (attribute)|Finding|false|false||moodnull|null|Attribute|false|false||moodnull|Affect (mental function)|Finding|false|false||affectnull|assessment of affect|Procedure|false|false||affectnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Physical Examination|Procedure|false|false||EXAMINATION
null|Medical Examination|Procedure|false|false||EXAMINATIONnull|Examination|Event|false|false||EXAMINATIONnull|Cancer/Testis Antigen|Drug|false|false||CTAnull|PCYT1A wt Allele|Finding|false|false||CTA
null|CERNA3 gene|Finding|false|false||CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false||CTAnull|Chest problem|Finding|false|false||CHESTnull|Chest|Anatomy|false|false||CHEST
null|Anterior thoracic region|Anatomy|false|false||CHESTnull|Contrast Media|Drug|false|false||CONTRASTnull|Contrast|Modifier|false|false||CONTRASTnull|Comparison|Event|false|false||COMPARISONnull|Chest CT|Procedure|false|false||Chest CTnull|Chest problem|Finding|false|false||Chestnull|Chest|Anatomy|false|false||Chest
null|Anterior thoracic region|Anatomy|false|false||Chestnull|findings aspects|Finding|false|false||FINDINGSnull|null|Attribute|false|false||FINDINGSnull|Malignant neoplasm of heart|Disorder|false|false||HEART
null|benign neoplasm of heart|Disorder|false|false||HEARTnull|HEART PROBLEM|Finding|false|false||HEARTnull|Chest>Heart|Anatomy|false|false||HEART
null|Heart|Anatomy|false|false||HEARTnull|Vasculature|Anatomy|false|false||VASCULATUREnull|Blood supply aspects|Modifier|false|false||VASCULATUREnull|Central brand of multivitamin with minerals|Drug|true|false||central
null|Central brand of multivitamin with minerals|Drug|true|false||centralnull|Central Minus|Procedure|true|false||centralnull|Central|Modifier|true|false||centralnull|Pulmonary Embolism|Finding|true|false||pulmonary embolismnull|Pulmonary (intended site)|Finding|true|false||pulmonarynull|Lung|Anatomy|true|false||pulmonarynull|null|Attribute|true|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|true|false||pulmonarynull|Embolism|Finding|true|false||embolism
null|Embolus|Finding|true|false||embolismnull|Dissecting Thoracic Aortic Aneurysm|Disorder|true|false||thoracicnull|Chest|Anatomy|true|false||thoracicnull|Procedure on aorta|Procedure|true|false||aortanull|Chest+Abdomen>Aorta|Anatomy|true|false||aorta
null|Aorta|Anatomy|true|false||aortanull|Diameter (qualifier value)|LabModifier|true|false||calibernull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Dissecting hemorrhage|Finding|true|false||dissectionnull|Tissue Dissection|Procedure|true|false||dissectionnull|Internal|Modifier|true|false||intramuralnull|Hematoma|Finding|false|false||hematomanull|Malignant neoplasm of heart|Disorder|false|false||heart
null|benign neoplasm of heart|Disorder|false|false||heartnull|HEART PROBLEM|Finding|false|false||heartnull|Chest>Heart|Anatomy|false|false||heart
null|Heart|Anatomy|false|false||heartnull|Pericardial sac structure|Anatomy|false|false||pericardiumnull|Structure of great blood vessel (organ)|Anatomy|false|false||great vesselsnull|RXFP2 gene|Finding|false|false||greatnull|Greater|LabModifier|false|false||great
null|Large|LabModifier|false|false||greatnull|Blood Vessel|Anatomy|false|false||vesselsnull|Limited (extensiveness)|Finding|false|false||limitsnull|Pericardial effusion|Disorder|true|false||pericardial effusionnull|Pericardial effusion body substance|Finding|true|false||pericardial effusionnull|Pericardial (qualifier value)|Anatomy|true|false||pericardial
null|Pericardial sac structure|Anatomy|true|false||pericardialnull|Effusion (substance)|Finding|true|false||effusion
null|null|Finding|true|false||effusion
null|effusion|Finding|true|false||effusionnull|Axilla|Anatomy|false|false||AXILLAnull|Neoplasm of uncertain or unknown behavior of mediastinum|Disorder|false|false||MEDIASTINUM
null|Benign tumor of mediastinum|Disorder|false|false||MEDIASTINUMnull|Chest>Mediastinum|Anatomy|false|false||MEDIASTINUM
null|Mediastinum|Anatomy|false|false||MEDIASTINUMnull|Collection Object - UML Entity|Finding|false|false||collection
null|Item Collection|Finding|false|false||collection
null|Collections (publication)|Finding|false|false||collection
null|Collection (action)|Finding|false|false||collectionnull|Left breast|Anatomy|false|false||left breastnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||breastnull|Breast problem|Finding|false|false||breastnull|Procedures on breast|Procedure|false|false||breastnull|Breast|Anatomy|false|false||breastnull|density|LabModifier|false|false||densitynull|Unit - NCI Thesaurus Property|LabModifier|false|false||units
null|Unit of Measure|LabModifier|false|false||units
null|Unit|LabModifier|false|false||unitsnull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|Hematoma|Finding|false|false||hematomanull|Focal|Modifier|false|false||foci ofnull|Foci|Finding|false|false||focinull|Focal|Modifier|false|false||focinull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false||air
null|AIRN gene|Finding|false|false||air
null|AI/RHEUM|Finding|false|false||airnull|Collection Object - UML Entity|Finding|false|false||collection
null|Item Collection|Finding|false|false||collection
null|Collections (publication)|Finding|false|false||collection
null|Collection (action)|Finding|false|false||collectionnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|null|Time|false|false||priornull|Respiratory Aspiration|Disorder|false|false||aspirationnull|Aspiration into respiratory tract|Finding|false|false||aspiration
null|Endotracheal aspiration|Finding|false|false||aspiration
null|Pulmonary aspiration|Finding|false|false||aspirationnull|null|Procedure|false|false||aspirationnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Punctate|Modifier|false|false||punctatenull|Axilla|Anatomy|true|false||axillarynull|Mediastinum|Anatomy|true|false||mediastinalnull|Mediastinal|Modifier|true|false||mediastinalnull|Hilar lymphadenopathy|Disorder|true|false||hilar lymphadenopathynull|Hilar|Modifier|true|false||hilarnull|Lymphadenopathy|Disorder|false|false||lymphadenopathynull|Swollen Lymph Node|Finding|false|false||lymphadenopathynull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Structure of right axillary region|Anatomy|true|false||right axillanull|Table Cell Horizontal Align - right|Finding|true|false||rightnull|Right sided|Modifier|true|false||right
null|Right|Modifier|true|false||rightnull|Axilla|Anatomy|true|false||axillanull|Study Object|Finding|true|false||studynull|Scientific Study|Procedure|true|false||study
null|Study|Procedure|true|false||study
null|Clinical Research|Procedure|true|false||studynull|Room of building - Study|Device|true|false||studynull|Mediastinal mass|Finding|true|false||mediastinal massnull|Mediastinum|Anatomy|true|false||mediastinalnull|Mediastinal|Modifier|true|false||mediastinalnull|Mass of body structure|Finding|true|false||mass
null|Morphology, Attenuation, Size, and Structure Criteria|Finding|true|false||mass
null|null|Finding|true|false||mass
null|FBN1 wt Allele|Finding|true|false||mass
null|FBN1 gene|Finding|true|false||mass
null|Mass of body region|Finding|true|false||massnull|Mass, a measure of quantity of matter|LabModifier|true|false||mass
null|Molecular Mass|LabModifier|true|false||massnull|Pleural cavity|Anatomy|false|false||PLEURAL SPACESnull|Pleural Diseases|Disorder|false|false||PLEURALnull|Pleura|Anatomy|false|false||PLEURALnull|Pleural|Modifier|false|false||PLEURALnull|Pleural effusion (disorder)|Finding|true|false||pleural effusion
null|Pleural effusion fluid|Finding|true|false||pleural effusion
null|null|Finding|true|false||pleural effusionnull|Pleural Diseases|Disorder|true|false||pleuralnull|Pleura|Anatomy|true|false||pleuralnull|Pleural|Modifier|true|false||pleuralnull|Effusion (substance)|Finding|true|false||effusion
null|null|Finding|true|false||effusion
null|effusion|Finding|true|false||effusionnull|Pneumothorax|Disorder|true|false||pneumothoraxnull|Lung|Anatomy|false|false||LUNGSnull|Airway structure|Anatomy|false|false||AIRWAYSnull|Artificial Airways|Device|false|false||AIRWAYSnull|Lung|Anatomy|true|false||lungsnull|Remote control command - Clear|Finding|true|false||clearnull|Clear|Modifier|true|false||clear
null|Transparent (qualitative concept)|Modifier|true|false||clearnull|Areas <Spilosomini>|Entity|true|false||areasnull|Area|Modifier|true|false||areasnull|Opacification|Modifier|false|false||opacificationnull|Airway structure|Anatomy|false|false||airwaysnull|Artificial Airways|Device|false|false||airwaysnull|Legal patent|Finding|false|false||patentnull|Open|Modifier|false|false||patentnull|Segmental|Modifier|false|false||segmentalnull|Bronchi|Anatomy|false|false||bronchinull|Base of neck|Anatomy|false|false||BASE OF NECKnull|nitrogenous base|Drug|false|false||BASE
null|Base|Drug|false|false||BASE
null|Dental Base|Drug|false|false||BASE
null|base - RoleClass|Drug|false|false||BASEnull|Base - General Qualifier|Finding|false|false||BASE
null|BPIFA4P gene|Finding|false|false||BASE
null|Base - RX Component Type|Finding|false|false||BASEnull|Anatomical base|Anatomy|false|false||BASEnull|Base - unit of product usage|LabModifier|false|false||BASEnull|Passive joint movement of neck (finding)|Finding|false|false||NECK
null|Neck problem|Finding|false|false||NECKnull|dendritic spine neck|Anatomy|false|false||NECK
null|Neck|Anatomy|false|false||NECKnull|Visual|Finding|false|false||Visualizednull|nitrogenous base|Drug|true|false||base
null|Base|Drug|true|false||base
null|Dental Base|Drug|true|false||base
null|base - RoleClass|Drug|true|false||basenull|Base - General Qualifier|Finding|true|false||base
null|BPIFA4P gene|Finding|true|false||base
null|Base - RX Component Type|Finding|true|false||basenull|Anatomical base|Anatomy|true|false||basenull|Base - unit of product usage|LabModifier|true|false||basenull|Passive joint movement of neck (finding)|Finding|true|false||neck
null|Neck problem|Finding|true|false||necknull|dendritic spine neck|Anatomy|true|false||neck
null|Neck|Anatomy|true|false||necknull|Show|Entity|true|false||shownull|Congenital Abnormality|Disorder|true|false||abnormalitynull|Abnormality|Finding|true|false||abnormalitynull|Skeletal bone|Anatomy|false|false||BONES
null|XXX bone|Anatomy|false|false||BONESnull|Suspicious|Modifier|true|false||suspiciousnull|Bone Tissue, Human|Anatomy|true|false||osseous
null|Skeletal bone|Anatomy|true|false||osseousnull|Congenital Abnormality|Disorder|true|false||abnormalitynull|Abnormality|Finding|true|false||abnormalitynull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|true|false||acutenull|Fracture|Disorder|true|false||fracturenull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Left breast|Anatomy|true|false||left breastnull|Table Cell Horizontal Align - left|Finding|true|false||leftnull|Left sided|Modifier|true|false||left
null|Left|Modifier|true|false||leftnull|Breast hematoma|Finding|true|false||breast hematomanull|Neoplasm of uncertain or unknown behavior of breast|Disorder|true|false||breastnull|Breast problem|Finding|true|false||breastnull|Procedures on breast|Procedure|true|false||breastnull|Breast|Anatomy|true|false||breastnull|Hematoma|Finding|true|false||hematomanull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Hemorrhage|Finding|true|false||bleednull|Timing, LOINC Axis 3|Finding|false|false||timingnull|Timing|Time|false|false||timingnull|Suboptimal|Modifier|false|false||suboptimalnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Due to|Finding|false|false||due
null|Due|Finding|false|false||duenull|Document Completion - incomplete|Finding|false|false||incompletenull|Incomplete|Modifier|false|false||incompletenull|Partial|LabModifier|false|false||incompletenull|Knowledge Field|Finding|false|false||field
null|Force Field|Finding|false|false||field
null|Field|Finding|false|false||fieldnull|field - patient encounter|Procedure|false|false||fieldnull|View|Modifier|false|false||viewnull|Initial (abbreviation)|Finding|false|false||initialnull|Initially|Time|false|false||initialnull|Firstly|Modifier|false|false||initialnull|density|LabModifier|false|false||densitynull|Collection Object - UML Entity|Finding|false|false||collection
null|Item Collection|Finding|false|false||collection
null|Collections (publication)|Finding|false|false||collection
null|Collection (action)|Finding|false|false||collectionnull|null|Finding|false|false||unchangednull|About The Same|Modifier|false|false||unchangednull|Series|LabModifier|false|false||seriesnull|BRIEF Health Literacy Screening Tool|Finding|false|false||Brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||Briefnull|Brief|Time|false|false||Briefnull|Shortened|Modifier|false|false||Briefnull|Hospital course|Finding|false|false||Hospital Coursenull|null|Attribute|false|false||Hospital Coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||Coursenull|Woman|Subject|false|false||woman
null|Human, Female adult|Subject|false|false||womannull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||breastnull|Breast problem|Finding|false|false||breastnull|Procedures on breast|Procedure|false|false||breastnull|Breast|Anatomy|false|false||breastnull|ActInformationPrivacyReason - service|Finding|false|false||servicenull|Software Service|Device|false|false||servicenull|Services|Event|false|false||servicenull|Lumpectomy of left breast|Procedure|false|false||left breast lumpectomynull|Left breast|Anatomy|false|false||left breastnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Lumpectomy of breast|Procedure|false|false||breast lumpectomynull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||breastnull|Breast problem|Finding|false|false||breastnull|Procedures on breast|Procedure|false|false||breastnull|Breast|Anatomy|false|false||breastnull|Lumpectomy of breast|Procedure|false|false||lumpectomy
null|Excision of mass (procedure)|Procedure|false|false||lumpectomynull|Invasive|Modifier|false|false||invasivenull|Carcinoma|Disorder|false|false||carcinomanull|Recurrent|Time|false|false||recurrent
null|Episodic|Time|false|false||recurrentnull|Left breast|Anatomy|false|false||left breastnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Breast hematoma|Finding|false|false||breast hematomanull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||breastnull|Breast problem|Finding|false|false||breastnull|Procedures on breast|Procedure|false|false||breastnull|Breast|Anatomy|false|false||breastnull|Hematoma|Finding|false|false||hematomanull|null|Procedure|false|false||needle aspirationnull|Aspiration needles|Device|false|false||needle aspirationnull|null|Finding|false|false||needlenull|Needle device|Device|false|false||needlenull|Needle Shape|Modifier|false|false||needlenull|Respiratory Aspiration|Disorder|false|false||aspirationnull|Aspiration into respiratory tract|Finding|false|false||aspiration
null|Endotracheal aspiration|Finding|false|false||aspiration
null|Pulmonary aspiration|Finding|false|false||aspirationnull|null|Procedure|false|false||aspirationnull|Clinic|Device|false|false||clinic
null|Ambulatory Care Facilities|Device|false|false||clinicnull|Clinic|Entity|false|false||clinic
null|Ambulatory Care Facilities|Entity|false|false||clinicnull|Patient location type - Clinic|Modifier|false|false||clinic
null|Person location type - Clinic|Modifier|false|false||clinicnull|Examination and observation for unspecified reason|Finding|false|false||observation
null|null|Finding|false|false||observation
null|null|Finding|false|false||observation
null|Observation (finding)|Finding|false|false||observationnull|Observation - diagnostic procedure|Procedure|false|false||observation
null|Observation in research|Procedure|false|false||observation
null|Patient observation|Procedure|false|false||observationnull|Operative Surgical Procedures|Procedure|false|false||surgical
null|Surgical service|Procedure|false|false||surgicalnull|Evacuation procedure|Procedure|false|false||evacuationnull|Hematoma|Finding|false|false||hematomanull|Operating Room|Device|false|false||operating roomnull|Operating Room|Entity|false|false||operating roomnull|Patient location type - Operating Room|Modifier|false|false||operating roomnull|Operating|Finding|false|false||operatingnull|Room - Patient location type|Modifier|false|false||room
null|Room|Modifier|false|false||roomnull|Evacuation procedure|Procedure|false|false||evacuationnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Hematoma|Finding|false|false||hematomanull|Clinical act of insertion|Procedure|false|false||placement
null|Implantation procedure|Procedure|false|false||placement
null|null|Procedure|false|false||placementnull|Placement|Modifier|false|false||placementnull|Surgical drains|Device|false|false||surgical drainnull|Operative Surgical Procedures|Procedure|false|false||surgical
null|Surgical service|Procedure|false|false||surgicalnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Hospital course|Finding|false|false||Hospital coursenull|null|Attribute|false|false||Hospital coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||coursenull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Oral pain|Finding|false|false||oral painnull|Oral Dosage Form|Drug|false|false||oralnull|Oral Route of Administration|Finding|false|false||oral
null|Oral (intended site)|Finding|false|false||oralnull|Oral cavity|Anatomy|false|false||oralnull|Oral|Modifier|false|false||oralnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Acetaminophen [EPC]|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophennull|Acetaminophen measurement|Procedure|false|false||acetaminophennull|tramadol|Drug|false|false||tramadol
null|tramadol|Drug|false|false||tramadolnull|Tramadol measurement (procedure)|Procedure|false|false||tramadolnull|Taking vital signs|Procedure|false|false||Vital signsnull|null|Attribute|false|false||Vital signs
null|Vital signs|Attribute|false|false||Vital signsnull|Vital High Nitrogen Enteral Nutrition|Drug|false|false||Vitalnull|Vital (qualifier value)|Modifier|false|false||Vitalnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|per protocol|Finding|false|false||per protocol
null|On Protocol Therapy|Finding|false|false||per protocolnull|Clinical trial protocol document|Finding|false|false||protocol
null|Study Protocol|Finding|false|false||protocol
null|Protocols documentation|Finding|false|false||protocol
null|Protocol - answer to question|Finding|false|false||protocol
null|Library Protocol|Finding|false|false||protocolnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Respiratory, thoracic and mediastinal disorders|Disorder|false|false||Respnull|Respiratory rate|Attribute|false|false||Respnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|albuterol|Drug|false|false||albuterol
null|albuterol|Drug|false|false||albuterolnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|null|Finding|false|false||regular dietnull|Regular|Modifier|false|false||regularnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|NPO - Nothing by mouth|Procedure|false|false||NPOnull|null|Entity|false|false||NPOnull|Operating Room|Device|false|false||operating roomnull|Operating Room|Entity|false|false||operating roomnull|Patient location type - Operating Room|Modifier|false|false||operating roomnull|Operating|Finding|false|false||operatingnull|Room - Patient location type|Modifier|false|false||room
null|Room|Modifier|false|false||roomnull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|Perioperative Period|Time|false|false||perioperative periodnull|perioperative|Time|false|false||perioperativenull|Menstruation|Finding|false|false||periodnull|Clinical Trial Period|Procedure|false|false||periodnull|per period (qualifier value)|Time|false|false||period
null|Time periods|Time|false|false||periodnull|Transaction counts and value totals - Period|LabModifier|false|false||periodnull|Issue (document)|Finding|true|false||issue
null|Problem|Finding|true|false||issuenull|Issue (action)|Event|true|false||issuenull|Hospital course|Finding|true|false||hospital coursenull|null|Attribute|true|false||hospital coursenull|Organization unit type - Hospital|Finding|true|false||hospitalnull|Hospitals|Device|true|false||hospitalnull|Hospitals|Entity|true|false||hospitalnull|Hospital environment|Modifier|true|false||hospitalnull|Course|Time|true|false||coursenull|Heme|Drug|false|false||Heme
null|Heme|Drug|false|false||Hemenull|Daily|Time|false|false||dailynull|Laboratory test finding|Lab|false|false||labsnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|ANTICOAGULATION (finding)|Finding|false|false||anticoagulation
null|Anticoagulation function|Finding|false|false||anticoagulation
null|Decreased Coagulation Activity [PE]|Finding|false|false||anticoagulationnull|Anticoagulation Therapy|Procedure|false|false||anticoagulationnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Course|Time|false|false||coursenull|Visit User Code - Home|Finding|true|false||home
null|Address type - Home|Finding|true|false||homenull|home health encounter|Procedure|true|false||homenull|Organization unit type - Home|Entity|true|false||homenull|Person location type - Home|Modifier|true|false||home
null|Home environment|Modifier|true|false||homenull|Unit dose|LabModifier|true|false||dose
null|Dosage|LabModifier|true|false||dosenull|warfarin|Drug|true|false||warfarin
null|warfarin|Drug|true|false||warfarin
null|warfarin|Drug|true|false||warfarinnull|Body Substance Discharge|Finding|true|false||discharge
null|Discharge Body Fluid|Finding|true|false||discharge
null|Body Fluid Discharge|Finding|true|false||discharge
null|null|Finding|true|false||dischargenull|Patient Discharge|Procedure|true|false||dischargenull|Lovenox|Drug|true|false||lovenox
null|Lovenox|Drug|true|false||lovenoxnull|Fixation of dental bridge|Procedure|true|false||bridgenull|Type of bridge device|Device|true|false||bridgenull|null|Finding|false|false||compression
null|Compressed structure|Finding|false|false||compressionnull|Compression Therapy|Procedure|false|false||compression
null|Data Compression|Procedure|false|false||compressionnull|Compression|Phenomenon|false|false||compressionnull|Boots|Device|false|false||bootsnull|Boots pharmaceutical company|Entity|false|false||bootsnull|Hospital course|Finding|false|false||hospital coursenull|null|Attribute|false|false||hospital coursenull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Course|Time|false|false||coursenull|Deep thrombophlebitis|Disorder|false|false||DVTsnull|Ancef|Drug|false|false||ancef
null|Ancef|Drug|false|false||ancefnull|Prophylactic treatment|Procedure|false|false||prophylaxisnull|prevention & control|Modifier|false|false||prophylaxisnull|Apyrexial|Finding|true|false||afebrilenull|Leukocytosis|Disorder|true|false||leukocytosisnull|Blood leukocyte number above reference range|Finding|true|false||leukocytosisnull|Hospital course|Finding|true|false||hospital coursenull|null|Attribute|true|false||hospital coursenull|Organization unit type - Hospital|Finding|true|false||hospitalnull|Hospitals|Device|true|false||hospitalnull|Hospitals|Entity|true|false||hospitalnull|Hospital environment|Modifier|true|false||hospitalnull|Course|Time|false|false||coursenull|Endocrine System Diseases|Disorder|false|false||Endo
null|Endometriosis|Disorder|false|false||Endonull|MANEA gene|Finding|false|false||Endonull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Metabolic Syndrome X|Disorder|false|false||metabolic syndromenull|Metabolic Process, Cellular|Finding|false|false||metabolic
null|Metabolic|Finding|false|false||metabolicnull|Multisection metabolic|Procedure|false|false||metabolicnull|Syndrome|Disorder|false|false||syndromenull|Prediabetes syndrome|Disorder|false|false||pre-diabetesnull|Constant - dosing instruction fragment|Finding|false|false||constantnull|Constant (qualifier)|Modifier|false|false||constantnull|Carbohydrate diet|Procedure|false|false||carbohydrate dietnull|Carbohydrates|Drug|false|false||carbohydratenull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|null|Finding|false|false||regular dietnull|Regular|Modifier|false|false||regularnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Emesis [PE]|Finding|false|false||emesis
null|Vomiting|Finding|false|false||emesis
null|Vomitus|Finding|false|false||emesisnull|Emesis <Emesidini>|Entity|false|false||emesis
null|Emesis <subgenus>|Entity|false|false||emesisnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Oral pain|Finding|false|false||oral painnull|Oral Dosage Form|Drug|false|false||oralnull|Oral Route of Administration|Finding|false|false||oral
null|Oral (intended site)|Finding|false|false||oralnull|Oral cavity|Anatomy|false|false||oralnull|Oral|Modifier|false|false||oralnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Apyrexial|Finding|true|false||afebrilenull|Leukocytosis|Disorder|true|false||leukocytosisnull|Blood leukocyte number above reference range|Finding|true|false||leukocytosisnull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|true|false||antibiotics
null|Antibiotics|Drug|true|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|true|false||antibiotics
null|Antibiotics, Gynecological|Drug|true|false||antibiotics
null|antibiotics, intestinal|Drug|true|false||antibiotics
null|Antibiotic throat preparations|Drug|true|false||antibiotics
null|Antibiotics, Antitubercular|Drug|true|false||antibiotics
null|Antibiotics for systemic use|Drug|true|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|true|false||antibioticsnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Disease Management|Procedure|false|false||managementnull|Management Occupations|Subject|false|false||managementnull|Management procedure|Event|false|false||management
null|Administration occupational activities|Event|false|false||managementnull|Close|Finding|false|false||close
null|Closed|Finding|false|false||closenull|Clinic|Device|false|false||clinic
null|Ambulatory Care Facilities|Device|false|false||clinicnull|Clinic|Entity|false|false||clinic
null|Ambulatory Care Facilities|Entity|false|false||clinicnull|Patient location type - Clinic|Modifier|false|false||clinic
null|Person location type - Clinic|Modifier|false|false||clinicnull|Removal of drain|Procedure|false|false||drain removalnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|removal technique|Procedure|false|false||removal
null|Excision|Procedure|false|false||removal
null|Extraction|Procedure|false|false||removalnull|Removing (action)|Event|false|false||removalnull|Clinic|Device|false|false||clinic
null|Ambulatory Care Facilities|Device|false|false||clinicnull|Clinic|Entity|false|false||clinic
null|Ambulatory Care Facilities|Entity|false|false||clinicnull|Patient location type - Clinic|Modifier|false|false||clinic
null|Person location type - Clinic|Modifier|false|false||clinicnull|Early|Time|false|false||earlynull|Extended Priority Codes - Routine|Finding|false|false||routine
null|Report priority - Routine|Finding|false|false||routine
null|Admission Type - Routine|Finding|false|false||routine
null|Level of Care - Routine|Finding|false|false||routine
null|Processing priority - Routine|Finding|false|false||routine
null|Referral priority - Routine|Finding|false|false||routinenull|Routine coag|Procedure|false|false||routinenull|Priority - Routine|Time|false|false||routinenull|Routine|Modifier|false|false||routinenull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|Active medication list|Finding|false|false||Active Medication listnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|prescription document|Finding|false|false||Prescriptionnull|Prescription (procedure)|Procedure|false|false||Prescriptionnull|Prescription (attribute)|Attribute|false|false||Prescriptionnull|albuterol sulfate|Drug|false|false||ALBUTEROL SULFATE
null|albuterol sulfate|Drug|false|false||ALBUTEROL SULFATEnull|albuterol|Drug|false|false||ALBUTEROL
null|albuterol|Drug|false|false||ALBUTEROLnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||SULFATE
null|Sulfates, Inorganic|Drug|false|false||SULFATE
null|sulfate ion|Drug|false|false||SULFATE
null|sulfate ion|Drug|false|false||SULFATE
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||SULFATEnull|albuterol sulfate|Drug|false|false||albuterol sulfate
null|albuterol sulfate|Drug|false|false||albuterol sulfatenull|albuterol|Drug|false|false||albuterol
null|albuterol|Drug|false|false||albuterolnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfate
null|Sulfates, Inorganic|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfatenull|Solution Dosage Form|Drug|false|false||solution
null|Solutions|Drug|false|false||solution
null|Pharmaceutical Solutions|Drug|false|false||solutionnull|Resolution|Finding|false|false||solutionnull|nebulization-mediated drug administration|Procedure|false|false||nebulizationnull|Four times daily|Time|false|false||four times a daynull|Four Times|LabModifier|false|false||four timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Wheezing|Finding|false|false||wheezenull|albuterol sulfate|Drug|false|false||ALBUTEROL SULFATE
null|albuterol sulfate|Drug|false|false||ALBUTEROL SULFATEnull|albuterol|Drug|false|false||ALBUTEROL
null|albuterol|Drug|false|false||ALBUTEROLnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||SULFATE
null|Sulfates, Inorganic|Drug|false|false||SULFATE
null|sulfate ion|Drug|false|false||SULFATE
null|sulfate ion|Drug|false|false||SULFATE
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||SULFATEnull|ProAir|Drug|false|false||PROAIR HFA
null|ProAir|Drug|false|false||PROAIR HFAnull|ProAir|Drug|false|false||PROAIR
null|ProAir|Drug|false|false||PROAIR
null|Pro-Air Procaterol|Drug|false|false||PROAIR
null|Pro-Air Procaterol|Drug|false|false||PROAIRnull|Facial Hemiatrophy|Disorder|false|false||HFAnull|High frequency audiometry|Procedure|false|false||HFAnull|ProAir|Drug|false|false||ProAir HFA
null|ProAir|Drug|false|false||ProAir HFAnull|ProAir|Drug|false|false||ProAir
null|ProAir|Drug|false|false||ProAir
null|Pro-Air Procaterol|Drug|false|false||ProAir
null|Pro-Air Procaterol|Drug|false|false||ProAirnull|Facial Hemiatrophy|Disorder|false|false||HFAnull|High frequency audiometry|Procedure|false|false||HFAnull|mcg/actuation|LabModifier|false|false||mcg/actuationnull|microgram|LabModifier|false|false||mcgnull|Actuation (unit of presentation)|LabModifier|false|false||actuationnull|Aerosol Dose Form|Drug|false|false||aerosolnull|Aerosols|Device|false|false||aerosolnull|Puff Dosing Unit|LabModifier|false|false||puffsnull|Inhalation Route of Administration|Finding|false|false||inhalation
null|Inspiration (function)|Finding|false|false||inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||inhalationnull|6 Hours|Time|false|false||6 hoursnull|Hour|Time|false|false||hoursnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Wheezing|Finding|false|false||wheezenull|atorvastatin|Drug|false|false||ATORVASTATIN
null|atorvastatin|Drug|false|false||ATORVASTATINnull|atorvastatin|Drug|false|false||atorvastatin
null|atorvastatin|Drug|false|false||atorvastatinnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Once a day, at bedtime|Time|false|false||at bedtimenull|Once a day, at bedtime|Time|false|false||bedtime
null|Bedtime (qualifier value)|Time|false|false||bedtimenull|Transaction counts and value totals - provider|Finding|false|false||Provider
null|Provider|Finding|false|false||Providernull|Unit dose|LabModifier|true|false||Dose
null|Dosage|LabModifier|true|false||Dosenull|Adjustment - classification term|Finding|true|false||adjustment
null|Personal Adjustment|Finding|true|false||adjustment
null|null|Finding|true|false||adjustment
null|Psychological adjustment|Finding|true|false||adjustment
null|Transaction Type - Adjustment|Finding|true|false||adjustmentnull|Query Status Code - new|Finding|true|false||new
null|Act Status - new|Finding|true|false||newnull|Newar Language|Entity|true|false||newnull|New|Modifier|true|false||newnull|enoxaparin|Drug|false|false||ENOXAPARIN
null|enoxaparin|Drug|false|false||ENOXAPARINnull|enoxaparin|Drug|false|false||enoxaparin
null|enoxaparin|Drug|false|false||enoxaparinnull|Kilogram per Cubic Meter|LabModifier|false|false||mg/mLnull|per milliliter|LabModifier|false|false||/mLnull|Subcutaneous Route of Administration|Finding|false|false||subcutaneousnull|subcutaneous|Modifier|false|false||subcutaneousnull|Syringes|Device|false|false||syringenull|Syringe (unit of presentation)|LabModifier|false|false||syringe
null|Syringe Dosing Unit|LabModifier|false|false||syringenull|Twice a day|Time|false|false||twice dailynull|Daily|Time|false|false||dailynull|Approximate|Modifier|false|false||approximatelynull|12 hours (qualifier value)|Time|false|false||12 hoursnull|Hour|Time|false|false||hoursnull|Last|Modifier|false|false||lastnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Transaction counts and value totals - provider|Finding|false|false||Provider
null|Provider|Finding|false|false||Providernull|Unit dose|LabModifier|true|false||Dose
null|Dosage|LabModifier|true|false||Dosenull|Adjustment - classification term|Finding|true|false||adjustment
null|Personal Adjustment|Finding|true|false||adjustment
null|null|Finding|true|false||adjustment
null|Psychological adjustment|Finding|true|false||adjustment
null|Transaction Type - Adjustment|Finding|true|false||adjustmentnull|Query Status Code - new|Finding|true|false||new
null|Act Status - new|Finding|true|false||newnull|Newar Language|Entity|true|false||newnull|New|Modifier|true|false||newnull|erythromycin|Drug|false|false||ERYTHROMYCIN
null|erythromycin|Drug|false|false||ERYTHROMYCINnull|erythromycin|Drug|false|false||erythromycin
null|erythromycin|Drug|false|false||erythromycinnull|gram|LabModifier|false|false||gramnull|Ophthalmic Ointment|Drug|false|false||eye ointmentnull|Carcinoma in situ of eye|Disorder|false|false||eye
null|Disorder of eye|Disorder|false|false||eyenull|Eye - Specimen Source Code|Finding|false|false||eye
null|Eye problem|Finding|false|false||eye
null|Eye Specimen|Finding|false|false||eyenull|Head>Eye|Anatomy|false|false||eye
null|Eye|Anatomy|false|false||eye
null|Orbital region|Anatomy|false|false||eyenull|Ointments|Drug|false|false||ointmentnull|Apply (administration method)|Finding|false|false||Apply
null|Apply (instruction)|Finding|false|false||Apply
null|null|Finding|false|false||Apply
null|Apply|Finding|false|false||Applynull|Inch Unit of Length|LabModifier|false|false||inchnull|Carcinoma in situ of eye|Disorder|false|false||eye
null|Disorder of eye|Disorder|false|false||eyenull|Eye - Specimen Source Code|Finding|false|false||eye
null|Eye problem|Finding|false|false||eye
null|Eye Specimen|Finding|false|false||eyenull|Head>Eye|Anatomy|false|false||eye
null|Eye|Anatomy|false|false||eye
null|Orbital region|Anatomy|false|false||eyenull|Four times daily|Time|false|false||four times a daynull|Four Times|LabModifier|false|false||four timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|furosemide|Drug|false|false||FUROSEMIDE
null|furosemide|Drug|false|false||FUROSEMIDEnull|furosemide|Drug|false|false||furosemide
null|furosemide|Drug|false|false||furosemidenull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Swelling of lower limb|Finding|false|false||leg swellingnull|Leg|Anatomy|false|false||leg
null|Lower Extremity|Anatomy|false|false||legnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|hydromorphone|Drug|false|false||HYDROMORPHONE
null|hydromorphone|Drug|false|false||HYDROMORPHONEnull|hydromorphone|Drug|false|false||hydromorphone
null|hydromorphone|Drug|false|false||hydromorphonenull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Hour|Time|true|false||hoursnull|Severe Extremity Pain|Finding|true|false||severe pain
null|Severe pain|Finding|true|false||severe pain
null|Neck Pain Score 6|Finding|true|false||severe painnull|Severe - Severity of Illness Code|Finding|true|false||severe
null|Intensity and Distress 5|Finding|true|false||severe
null|Severe - Triage Code|Finding|true|false||severe
null|Severe (severity modifier)|Finding|true|false||severe
null|Allergy Severity - Severe|Finding|true|false||severenull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Drink (dietary substance)|Drug|true|false||drinknull|Alcohols|Drug|true|false||alcohol
null|Alcohols|Drug|true|false||alcohol
null|ethanol|Drug|true|false||alcohol
null|ethanol|Drug|true|false||alcoholnull|Alcohol - Recreational Drug Use Code|Finding|true|false||alcoholnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Nebulizers|Device|false|false||NEBULIZERnull|Compressor Air Pump Device|Device|false|false||COMPRESSORnull|Portable nebuliser system|Device|false|false||PORTABLE NEBULIZER SYSTEMnull|Portable|Modifier|false|false||PORTABLEnull|Nebulizers|Device|false|false||NEBULIZERnull|System (basic dose form)|Drug|false|false||SYSTEMnull|System, LOINC Axis 4|Finding|false|false||SYSTEM
null|System|Finding|false|false||SYSTEMnull|Device system|Device|false|false||SYSTEM
null|System - kit|Device|false|false||SYSTEMnull|System (unit of presentation)|LabModifier|false|false||SYSTEMnull|Portable|Modifier|false|false||Portablenull|Nebulizers|Device|false|false||Nebulizernull|System (basic dose form)|Drug|false|false||Systemnull|System, LOINC Axis 4|Finding|false|false||System
null|System|Finding|false|false||Systemnull|Device system|Device|false|false||System
null|System - kit|Device|false|false||Systemnull|System (unit of presentation)|LabModifier|false|false||Systemnull|Use - dosing instruction imperative|Finding|false|false||Use
null|utilization qualifier|Finding|false|false||Use
null|Usage|Finding|false|false||Usenull|albuterol|Drug|false|false||albuterol
null|albuterol|Drug|false|false||albuterolnull|Nebulizers|Device|false|false||nebulizernull|Four Times|LabModifier|false|false||four timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Wheezing|Finding|false|false||wheezenull|omeprazole|Drug|false|false||OMEPRAZOLE
null|omeprazole|Drug|false|false||OMEPRAZOLEnull|omeprazole|Drug|false|false||omeprazole
null|omeprazole|Drug|false|false||omeprazolenull|capsule (pharmacologic)|Drug|false|false||capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||capsule
null|Structure of organ capsule|Anatomy|false|false||capsulenull|Capsule Shape|Modifier|false|false||capsulenull|Capsule (unit of presentation)|LabModifier|false|false||capsule
null|Capsule Dosing Unit|LabModifier|false|false||capsulenull|Release - action (qualifier value)|Finding|false|false||release
null|Released (action)|Finding|false|false||releasenull|Discharge (release)|Procedure|false|false||release
null|Release (procedure)|Procedure|false|false||release
null|Patient Discharge|Procedure|false|false||releasenull|capsule (pharmacologic)|Drug|false|false||CAPSULEnull|Microbial anatomical capsule structure|Anatomy|false|false||CAPSULE
null|Structure of organ capsule|Anatomy|false|false||CAPSULEnull|Capsule Shape|Modifier|false|false||CAPSULEnull|Capsule (unit of presentation)|LabModifier|false|false||CAPSULE
null|Capsule Dosing Unit|LabModifier|false|false||CAPSULEnull|Twice a day|Time|false|false||TWICE DAILYnull|Daily|Time|false|false||DAILYnull|gastroesophageal|Anatomy|false|false||GASTROESOPHAGEALnull|sertraline|Drug|false|false||SERTRALINE
null|sertraline|Drug|false|false||SERTRALINEnull|sertraline|Drug|false|false||sertraline
null|sertraline|Drug|false|false||sertralinenull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|tramadol|Drug|false|false||TRAMADOL
null|tramadol|Drug|false|false||TRAMADOLnull|Tramadol measurement (procedure)|Procedure|false|false||TRAMADOLnull|tramadol|Drug|false|false||tramadol
null|tramadol|Drug|false|false||tramadolnull|Tramadol measurement (procedure)|Procedure|false|false||tramadolnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|trazodone|Drug|false|false||TRAZODONE
null|trazodone|Drug|false|false||TRAZODONEnull|trazodone|Drug|false|false||trazodone
null|trazodone|Drug|false|false||trazodonenull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Bedtime (qualifier value)|Time|false|false||bedtime
null|Once a day, at bedtime|Time|false|false||bedtimenull|warfarin|Drug|false|false||WARFARIN
null|warfarin|Drug|false|false||WARFARIN
null|warfarin|Drug|false|false||WARFARINnull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Five times weekly|Time|false|false||5 times a weeknull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Last|Modifier|false|false||lastnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|PROGRESSIVE ENCEPHALOMYELITIS WITH RIGIDITY|Disorder|false|false||pernull|Per - dosing instruction fragment|Finding|false|false||per
null|PER1 gene|Finding|false|false||per
null|Follow|Finding|false|false||per
null|PER1 wt Allele|Finding|false|false||pernull|PER (body structure)|Anatomy|false|false||pernull|Per (qualifier)|Modifier|false|false||pernull|Clinic|Device|false|false||clinic
null|Ambulatory Care Facilities|Device|false|false||clinicnull|Clinic|Entity|false|false||clinic
null|Ambulatory Care Facilities|Entity|false|false||clinicnull|Patient location type - Clinic|Modifier|false|false||clinic
null|Person location type - Clinic|Modifier|false|false||clinicnull|Transaction counts and value totals - provider|Finding|false|false||Provider
null|Provider|Finding|false|false||Providernull|Unit dose|LabModifier|true|false||Dose
null|Dosage|LabModifier|true|false||Dosenull|Adjustment - classification term|Finding|true|false||adjustment
null|Personal Adjustment|Finding|true|false||adjustment
null|null|Finding|true|false||adjustment
null|Psychological adjustment|Finding|true|false||adjustment
null|Transaction Type - Adjustment|Finding|true|false||adjustmentnull|Query Status Code - new|Finding|true|false||new
null|Act Status - new|Finding|true|false||newnull|Newar Language|Entity|true|false||newnull|New|Modifier|true|false||newnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|Drugs, Non-Prescription|Drug|false|false||OTCnull|OTC gene|Finding|false|false||OTCnull|Acetaminophen [EPC]|Drug|false|false||ACETAMINOPHEN
null|acetaminophen|Drug|false|false||ACETAMINOPHEN
null|acetaminophen|Drug|false|false||ACETAMINOPHENnull|Acetaminophen measurement|Procedure|false|false||ACETAMINOPHENnull|Acetaminophen [EPC]|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophennull|Acetaminophen measurement|Procedure|false|false||acetaminophennull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|3 times|Finding|false|false||3 timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Daily|Time|false|false||dailynull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Multiple Epiphyseal Dysplasia|Disorder|false|false||mednull|Master of Education|Finding|false|false||med
null|COMP wt Allele|Finding|false|false||med
null|COL9A3 gene|Finding|false|false||med
null|SCN8A wt Allele|Finding|false|false||med
null|COL9A2 gene|Finding|false|false||med
null|COMP gene|Finding|false|false||med
null|SCN8A gene|Finding|false|false||mednull|ZDHHC2 protein, human|Drug|false|false||rec
null|ZDHHC2 protein, human|Drug|false|false||recnull|RBPJP4 gene|Finding|false|false||rec
null|MCM8 gene|Finding|false|false||recnull|cholecalciferol|Drug|false|false||CHOLECALCIFEROL (VITAMIN D3)
null|cholecalciferol|Drug|false|false||CHOLECALCIFEROL (VITAMIN D3)
null|cholecalciferol|Drug|false|false||CHOLECALCIFEROL (VITAMIN D3)null|cholecalciferol|Drug|false|false||CHOLECALCIFEROL
null|cholecalciferol|Drug|false|false||CHOLECALCIFEROL
null|cholecalciferol|Drug|false|false||CHOLECALCIFEROLnull|vitamin D3|Drug|false|false||VITAMIN D3
null|vitamin D3|Drug|false|false||VITAMIN D3
null|cholecalciferol|Drug|false|false||VITAMIN D3
null|cholecalciferol|Drug|false|false||VITAMIN D3
null|cholecalciferol|Drug|false|false||VITAMIN D3null|Vitamins|Drug|false|false||VITAMIN
null|Vitamins|Drug|false|false||VITAMIN
null|Vitamins|Drug|false|false||VITAMINnull|cholecalciferol|Drug|false|false||cholecalciferol (vitamin D3)
null|cholecalciferol|Drug|false|false||cholecalciferol (vitamin D3)
null|cholecalciferol|Drug|false|false||cholecalciferol (vitamin D3)null|cholecalciferol|Drug|false|false||cholecalciferol
null|cholecalciferol|Drug|false|false||cholecalciferol
null|cholecalciferol|Drug|false|false||cholecalciferolnull|vitamin D3|Drug|false|false||vitamin D3
null|vitamin D3|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitaminnull|Storage Unit|Device|false|false||unit
null|Unit device|Device|false|false||unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||unit
null|Unit of Measure|LabModifier|false|false||unit
null|Unit|LabModifier|false|false||unit
null|Enzyme Unit|LabModifier|false|false||unitnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Drugs, Non-Prescription|Drug|false|false||OTCnull|OTC gene|Finding|false|false||OTCnull|polyethylene glycol 3350|Drug|false|false||POLYETHYLENE GLYCOL 3350
null|polyethylene glycol 3350|Drug|false|false||POLYETHYLENE GLYCOL 3350null|polyethylene glycols|Drug|false|false||POLYETHYLENE GLYCOL
null|polyethylene glycols|Drug|false|false||POLYETHYLENE GLYCOLnull|high-density polyethylene|Drug|false|false||POLYETHYLENE
null|high-density polyethylene|Drug|false|false||POLYETHYLENE
null|polyethylenes|Drug|false|false||POLYETHYLENE
null|polyethylenes|Drug|false|false||POLYETHYLENE
null|Polyethylene|Drug|false|false||POLYETHYLENE
null|Polyethylene|Drug|false|false||POLYETHYLENEnull|ethylene glycol|Drug|false|false||GLYCOL
null|Glycol|Drug|false|false||GLYCOL
null|ethylene glycol|Drug|false|false||GLYCOL
null|Glycols|Drug|false|false||GLYCOLnull|Miralax|Drug|false|false||MIRALAX
null|Miralax|Drug|false|false||MIRALAXnull|Miralax|Drug|false|false||Miralax
null|Miralax|Drug|false|false||Miralaxnull|gram|LabModifier|false|false||gramnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Oral Dosage Form|Drug|false|false||oralnull|Oral Route of Administration|Finding|false|false||oral
null|Oral (intended site)|Finding|false|false||oralnull|Oral cavity|Anatomy|false|false||oralnull|Oral|Modifier|false|false||oralnull|powder physical state|Drug|false|false||powder
null|Powder dose form|Drug|false|false||powdernull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Constipation|Finding|false|false||constipationnull|Transaction counts and value totals - provider|Finding|false|false||Provider
null|Provider|Finding|false|false||Providernull|Dose Adjustment|Procedure|true|false||Dose adjustmentnull|Unit dose|LabModifier|true|false||Dose
null|Dosage|LabModifier|true|false||Dosenull|Adjustment - classification term|Finding|true|false||adjustment
null|Personal Adjustment|Finding|true|false||adjustment
null|null|Finding|true|false||adjustment
null|Psychological adjustment|Finding|true|false||adjustment
null|Transaction Type - Adjustment|Finding|true|false||adjustmentnull|Query Status Code - new|Finding|true|false||new
null|Act Status - new|Finding|true|false||newnull|Newar Language|Entity|true|false||newnull|New|Modifier|true|false||newnull|sennosides, USP|Drug|false|false||SENNOSIDES
null|sennosides, USP|Drug|false|false||SENNOSIDESnull|sennosides, USP|Drug|false|false||SENNA
null|sennosides, USP|Drug|false|false||SENNAnull|Senna alexandrina|Entity|false|false||SENNA
null|Senna Plant|Entity|false|false||SENNAnull|sennosides, USP|Drug|false|false||senna
null|sennosides, USP|Drug|false|false||sennanull|Senna alexandrina|Entity|false|false||senna
null|Senna Plant|Entity|false|false||sennanull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Constipation|Finding|false|false||constipationnull|Drugs, Non-Prescription|Drug|false|false||OTCnull|OTC gene|Finding|false|false||OTCnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|tramadol|Drug|false|false||TraMADol
null|tramadol|Drug|false|false||TraMADolnull|Tramadol measurement (procedure)|Procedure|false|false||TraMADolnull|Every four hours|Time|false|false||Q4Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Moderate - Severity of Illness Code|Finding|false|false||Moderate
null|Moderate|Finding|false|false||Moderatenull|Moderate (severity modifier)|Modifier|false|false||Moderate
null|Moderate - Allergy Severity|Modifier|false|false||Moderate
null|Moderation|Modifier|false|false||Moderatenull|Indication of (contextual qualifier)|Finding|false|false||Reason fornull|Indication of (contextual qualifier)|Finding|false|false||Reasonnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Duplicate component (foundation metadata concept)|Finding|false|false||duplicate
null|Double (qualifier value)|Finding|false|false||duplicatenull|Replicate|Event|false|false||duplicatenull|Duplicate|Modifier|false|false||duplicatenull|Override|Finding|false|false||overridenull|Similarity|Modifier|false|false||similarnull|With intensity|Modifier|false|false||severity
null|Severities|Modifier|false|false||severitynull|tramadol|Drug|false|false||tramadol
null|tramadol|Drug|false|false||tramadolnull|Tramadol measurement (procedure)|Procedure|false|false||tramadolnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|CIAO3 gene|Finding|false|false||prnnull|As required|Time|false|false||prn
null|Pro Re Nata|Time|false|false||prnnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|omeprazole|Drug|false|false||Omeprazole
null|omeprazole|Drug|false|false||Omeprazolenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|sennosides, USP|Drug|false|false||Senna
null|sennosides, USP|Drug|false|false||Sennanull|Senna alexandrina|Entity|false|false||Senna
null|Senna Plant|Entity|false|false||Sennanull|sertraline|Drug|false|false||Sertraline
null|sertraline|Drug|false|false||Sertralinenull|Daily|Time|false|false||DAILYnull|trazodone|Drug|false|false||TraZODone
null|trazodone|Drug|false|false||TraZODonenull|Once a day, at bedtime|Time|false|false||QHSnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleep
null|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleepnull|Sleep|Finding|false|false||sleepnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Breast hematoma|Finding|false|false||breast hematomanull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||breastnull|Breast problem|Finding|false|false||breastnull|Procedures on breast|Procedure|false|false||breastnull|Breast|Anatomy|false|false||breastnull|Hematoma|Finding|false|false||hematomanull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Disease|Disorder|false|false||Conditionnull|Logical Condition|Finding|false|false||Conditionnull|null|Attribute|false|false||Conditionnull|Condition|Modifier|false|false||Conditionnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|Discharge instructions|Finding|false|false||Discharge Instructionsnull|hospital discharge instructions (treatment)|Procedure|false|false||Discharge Instructionsnull|null|Attribute|false|false||Discharge Instructionsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|Self-care interventions|Finding|false|false||Personal Carenull|Personal Attribute|Subject|false|false||Personalnull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|Surgical incisions|Procedure|false|false||incisionsnull|Open|Modifier|false|false||opennull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false||air
null|AIRN gene|Finding|false|false||air
null|AI/RHEUM|Finding|false|false||airnull|Cleaning (activity)|Event|false|false||cleannull|Sterility, Reproductive|Finding|false|false||sterile
null|Infertility|Finding|false|false||sterilenull|Sterile (qualifier value)|Modifier|false|false||sterilenull|Gauzes|Device|false|false||gauzenull|Daily|Time|false|false||dailynull|Cleaning (activity)|Event|false|false||Cleannull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|null|Finding|false|false||sitenull|Anatomic Site|Anatomy|false|false||sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Tubing|Device|false|false||tubingnull|Skin and subcutaneous tissue disorders|Disorder|false|false||skin
null|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||skinnull|Skin Specimen Source Code|Finding|false|false||skin
null|Skin Specimen|Finding|false|false||skinnull|Skin, Human|Anatomy|false|false||skin
null|Skin|Anatomy|false|false||skinnull|Soap Dosage Form|Drug|false|false||soapnull|Soap|Device|false|false||soapnull|Water Specimen|Drug|false|false||water
null|water|Drug|false|false||water
null|water|Drug|false|false||waternull|Water - Specimen Source Codes|Finding|false|false||waternull|Hydrotherapy|Procedure|false|false||waternull|Compliance Package - Strip|Drug|false|false||Strip
null|Strip Dosage Form|Drug|false|false||Stripnull|strip medical device|Device|false|false||Stripnull|Strip - unit of product usage|LabModifier|false|false||Strip
null|Strip (unit of presentation)|LabModifier|false|false||Strip
null|Strip Dosing Unit|LabModifier|false|false||Stripnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Tubing|Device|false|false||tubingnull|Exhausted|Finding|false|false||emptynull|Empty (qualifier)|Modifier|false|false||emptynull|anatomical bulb|Anatomy|false|false||bulb
null|Medulla Oblongata|Anatomy|false|false||bulbnull|plant bulb|Entity|false|false||bulbnull|Records|Finding|false|false||recordnull|Record - QueryRequestLimit|LabModifier|false|false||recordnull|system output|Finding|false|false||outputnull|Measurement of fluid output|Procedure|false|false||outputnull|times/day|LabModifier|false|false||times per daynull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|per day|Time|false|false||per daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|written - ParticipationMode|Finding|false|false||written
null|Written - Consent Mode|Finding|false|false||writtennull|Record of (contextual qualifier)|Modifier|false|false||record ofnull|Records|Finding|false|false||recordnull|Record - QueryRequestLimit|LabModifier|false|false||recordnull|Daily|Time|false|false||dailynull|system output|Finding|false|false||outputnull|Measurement of fluid output|Procedure|false|false||outputnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Follow-up status|Finding|false|false||follow-upnull|follow-up|Procedure|false|false||follow-upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|Appointments|Event|false|false||appointmentnull|Drain device|Device|false|false||drainsnull|As soon as possible|Time|false|false||as soon as possiblenull|Possible|Finding|false|false||possiblenull|Possibly Related to Intervention|Modifier|false|false||possible
null|Possible diagnosis|Modifier|false|false||possiblenull|Daily|Time|false|false||dailynull|system output|Finding|false|false||outputnull|Measurement of fluid output|Procedure|false|false||outputnull|Acceptable (foundation metadata concept)|Modifier|false|false||acceptable
null|Acceptable|Modifier|false|false||acceptablenull|Amount class - Amount|Finding|false|false||amountnull|Quantity|LabModifier|false|false||amountnull|Operative Surgical Procedures|Procedure|false|false||surgical
null|Surgical service|Procedure|false|false||surgicalnull|Brain|Anatomy|false|false||branull|Brassiere|Device|false|false||branull|Braj Language|Entity|false|false||branull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|Loose|Modifier|false|false||loosenull|Camisole|Device|false|false||camisolenull|Comfort brand of hydroxyethyl cellulose|Drug|false|false||comfort
null|Comfort brand of hydroxyethyl cellulose|Drug|false|false||comfortnull|Comfort|Finding|false|false||comfortnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|DERMABOND|Drug|false|false||Dermabond
null|DERMABOND|Drug|false|false||Dermabondnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false||skinnull|Skin Specimen Source Code|Finding|false|false||skin
null|Skin Specimen|Finding|false|false||skinnull|Skin, Human|Anatomy|false|false||skin
null|Skin|Anatomy|false|false||skinnull|Glues|Drug|false|false||gluenull|day|Time|false|false||daysnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|null|Finding|false|false||regular dietnull|Regular|Modifier|false|false||regularnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Walking (function)|Finding|false|false||Walknull|More than once a day|Time|false|false||several times a daynull|Several|LabModifier|false|false||severalnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Pounds|LabModifier|true|false||poundsnull|Strenuous Exercise|Finding|false|false||strenuous activitynull|Strenuous|Modifier|false|false||strenuousnull|Activity (animal life circumstance)|Finding|false|false||activity
null|Physical activity|Finding|false|false||activitynull|Activities|Event|false|false||activitynull|null|Modifier|false|false||activitynull|6 weeks|Time|false|false||6 weeksnull|week|Time|false|false||weeksnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|Resume - Remote control command|Finding|false|false||Resume
null|Curriculum Vitae|Finding|false|false||Resume
null|resume - DataOperation|Finding|false|false||Resumenull|Regular|Modifier|false|false||regularnull|Pharmaceutical Preparations|Drug|true|false||medicationsnull|Medications|Finding|true|false||medicationsnull|null|Attribute|true|false||medications
null|null|Attribute|true|false||medicationsnull|Query Status Code - new|Finding|true|false||new
null|Act Status - new|Finding|true|false||newnull|Newar Language|Entity|true|false||newnull|New|Modifier|true|false||newnull|MICROCEPHALY, EPILEPSY, AND DIABETES SYNDROME 1|Disorder|true|false||medsnull|Medications|Finding|true|false||medsnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Moderate - Severity of Illness Code|Finding|false|false||moderate
null|Moderate|Finding|false|false||moderatenull|Moderate (severity modifier)|Modifier|false|false||moderate
null|Moderate - Allergy Severity|Modifier|false|false||moderate
null|Moderation|Modifier|false|false||moderatenull|Severe Extremity Pain|Finding|false|false||severe pain
null|Severe pain|Finding|false|false||severe pain
null|Neck Pain Score 6|Finding|false|false||severe painnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Tylenol|Drug|false|false||Tylenol
null|Tylenol|Drug|false|false||Tylenolnull|Tylenol Extra Strength|Drug|false|false||Extra Strength Tylenol
null|Tylenol Extra Strength|Drug|false|false||Extra Strength Tylenolnull|Strength (attribute)|Finding|false|false||Strengthnull|Pharmaceutical Strength|LabModifier|false|false||Strength
null|Physical Strength|LabModifier|false|false||Strengthnull|Tylenol|Drug|false|false||Tylenol
null|Tylenol|Drug|false|false||Tylenolnull|Mild pain|Finding|false|false||mild pain
null|Neck Pain Score 2|Finding|false|false||mild painnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Packaging Materials|Device|false|false||packaging
null|Drug Packaging|Device|false|false||packagingnull|Packaging|Phenomenon|false|false||packagingnull|Packing (action)|Event|false|false||packagingnull|Percocet|Drug|false|false||Percocet
null|Percocet|Drug|false|false||Percocetnull|Vicodin|Drug|false|false||Vicodin
null|Vicodin|Drug|false|false||Vicodinnull|Tylenol|Drug|false|false||Tylenol
null|Tylenol|Drug|false|false||Tylenolnull|Active ingredient|Drug|true|false||active ingredientnull|Has active ingredient|Modifier|true|false||active ingredientnull|Ingredient|Drug|true|false||ingredientnull|MICROCEPHALY, EPILEPSY, AND DIABETES SYNDROME 1|Disorder|true|false||medsnull|Medications|Finding|true|false||medsnull|Additional|Finding|true|false||additionalnull|Tylenol|Drug|true|false||Tylenol
null|Tylenol|Drug|true|false||Tylenolnull|prescription document|Finding|true|false||prescriptionnull|Prescription (procedure)|Procedure|true|false||prescriptionnull|Prescription (attribute)|Attribute|true|false||prescriptionnull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Pharmaceutical Preparations|Drug|true|false||medicationsnull|Medications|Finding|true|false||medicationsnull|null|Attribute|true|false||medications
null|null|Attribute|true|false||medicationsnull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Tylenol|Drug|true|false||Tylenol
null|Tylenol|Drug|true|false||Tylenolnull|Colace|Drug|false|false||Colace
null|Colace|Drug|false|false||Colacenull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|2 times per day|Finding|false|false||2 times per daynull|2 times|Finding|false|false||2 timesnull|times/day|LabModifier|false|false||times per daynull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|per day|Time|false|false||per daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|prescription document|Finding|false|false||prescriptionnull|Prescription (procedure)|Procedure|false|false||prescriptionnull|Prescription (attribute)|Attribute|false|false||prescriptionnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Different|Modifier|false|false||differentnull|Counter brand of Terbufos|Drug|false|false||counter
null|Counter brand of Terbufos|Drug|false|false||counternull|Counter device|Device|false|false||counternull|Stool Softener brand of docusate sodium|Drug|false|false||stool softener
null|Stool Softener brand of docusate sodium|Drug|false|false||stool softener
null|Stool Softener|Drug|false|false||stool softenernull|Feces|Finding|false|false||stoolnull|Stool seat|Device|false|false||stoolnull|heavy machinery|Device|true|false||heavy machinerynull|Heavy (weight) (qualifier value)|Modifier|true|false||heavy
null|Heavy (amount)|Modifier|true|false||heavynull|Contact with machinery|Disorder|true|false||machinerynull|Industrial machine|Device|true|false||machinerynull|Narcotics|Drug|true|false||narcotic
null|Narcotics|Drug|true|false||narcoticnull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Pharmaceutical Preparations|Drug|true|false||medicationnull|medication - HL7 publishing domain|Finding|true|false||medication
null|Medications|Finding|true|false||medicationnull|Have Constipation|Finding|false|false||have constipationnull|Constipation|Finding|false|false||constipationnull|Narcotics|Drug|false|false||narcotic
null|Narcotics|Drug|false|false||narcoticnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|oxycodone|Drug|false|false||oxycodone
null|oxycodone|Drug|false|false||oxycodonenull|Oxycodone measurement|Procedure|false|false||oxycodonenull|Percocet|Drug|false|false||percocet
null|Percocet|Drug|false|false||percocetnull|Vicodin|Drug|false|false||vicodin
null|Vicodin|Drug|false|false||vicodinnull|hydrocodone|Drug|false|false||hydrocodone
null|hydrocodone|Drug|false|false||hydrocodonenull|Dilaudid|Drug|false|false||dilaudid
null|Dilaudid|Drug|false|false||dilaudidnull|Etc.|Finding|false|false||etcnull|Drinking (function)|Finding|false|false||drinking
null|Alcohol consumption|Finding|false|false||drinkingnull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|Stool Softener|Drug|false|false||stool softenersnull|Feces|Finding|false|false||stoolnull|Stool seat|Device|false|false||stoolnull|Food|Drug|false|false||foodsnull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Fiber brand of calcium polycarbophil|Drug|false|false||fiber
null|fiber|Drug|false|false||fiber
null|fiber|Drug|false|false||fiber
null|Fiber brand of calcium polycarbophil|Drug|false|false||fibernull|Tissue fiber|Anatomy|false|false||fibernull|Fiber Device|Device|false|false||fibernull|Animal in fiber production|Entity|false|false||fiber
null|Plant fiber|Entity|false|false||fibernull|Address type - Office|Finding|false|false||officenull|Office|Device|false|false||officenull|Organization unit type - Office|Entity|false|false||officenull|Stat (do immediately)|Time|false|false||IMMEDIATELYnull|Following|Time|true|false||following
null|Status post|Time|true|false||followingnull|Aspects of signs|Finding|false|false||Signs
null|Physical findings|Finding|false|false||Signsnull|Manufactured sign|Device|false|false||Signsnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Fever with chills|Finding|false|false||fever with chillsnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Chills|Finding|false|false||chillsnull|Erythema|Disorder|false|false||rednessnull|Redness|Finding|false|false||rednessnull|Red color|Modifier|false|false||rednessnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Physiologic warmth|Finding|false|false||warmth
null|Social warmth|Finding|false|false||warmthnull|Emotional tenderness|Finding|false|false||tenderness
null|Sore to touch|Finding|false|false||tendernessnull|Operative site|Modifier|false|false||surgical sitenull|Operative Surgical Procedures|Procedure|false|false||surgical
null|Surgical service|Procedure|false|false||surgicalnull|null|Finding|false|false||sitenull|Anatomic Site|Anatomy|false|false||sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Unusual|Modifier|false|false||unusualnull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|Surgical wound|Disorder|false|false||incisionnull|Surgical incisions|Procedure|false|false||incisionnull|Cranial incision point|Anatomy|false|false||incisionnull|Large amount|LabModifier|false|false||large amountnull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|Amount class - Amount|Finding|false|false||amountnull|Quantity|LabModifier|false|false||amountnull|Hemorrhage|Finding|false|false||bleedingnull|Surgical wound|Disorder|false|false||incisionnull|Surgical incisions|Procedure|false|false||incisionnull|Cranial incision point|Anatomy|false|false||incisionnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Fever symptoms (finding)|Finding|false|false||Fever
null|Fever|Finding|false|false||Fevernull|Greater Than|LabModifier|true|false||greater thannull|Greater|LabModifier|false|false||greaternull|Severe Extremity Pain|Finding|true|false||Severe pain
null|Severe pain|Finding|true|false||Severe pain
null|Neck Pain Score 6|Finding|true|false||Severe painnull|Severe - Severity of Illness Code|Finding|true|false||Severe
null|Intensity and Distress 5|Finding|true|false||Severe
null|Severe - Triage Code|Finding|true|false||Severe
null|Severe (severity modifier)|Finding|true|false||Severe
null|Allergy Severity - Severe|Finding|true|false||Severenull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Pharmaceutical Preparations|Drug|true|false||medicationnull|medication - HL7 publishing domain|Finding|true|false||medication
null|Medications|Finding|true|false||medicationnull|Vomiting|Finding|true|false||vomitingnull|Liquid substance|Drug|true|false||fluidsnull|Mouse Body Fluid or Substance|Finding|true|false||fluidsnull|Fluid Therapy|Procedure|true|false||fluidsnull|Pharmaceutical Preparations|Drug|true|false||medicationsnull|Medications|Finding|true|false||medicationsnull|null|Attribute|true|false||medications
null|null|Attribute|true|false||medicationsnull|Chills|Finding|false|false||chillsnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Greater Than|LabModifier|false|false||greater thannull|Greater|LabModifier|false|false||greaternull|Academic degree|Finding|false|false||degreesnull|Degree or extent|LabModifier|false|false||degreesnull|Academic degree|Finding|false|false||degreesnull|Degree or extent|LabModifier|false|false||degreesnull|Increased (finding)|Finding|false|false||increased
null|Increase|Finding|false|false||increasednull|Increased|LabModifier|false|false||increasednull|Erythema|Disorder|false|false||rednessnull|Redness|Finding|false|false||rednessnull|Red color|Modifier|false|false||rednessnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Surgical wound|Disorder|false|false||incisionnull|Surgical incisions|Procedure|false|false||incisionnull|Cranial incision point|Anatomy|false|false||incisionnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Dyspnea|Finding|false|false||shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false||breathnull|Else|Finding|false|false||elsenull|Equipment Alert Level - Serious|Finding|true|false||serious
null|Device Alert Level - Serious|Finding|true|false||serious
null|Alert level - Serious|Finding|true|false||seriousnull|Serious|Modifier|true|false||seriousnull|Changing|Finding|true|false||change innull|Changed status|LabModifier|true|false||change innull|Changing|Finding|true|false||changenull|Change - procedure|Procedure|true|false||changenull|Delta (difference)|LabModifier|true|false||change
null|Changed status|LabModifier|true|false||changenull|Symptoms aspect|Finding|true|false||symptoms
null|Symptoms|Finding|true|false||symptomsnull|Query Status Code - new|Finding|true|false||new
null|Act Status - new|Finding|true|false||newnull|Newar Language|Entity|true|false||newnull|New|Modifier|true|false||newnull|Symptoms aspect|Finding|true|false||symptoms
null|Symptoms|Finding|true|false||symptomsnull|Concern|Finding|true|false||concernnull|ANTICOAGULATION (finding)|Finding|false|false||ANTICOAGULATION
null|Anticoagulation function|Finding|false|false||ANTICOAGULATION
null|Decreased Coagulation Activity [PE]|Finding|false|false||ANTICOAGULATIONnull|Anticoagulation Therapy|Procedure|false|false||ANTICOAGULATIONnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|warfarin dose|Procedure|false|false||warfarin dosenull|null|Attribute|false|false||warfarin dosenull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Evening|Time|false|false||eveningnull|Resume - Remote control command|Finding|false|false||resume
null|Curriculum Vitae|Finding|false|false||resume
null|resume - DataOperation|Finding|false|false||resumenull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|Regular|Modifier|false|false||regularnull|Dosage|LabModifier|false|false||dosesnull|Bridge Therapy|Procedure|true|false||bridge therapynull|Fixation of dental bridge|Procedure|true|false||bridgenull|Type of bridge device|Device|true|false||bridgenull|Therapy Object (animal model)|Finding|true|false||therapy
null|therapeutic aspects|Finding|true|false||therapynull|Therapeutic procedure|Procedure|true|false||therapynull|warfarin|Drug|true|false||warfarin
null|warfarin|Drug|true|false||warfarin
null|warfarin|Drug|true|false||warfarinnull|Drain - SpecimenType|Drug|false|false||DRAINnull|Drain Specimen Code|Finding|false|false||DRAINnull|Drain device|Device|false|false||DRAINnull|Discharge instructions|Finding|false|false||DISCHARGE INSTRUCTIONSnull|hospital discharge instructions (treatment)|Procedure|false|false||DISCHARGE INSTRUCTIONSnull|null|Attribute|false|false||DISCHARGE INSTRUCTIONSnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Instructions|Finding|false|false||INSTRUCTIONS
null|Instruction [Publication Type]|Finding|false|false||INSTRUCTIONSnull|null|Attribute|false|false||INSTRUCTIONSnull|Drain device|Device|false|false||drainsnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Drain - SpecimenType|Drug|false|false||Drainnull|Drain Specimen Code|Finding|false|false||Drainnull|Drain device|Device|false|false||Drainnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Cleaning (activity)|Event|false|false||cleannull|Procedure (set of actions)|Finding|false|false||procedurenull|Interventional procedure|Procedure|false|false||procedurenull|null|Attribute|false|false||procedurenull|Act Class - procedure|Event|false|false||procedurenull|Hand|Anatomy|false|false||handsnull|Thoroughly|Finding|false|false||thoroughlynull|Soap Dosage Form|Drug|false|false||soapnull|Soap|Device|false|false||soapnull|Feels warm|Finding|false|false||warmnull|warming process|Phenomenon|false|false||warmnull|Water Specimen|Drug|false|false||water
null|water|Drug|false|false||water
null|water|Drug|false|false||waternull|Water - Specimen Source Codes|Finding|false|false||waternull|Hydrotherapy|Procedure|false|false||waternull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Exhausted|Finding|false|false||emptynull|Empty (qualifier)|Modifier|false|false||emptynull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Daily|Time|false|false||each daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Does pull|Finding|false|false||Pullnull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|null|Device|false|false||bottlenull|Bottle (unit of presentation)|LabModifier|false|false||bottle
null|Bottle Dosing Unit|LabModifier|false|false||bottlenull|Exhausted|Finding|false|false||emptynull|Empty (qualifier)|Modifier|false|false||emptynull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Carcinoma of unknown primary|Disorder|false|false||cupnull|Cup (physical object)|Device|false|false||cup
null|Cup Device|Device|false|false||cupnull|Cup (unit of presentation)|LabModifier|false|false||cup
null|Cup Dosing Unit|LabModifier|false|false||cupnull|Amount class - Amount|Finding|false|false||amountnull|Quantity|LabModifier|false|false||amountnull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Records|Finding|false|false||recordnull|Record - QueryRequestLimit|LabModifier|false|false||recordnull|Suction drain|Device|false|false||drain suctionnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Suction drainage|Procedure|false|false||suctionnull|Location Equipment - Suction|Modifier|false|false||suctionnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Daily|Time|false|false||dailynull|Event Log|Finding|false|false||lognull|lateral occipital gyrus (human only)|Anatomy|false|false||lognull|Logarithm|LabModifier|false|false||lognull|Individual - insurance coverage level|Finding|false|false||individualnull|Individual|Subject|false|false||individual
null|Persons|Subject|false|false||individualnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Appointments|Event|false|false||appointmentnull|null|Attribute|false|false||surgeonnull|Surgeon|Subject|false|false||surgeonnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions